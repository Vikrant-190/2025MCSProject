* File: netlist.sp
* Created: Sat Jun 14 09:12:51 2025
* Program "Calibre xRC"
* Version "v2019.2_26.18"
* 
.include "netlist.sp.pex"
.subckt SRAMnSA_1  VSS BL<15> VDD BLN<15> BL<14> BLN<14> BL<13> BLN<13> BL<12>
+ BLN<12> BL_S<15> BL_S<14> BL_S<13> BL_S<12> BLN_S<15> BLN_S<14> BLN_S<13>
+ BLN_S<12> BL<11> BLN<11> BL<10> BLN<10> BL<9> BLN<9> BL<8> BLN<8> BL_S<11>
+ BL_S<10> BL_S<9> BL_S<8> BLN_S<11> BLN_S<10> BLN_S<9> BLN_S<8> BL<7> BLN<7>
+ BL<6> BLN<6> BL<5> BLN<5> BL<4> BLN<4> BL_S<7> BL_S<6> BL_S<5> BL_S<4>
+ BLN_S<7> BLN_S<6> BLN_S<5> BLN_S<4> BL<3> BLN<3> BL<2> BLN<2> BL<1> BLN<1>
+ BL<0> BLN<0> BL_S<3> BL_S<2> BL_S<1> BL_S<0> BLN_S<3> BLN_S<2> BLN_S<1>
+ BLN_S<0> SA_EN WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> WL<6> WL<7> WL<8> WL<9>
+ WL<10> WL<11> WL<12> WL<13> WL<14> WL<15> WL<16> WL<17> WL<18> WL<19> WL<20>
+ WL<21> WL<22> WL<23> WL<24> WL<25> WL<26> WL<27> WL<28> WL<29> WL<30> WL<31>
+ WL<32> WL<33> WL<34> WL<35> WL<36> WL<37> WL<38> WL<39> WL<40> WL<41> WL<42>
+ WL<43> WL<44> WL<45> WL<46> WL<47> WL<48> WL<49> WL<50> WL<51> WL<52> WL<53>
+ WL<54> WL<55> WL<56> WL<57> WL<58> WL<59> WL<60> WL<61> WL<62> WL<63> WL<64>
+ WL<65> WL<66> WL<67> WL<68> WL<69> WL<70> WL<71> WL<72> WL<73> WL<74> WL<75>
+ WL<76> WL<77> WL<78> WL<79> WL<80> WL<81> WL<82> WL<83> WL<84> WL<85> WL<86>
+ WL<87> WL<88> WL<89> WL<90> WL<91> WL<92> WL<93> WL<94> WL<95> WL<96> WL<97>
+ WL<98> WL<99> WL<100> WL<101> WL<102> WL<103> WL<104> WL<105> WL<106> WL<107>
+ WL<108> WL<109> WL<110> WL<111> WL<112> WL<113> WL<114> WL<115> WL<116>
+ WL<117> WL<118> WL<119> WL<120> WL<121> WL<122> WL<123> WL<124> WL<125>
+ WL<126> WL<127>
* 
* WL<127>	WL<127>
* WL<126>	WL<126>
* WL<125>	WL<125>
* WL<124>	WL<124>
* WL<123>	WL<123>
* WL<122>	WL<122>
* WL<121>	WL<121>
* WL<120>	WL<120>
* WL<119>	WL<119>
* WL<118>	WL<118>
* WL<117>	WL<117>
* WL<116>	WL<116>
* WL<115>	WL<115>
* WL<114>	WL<114>
* WL<113>	WL<113>
* WL<112>	WL<112>
* WL<111>	WL<111>
* WL<110>	WL<110>
* WL<109>	WL<109>
* WL<108>	WL<108>
* WL<107>	WL<107>
* WL<106>	WL<106>
* WL<105>	WL<105>
* WL<104>	WL<104>
* WL<103>	WL<103>
* WL<102>	WL<102>
* WL<101>	WL<101>
* WL<100>	WL<100>
* WL<99>	WL<99>
* WL<98>	WL<98>
* WL<97>	WL<97>
* WL<96>	WL<96>
* WL<95>	WL<95>
* WL<94>	WL<94>
* WL<93>	WL<93>
* WL<92>	WL<92>
* WL<91>	WL<91>
* WL<90>	WL<90>
* WL<89>	WL<89>
* WL<88>	WL<88>
* WL<87>	WL<87>
* WL<86>	WL<86>
* WL<85>	WL<85>
* WL<84>	WL<84>
* WL<83>	WL<83>
* WL<82>	WL<82>
* WL<81>	WL<81>
* WL<80>	WL<80>
* WL<79>	WL<79>
* WL<78>	WL<78>
* WL<77>	WL<77>
* WL<76>	WL<76>
* WL<75>	WL<75>
* WL<74>	WL<74>
* WL<73>	WL<73>
* WL<72>	WL<72>
* WL<71>	WL<71>
* WL<70>	WL<70>
* WL<69>	WL<69>
* WL<68>	WL<68>
* WL<67>	WL<67>
* WL<66>	WL<66>
* WL<65>	WL<65>
* WL<64>	WL<64>
* WL<63>	WL<63>
* WL<62>	WL<62>
* WL<61>	WL<61>
* WL<60>	WL<60>
* WL<59>	WL<59>
* WL<58>	WL<58>
* WL<57>	WL<57>
* WL<56>	WL<56>
* WL<55>	WL<55>
* WL<54>	WL<54>
* WL<53>	WL<53>
* WL<52>	WL<52>
* WL<51>	WL<51>
* WL<50>	WL<50>
* WL<49>	WL<49>
* WL<48>	WL<48>
* WL<47>	WL<47>
* WL<46>	WL<46>
* WL<45>	WL<45>
* WL<44>	WL<44>
* WL<43>	WL<43>
* WL<42>	WL<42>
* WL<41>	WL<41>
* WL<40>	WL<40>
* WL<39>	WL<39>
* WL<38>	WL<38>
* WL<37>	WL<37>
* WL<36>	WL<36>
* WL<35>	WL<35>
* WL<34>	WL<34>
* WL<33>	WL<33>
* WL<32>	WL<32>
* WL<31>	WL<31>
* WL<30>	WL<30>
* WL<29>	WL<29>
* WL<28>	WL<28>
* WL<27>	WL<27>
* WL<26>	WL<26>
* WL<25>	WL<25>
* WL<24>	WL<24>
* WL<23>	WL<23>
* WL<22>	WL<22>
* WL<21>	WL<21>
* WL<20>	WL<20>
* WL<19>	WL<19>
* WL<18>	WL<18>
* WL<17>	WL<17>
* WL<16>	WL<16>
* WL<15>	WL<15>
* WL<14>	WL<14>
* WL<13>	WL<13>
* WL<12>	WL<12>
* WL<11>	WL<11>
* WL<10>	WL<10>
* WL<9>	WL<9>
* WL<8>	WL<8>
* WL<7>	WL<7>
* WL<6>	WL<6>
* WL<5>	WL<5>
* WL<4>	WL<4>
* WL<3>	WL<3>
* WL<2>	WL<2>
* WL<1>	WL<1>
* WL<0>	WL<0>
* SA_EN	SA_EN
* BLN_S<0>	BLN_S<0>
* BLN_S<1>	BLN_S<1>
* BLN_S<2>	BLN_S<2>
* BLN_S<3>	BLN_S<3>
* BL_S<0>	BL_S<0>
* BL_S<1>	BL_S<1>
* BL_S<2>	BL_S<2>
* BL_S<3>	BL_S<3>
* BLN<0>	BLN<0>
* BL<0>	BL<0>
* BLN<1>	BLN<1>
* BL<1>	BL<1>
* BLN<2>	BLN<2>
* BL<2>	BL<2>
* BLN<3>	BLN<3>
* BL<3>	BL<3>
* BLN_S<4>	BLN_S<4>
* BLN_S<5>	BLN_S<5>
* BLN_S<6>	BLN_S<6>
* BLN_S<7>	BLN_S<7>
* BL_S<4>	BL_S<4>
* BL_S<5>	BL_S<5>
* BL_S<6>	BL_S<6>
* BL_S<7>	BL_S<7>
* BLN<4>	BLN<4>
* BL<4>	BL<4>
* BLN<5>	BLN<5>
* BL<5>	BL<5>
* BLN<6>	BLN<6>
* BL<6>	BL<6>
* BLN<7>	BLN<7>
* BL<7>	BL<7>
* BLN_S<8>	BLN_S<8>
* BLN_S<9>	BLN_S<9>
* BLN_S<10>	BLN_S<10>
* BLN_S<11>	BLN_S<11>
* BL_S<8>	BL_S<8>
* BL_S<9>	BL_S<9>
* BL_S<10>	BL_S<10>
* BL_S<11>	BL_S<11>
* BLN<8>	BLN<8>
* BL<8>	BL<8>
* BLN<9>	BLN<9>
* BL<9>	BL<9>
* BLN<10>	BLN<10>
* BL<10>	BL<10>
* BLN<11>	BLN<11>
* BL<11>	BL<11>
* BLN_S<12>	BLN_S<12>
* BLN_S<13>	BLN_S<13>
* BLN_S<14>	BLN_S<14>
* BLN_S<15>	BLN_S<15>
* BL_S<12>	BL_S<12>
* BL_S<13>	BL_S<13>
* BL_S<14>	BL_S<14>
* BL_S<15>	BL_S<15>
* BLN<12>	BLN<12>
* BL<12>	BL<12>
* BLN<13>	BLN<13>
* BL<13>	BL<13>
* BLN<14>	BLN<14>
* BL<14>	BL<14>
* BLN<15>	BLN<15>
* VDD	VDD
* BL<15>	BL<15>
* VSS	VSS
mXI1/XI0/MM1 N_BLN_S<15>_XI1/XI0/MM1_d N_BL_S<15>_XI1/XI0/MM1_g
+ N_XI1/XI0/NET3_XI1/XI0/MM1_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI0/MM0 N_BL_S<15>_XI1/XI0/MM0_d N_BLN_S<15>_XI1/XI0/MM0_g
+ N_XI1/XI0/NET3_XI1/XI0/MM0_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI0/MM2 N_XI1/XI0/NET3_XI1/XI0/MM2_d N_SA_EN_XI1/XI0/MM2_g
+ N_VSS_XI1/XI0/MM2_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM6 N_BL_S<15>_XI1/XI0/MM6_d N_SA_EN_XI1/XI0/MM6_g
+ N_BL<15>_XI1/XI0/MM6_s N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM4 N_BLN_S<15>_XI1/XI0/MM4_d N_BL_S<15>_XI1/XI0/MM4_g
+ N_VDD_XI1/XI0/MM4_s N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM3 N_BL_S<15>_XI1/XI0/MM3_d N_BLN_S<15>_XI1/XI0/MM3_g
+ N_VDD_XI1/XI0/MM3_s N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM5 N_BLN_S<15>_XI1/XI0/MM5_d N_SA_EN_XI1/XI0/MM5_g
+ N_BLN<15>_XI1/XI0/MM5_s N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM1 N_BLN_S<14>_XI1/XI4/MM1_d N_BL_S<14>_XI1/XI4/MM1_g
+ N_XI1/XI4/NET3_XI1/XI4/MM1_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI4/MM0 N_BL_S<14>_XI1/XI4/MM0_d N_BLN_S<14>_XI1/XI4/MM0_g
+ N_XI1/XI4/NET3_XI1/XI4/MM0_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI4/MM2 N_XI1/XI4/NET3_XI1/XI4/MM2_d N_SA_EN_XI1/XI4/MM2_g
+ N_VSS_XI1/XI4/MM2_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM6 N_BL_S<14>_XI1/XI4/MM6_d N_SA_EN_XI1/XI4/MM6_g
+ N_BL<14>_XI1/XI4/MM6_s N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM4 N_BLN_S<14>_XI1/XI4/MM4_d N_BL_S<14>_XI1/XI4/MM4_g
+ N_VDD_XI1/XI4/MM4_s N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM3 N_BL_S<14>_XI1/XI4/MM3_d N_BLN_S<14>_XI1/XI4/MM3_g
+ N_VDD_XI1/XI4/MM3_s N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM5 N_BLN_S<14>_XI1/XI4/MM5_d N_SA_EN_XI1/XI4/MM5_g
+ N_BLN<14>_XI1/XI4/MM5_s N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM1 N_BLN_S<13>_XI1/XI8/MM1_d N_BL_S<13>_XI1/XI8/MM1_g
+ N_XI1/XI8/NET3_XI1/XI8/MM1_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI8/MM0 N_BL_S<13>_XI1/XI8/MM0_d N_BLN_S<13>_XI1/XI8/MM0_g
+ N_XI1/XI8/NET3_XI1/XI8/MM0_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI8/MM2 N_XI1/XI8/NET3_XI1/XI8/MM2_d N_SA_EN_XI1/XI8/MM2_g
+ N_VSS_XI1/XI8/MM2_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM6 N_BL_S<13>_XI1/XI8/MM6_d N_SA_EN_XI1/XI8/MM6_g
+ N_BL<13>_XI1/XI8/MM6_s N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM4 N_BLN_S<13>_XI1/XI8/MM4_d N_BL_S<13>_XI1/XI8/MM4_g
+ N_VDD_XI1/XI8/MM4_s N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM3 N_BL_S<13>_XI1/XI8/MM3_d N_BLN_S<13>_XI1/XI8/MM3_g
+ N_VDD_XI1/XI8/MM3_s N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM5 N_BLN_S<13>_XI1/XI8/MM5_d N_SA_EN_XI1/XI8/MM5_g
+ N_BLN<13>_XI1/XI8/MM5_s N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM1 N_BLN_S<12>_XI1/XI12/MM1_d N_BL_S<12>_XI1/XI12/MM1_g
+ N_XI1/XI12/NET3_XI1/XI12/MM1_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI12/MM0 N_BL_S<12>_XI1/XI12/MM0_d N_BLN_S<12>_XI1/XI12/MM0_g
+ N_XI1/XI12/NET3_XI1/XI12/MM0_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI12/MM2 N_XI1/XI12/NET3_XI1/XI12/MM2_d N_SA_EN_XI1/XI12/MM2_g
+ N_VSS_XI1/XI12/MM2_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM6 N_BL_S<12>_XI1/XI12/MM6_d N_SA_EN_XI1/XI12/MM6_g
+ N_BL<12>_XI1/XI12/MM6_s N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI12/MM4 N_BLN_S<12>_XI1/XI12/MM4_d N_BL_S<12>_XI1/XI12/MM4_g
+ N_VDD_XI1/XI12/MM4_s N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM3 N_BL_S<12>_XI1/XI12/MM3_d N_BLN_S<12>_XI1/XI12/MM3_g
+ N_VDD_XI1/XI12/MM3_s N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM5 N_BLN_S<12>_XI1/XI12/MM5_d N_SA_EN_XI1/XI12/MM5_g
+ N_BLN<12>_XI1/XI12/MM5_s N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI1/MM1 N_BLN_S<11>_XI1/XI1/MM1_d N_BL_S<11>_XI1/XI1/MM1_g
+ N_XI1/XI1/NET3_XI1/XI1/MM1_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI1/MM0 N_BL_S<11>_XI1/XI1/MM0_d N_BLN_S<11>_XI1/XI1/MM0_g
+ N_XI1/XI1/NET3_XI1/XI1/MM0_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI1/MM2 N_XI1/XI1/NET3_XI1/XI1/MM2_d N_SA_EN_XI1/XI1/MM2_g
+ N_VSS_XI1/XI1/MM2_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM6 N_BL_S<11>_XI1/XI1/MM6_d N_SA_EN_XI1/XI1/MM6_g
+ N_BL<11>_XI1/XI1/MM6_s N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM4 N_BLN_S<11>_XI1/XI1/MM4_d N_BL_S<11>_XI1/XI1/MM4_g
+ N_VDD_XI1/XI1/MM4_s N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM3 N_BL_S<11>_XI1/XI1/MM3_d N_BLN_S<11>_XI1/XI1/MM3_g
+ N_VDD_XI1/XI1/MM3_s N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM5 N_BLN_S<11>_XI1/XI1/MM5_d N_SA_EN_XI1/XI1/MM5_g
+ N_BLN<11>_XI1/XI1/MM5_s N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM1 N_BLN_S<10>_XI1/XI5/MM1_d N_BL_S<10>_XI1/XI5/MM1_g
+ N_XI1/XI5/NET3_XI1/XI5/MM1_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI5/MM0 N_BL_S<10>_XI1/XI5/MM0_d N_BLN_S<10>_XI1/XI5/MM0_g
+ N_XI1/XI5/NET3_XI1/XI5/MM0_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI5/MM2 N_XI1/XI5/NET3_XI1/XI5/MM2_d N_SA_EN_XI1/XI5/MM2_g
+ N_VSS_XI1/XI5/MM2_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM6 N_BL_S<10>_XI1/XI5/MM6_d N_SA_EN_XI1/XI5/MM6_g
+ N_BL<10>_XI1/XI5/MM6_s N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM4 N_BLN_S<10>_XI1/XI5/MM4_d N_BL_S<10>_XI1/XI5/MM4_g
+ N_VDD_XI1/XI5/MM4_s N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM3 N_BL_S<10>_XI1/XI5/MM3_d N_BLN_S<10>_XI1/XI5/MM3_g
+ N_VDD_XI1/XI5/MM3_s N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM5 N_BLN_S<10>_XI1/XI5/MM5_d N_SA_EN_XI1/XI5/MM5_g
+ N_BLN<10>_XI1/XI5/MM5_s N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM1 N_BLN_S<9>_XI1/XI9/MM1_d N_BL_S<9>_XI1/XI9/MM1_g
+ N_XI1/XI9/NET3_XI1/XI9/MM1_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI9/MM0 N_BL_S<9>_XI1/XI9/MM0_d N_BLN_S<9>_XI1/XI9/MM0_g
+ N_XI1/XI9/NET3_XI1/XI9/MM0_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI9/MM2 N_XI1/XI9/NET3_XI1/XI9/MM2_d N_SA_EN_XI1/XI9/MM2_g
+ N_VSS_XI1/XI9/MM2_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM6 N_BL_S<9>_XI1/XI9/MM6_d N_SA_EN_XI1/XI9/MM6_g N_BL<9>_XI1/XI9/MM6_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM4 N_BLN_S<9>_XI1/XI9/MM4_d N_BL_S<9>_XI1/XI9/MM4_g
+ N_VDD_XI1/XI9/MM4_s N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM3 N_BL_S<9>_XI1/XI9/MM3_d N_BLN_S<9>_XI1/XI9/MM3_g
+ N_VDD_XI1/XI9/MM3_s N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM5 N_BLN_S<9>_XI1/XI9/MM5_d N_SA_EN_XI1/XI9/MM5_g
+ N_BLN<9>_XI1/XI9/MM5_s N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM1 N_BLN_S<8>_XI1/XI13/MM1_d N_BL_S<8>_XI1/XI13/MM1_g
+ N_XI1/XI13/NET3_XI1/XI13/MM1_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI13/MM0 N_BL_S<8>_XI1/XI13/MM0_d N_BLN_S<8>_XI1/XI13/MM0_g
+ N_XI1/XI13/NET3_XI1/XI13/MM0_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI13/MM2 N_XI1/XI13/NET3_XI1/XI13/MM2_d N_SA_EN_XI1/XI13/MM2_g
+ N_VSS_XI1/XI13/MM2_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM6 N_BL_S<8>_XI1/XI13/MM6_d N_SA_EN_XI1/XI13/MM6_g
+ N_BL<8>_XI1/XI13/MM6_s N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM4 N_BLN_S<8>_XI1/XI13/MM4_d N_BL_S<8>_XI1/XI13/MM4_g
+ N_VDD_XI1/XI13/MM4_s N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM3 N_BL_S<8>_XI1/XI13/MM3_d N_BLN_S<8>_XI1/XI13/MM3_g
+ N_VDD_XI1/XI13/MM3_s N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM5 N_BLN_S<8>_XI1/XI13/MM5_d N_SA_EN_XI1/XI13/MM5_g
+ N_BLN<8>_XI1/XI13/MM5_s N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI2/MM1 N_BLN_S<7>_XI1/XI2/MM1_d N_BL_S<7>_XI1/XI2/MM1_g
+ N_XI1/XI2/NET3_XI1/XI2/MM1_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI2/MM0 N_BL_S<7>_XI1/XI2/MM0_d N_BLN_S<7>_XI1/XI2/MM0_g
+ N_XI1/XI2/NET3_XI1/XI2/MM0_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI2/MM2 N_XI1/XI2/NET3_XI1/XI2/MM2_d N_SA_EN_XI1/XI2/MM2_g
+ N_VSS_XI1/XI2/MM2_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM6 N_BL_S<7>_XI1/XI2/MM6_d N_SA_EN_XI1/XI2/MM6_g N_BL<7>_XI1/XI2/MM6_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM4 N_BLN_S<7>_XI1/XI2/MM4_d N_BL_S<7>_XI1/XI2/MM4_g
+ N_VDD_XI1/XI2/MM4_s N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM3 N_BL_S<7>_XI1/XI2/MM3_d N_BLN_S<7>_XI1/XI2/MM3_g
+ N_VDD_XI1/XI2/MM3_s N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM5 N_BLN_S<7>_XI1/XI2/MM5_d N_SA_EN_XI1/XI2/MM5_g
+ N_BLN<7>_XI1/XI2/MM5_s N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM1 N_BLN_S<6>_XI1/XI6/MM1_d N_BL_S<6>_XI1/XI6/MM1_g
+ N_XI1/XI6/NET3_XI1/XI6/MM1_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI6/MM0 N_BL_S<6>_XI1/XI6/MM0_d N_BLN_S<6>_XI1/XI6/MM0_g
+ N_XI1/XI6/NET3_XI1/XI6/MM0_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI6/MM2 N_XI1/XI6/NET3_XI1/XI6/MM2_d N_SA_EN_XI1/XI6/MM2_g
+ N_VSS_XI1/XI6/MM2_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM6 N_BL_S<6>_XI1/XI6/MM6_d N_SA_EN_XI1/XI6/MM6_g N_BL<6>_XI1/XI6/MM6_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM4 N_BLN_S<6>_XI1/XI6/MM4_d N_BL_S<6>_XI1/XI6/MM4_g
+ N_VDD_XI1/XI6/MM4_s N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM3 N_BL_S<6>_XI1/XI6/MM3_d N_BLN_S<6>_XI1/XI6/MM3_g
+ N_VDD_XI1/XI6/MM3_s N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM5 N_BLN_S<6>_XI1/XI6/MM5_d N_SA_EN_XI1/XI6/MM5_g
+ N_BLN<6>_XI1/XI6/MM5_s N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM1 N_BLN_S<5>_XI1/XI10/MM1_d N_BL_S<5>_XI1/XI10/MM1_g
+ N_XI1/XI10/NET3_XI1/XI10/MM1_s N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI10/MM0 N_BL_S<5>_XI1/XI10/MM0_d N_BLN_S<5>_XI1/XI10/MM0_g
+ N_XI1/XI10/NET3_XI1/XI10/MM0_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI10/MM2 N_XI1/XI10/NET3_XI1/XI10/MM2_d N_SA_EN_XI1/XI10/MM2_g
+ N_VSS_XI1/XI10/MM2_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM6 N_BL_S<5>_XI1/XI10/MM6_d N_SA_EN_XI1/XI10/MM6_g
+ N_BL<5>_XI1/XI10/MM6_s N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM4 N_BLN_S<5>_XI1/XI10/MM4_d N_BL_S<5>_XI1/XI10/MM4_g
+ N_VDD_XI1/XI10/MM4_s N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM3 N_BL_S<5>_XI1/XI10/MM3_d N_BLN_S<5>_XI1/XI10/MM3_g
+ N_VDD_XI1/XI10/MM3_s N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM5 N_BLN_S<5>_XI1/XI10/MM5_d N_SA_EN_XI1/XI10/MM5_g
+ N_BLN<5>_XI1/XI10/MM5_s N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI14/MM1 N_BLN_S<4>_XI1/XI14/MM1_d N_BL_S<4>_XI1/XI14/MM1_g
+ N_XI1/XI14/NET3_XI1/XI14/MM1_s N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI14/MM0 N_BL_S<4>_XI1/XI14/MM0_d N_BLN_S<4>_XI1/XI14/MM0_g
+ N_XI1/XI14/NET3_XI1/XI14/MM0_s N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI14/MM2 N_XI1/XI14/NET3_XI1/XI14/MM2_d N_SA_EN_XI1/XI14/MM2_g
+ N_VSS_XI1/XI14/MM2_s N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM6 N_BL_S<4>_XI1/XI14/MM6_d N_SA_EN_XI1/XI14/MM6_g
+ N_BL<4>_XI1/XI14/MM6_s N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM4 N_BLN_S<4>_XI1/XI14/MM4_d N_BL_S<4>_XI1/XI14/MM4_g
+ N_VDD_XI1/XI14/MM4_s N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM3 N_BL_S<4>_XI1/XI14/MM3_d N_BLN_S<4>_XI1/XI14/MM3_g
+ N_VDD_XI1/XI14/MM3_s N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM5 N_BLN_S<4>_XI1/XI14/MM5_d N_SA_EN_XI1/XI14/MM5_g
+ N_BLN<4>_XI1/XI14/MM5_s N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI3/MM1 N_BLN_S<3>_XI1/XI3/MM1_d N_BL_S<3>_XI1/XI3/MM1_g
+ N_XI1/XI3/NET3_XI1/XI3/MM1_s N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI3/MM0 N_BL_S<3>_XI1/XI3/MM0_d N_BLN_S<3>_XI1/XI3/MM0_g
+ N_XI1/XI3/NET3_XI1/XI3/MM0_s N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI3/MM2 N_XI1/XI3/NET3_XI1/XI3/MM2_d N_SA_EN_XI1/XI3/MM2_g
+ N_VSS_XI1/XI3/MM2_s N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM6 N_BL_S<3>_XI1/XI3/MM6_d N_SA_EN_XI1/XI3/MM6_g N_BL<3>_XI1/XI3/MM6_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM4 N_BLN_S<3>_XI1/XI3/MM4_d N_BL_S<3>_XI1/XI3/MM4_g
+ N_VDD_XI1/XI3/MM4_s N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM3 N_BL_S<3>_XI1/XI3/MM3_d N_BLN_S<3>_XI1/XI3/MM3_g
+ N_VDD_XI1/XI3/MM3_s N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM5 N_BLN_S<3>_XI1/XI3/MM5_d N_SA_EN_XI1/XI3/MM5_g
+ N_BLN<3>_XI1/XI3/MM5_s N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM1 N_BLN_S<2>_XI1/XI7/MM1_d N_BL_S<2>_XI1/XI7/MM1_g
+ N_XI1/XI7/NET3_XI1/XI7/MM1_s N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI7/MM0 N_BL_S<2>_XI1/XI7/MM0_d N_BLN_S<2>_XI1/XI7/MM0_g
+ N_XI1/XI7/NET3_XI1/XI7/MM0_s N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI7/MM2 N_XI1/XI7/NET3_XI1/XI7/MM2_d N_SA_EN_XI1/XI7/MM2_g
+ N_VSS_XI1/XI7/MM2_s N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM6 N_BL_S<2>_XI1/XI7/MM6_d N_SA_EN_XI1/XI7/MM6_g N_BL<2>_XI1/XI7/MM6_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM4 N_BLN_S<2>_XI1/XI7/MM4_d N_BL_S<2>_XI1/XI7/MM4_g
+ N_VDD_XI1/XI7/MM4_s N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM3 N_BL_S<2>_XI1/XI7/MM3_d N_BLN_S<2>_XI1/XI7/MM3_g
+ N_VDD_XI1/XI7/MM3_s N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM5 N_BLN_S<2>_XI1/XI7/MM5_d N_SA_EN_XI1/XI7/MM5_g
+ N_BLN<2>_XI1/XI7/MM5_s N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM1 N_BLN_S<1>_XI1/XI11/MM1_d N_BL_S<1>_XI1/XI11/MM1_g
+ N_XI1/XI11/NET3_XI1/XI11/MM1_s N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI11/MM0 N_BL_S<1>_XI1/XI11/MM0_d N_BLN_S<1>_XI1/XI11/MM0_g
+ N_XI1/XI11/NET3_XI1/XI11/MM0_s N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI11/MM2 N_XI1/XI11/NET3_XI1/XI11/MM2_d N_SA_EN_XI1/XI11/MM2_g
+ N_VSS_XI1/XI11/MM2_s N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM6 N_BL_S<1>_XI1/XI11/MM6_d N_SA_EN_XI1/XI11/MM6_g
+ N_BL<1>_XI1/XI11/MM6_s N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM4 N_BLN_S<1>_XI1/XI11/MM4_d N_BL_S<1>_XI1/XI11/MM4_g
+ N_VDD_XI1/XI11/MM4_s N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM3 N_BL_S<1>_XI1/XI11/MM3_d N_BLN_S<1>_XI1/XI11/MM3_g
+ N_VDD_XI1/XI11/MM3_s N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM5 N_BLN_S<1>_XI1/XI11/MM5_d N_SA_EN_XI1/XI11/MM5_g
+ N_BLN<1>_XI1/XI11/MM5_s N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI1/XI15/MM1 N_BLN_S<0>_XI1/XI15/MM1_d N_BL_S<0>_XI1/XI15/MM1_g
+ N_XI1/XI15/NET3_XI1/XI15/MM1_s N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI15/MM0 N_BL_S<0>_XI1/XI15/MM0_d N_BLN_S<0>_XI1/XI15/MM0_g
+ N_XI1/XI15/NET3_XI1/XI15/MM0_s N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
mXI1/XI15/MM2 N_XI1/XI15/NET3_XI1/XI15/MM2_d N_SA_EN_XI1/XI15/MM2_g
+ N_VSS_XI1/XI15/MM2_s N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM6 N_BL_S<0>_XI1/XI15/MM6_d N_SA_EN_XI1/XI15/MM6_g
+ N_BL<0>_XI1/XI15/MM6_s N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM4 N_BLN_S<0>_XI1/XI15/MM4_d N_BL_S<0>_XI1/XI15/MM4_g
+ N_VDD_XI1/XI15/MM4_s N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM3 N_BL_S<0>_XI1/XI15/MM3_d N_BLN_S<0>_XI1/XI15/MM3_g
+ N_VDD_XI1/XI15/MM3_s N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM5 N_BLN_S<0>_XI1/XI15/MM5_d N_SA_EN_XI1/XI15/MM5_g
+ N_BLN<0>_XI1/XI15/MM5_s N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08
+ NFIN=1
mXI0/XI0/XI0/MM2 N_XI0/XI0/XI0/NET34_XI0/XI0/XI0/MM2_d
+ N_XI0/XI0/XI0/NET33_XI0/XI0/XI0/MM2_g N_VSS_XI0/XI0/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI0/MM3 N_XI0/XI0/XI0/NET33_XI0/XI0/XI0/MM3_d N_WL<0>_XI0/XI0/XI0/MM3_g
+ N_BLN<15>_XI0/XI0/XI0/MM3_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI0/MM0 N_XI0/XI0/XI0/NET34_XI0/XI0/XI0/MM0_d N_WL<0>_XI0/XI0/XI0/MM0_g
+ N_BL<15>_XI0/XI0/XI0/MM0_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI0/MM1 N_XI0/XI0/XI0/NET33_XI0/XI0/XI0/MM1_d
+ N_XI0/XI0/XI0/NET34_XI0/XI0/XI0/MM1_g N_VSS_XI0/XI0/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI0/MM9 N_XI0/XI0/XI0/NET36_XI0/XI0/XI0/MM9_d N_WL<1>_XI0/XI0/XI0/MM9_g
+ N_BL<15>_XI0/XI0/XI0/MM9_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI0/MM6 N_XI0/XI0/XI0/NET35_XI0/XI0/XI0/MM6_d
+ N_XI0/XI0/XI0/NET36_XI0/XI0/XI0/MM6_g N_VSS_XI0/XI0/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI0/MM7 N_XI0/XI0/XI0/NET36_XI0/XI0/XI0/MM7_d
+ N_XI0/XI0/XI0/NET35_XI0/XI0/XI0/MM7_g N_VSS_XI0/XI0/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI0/MM8 N_XI0/XI0/XI0/NET35_XI0/XI0/XI0/MM8_d N_WL<1>_XI0/XI0/XI0/MM8_g
+ N_BLN<15>_XI0/XI0/XI0/MM8_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI0/MM5 N_XI0/XI0/XI0/NET34_XI0/XI0/XI0/MM5_d
+ N_XI0/XI0/XI0/NET33_XI0/XI0/XI0/MM5_g N_VDD_XI0/XI0/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI0/MM4 N_XI0/XI0/XI0/NET33_XI0/XI0/XI0/MM4_d
+ N_XI0/XI0/XI0/NET34_XI0/XI0/XI0/MM4_g N_VDD_XI0/XI0/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI0/MM10 N_XI0/XI0/XI0/NET35_XI0/XI0/XI0/MM10_d
+ N_XI0/XI0/XI0/NET36_XI0/XI0/XI0/MM10_g N_VDD_XI0/XI0/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI0/MM11 N_XI0/XI0/XI0/NET36_XI0/XI0/XI0/MM11_d
+ N_XI0/XI0/XI0/NET35_XI0/XI0/XI0/MM11_g N_VDD_XI0/XI0/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI1/MM2 N_XI0/XI0/XI1/NET34_XI0/XI0/XI1/MM2_d
+ N_XI0/XI0/XI1/NET33_XI0/XI0/XI1/MM2_g N_VSS_XI0/XI0/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI1/MM3 N_XI0/XI0/XI1/NET33_XI0/XI0/XI1/MM3_d N_WL<0>_XI0/XI0/XI1/MM3_g
+ N_BLN<14>_XI0/XI0/XI1/MM3_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI1/MM0 N_XI0/XI0/XI1/NET34_XI0/XI0/XI1/MM0_d N_WL<0>_XI0/XI0/XI1/MM0_g
+ N_BL<14>_XI0/XI0/XI1/MM0_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI1/MM1 N_XI0/XI0/XI1/NET33_XI0/XI0/XI1/MM1_d
+ N_XI0/XI0/XI1/NET34_XI0/XI0/XI1/MM1_g N_VSS_XI0/XI0/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI1/MM9 N_XI0/XI0/XI1/NET36_XI0/XI0/XI1/MM9_d N_WL<1>_XI0/XI0/XI1/MM9_g
+ N_BL<14>_XI0/XI0/XI1/MM9_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI1/MM6 N_XI0/XI0/XI1/NET35_XI0/XI0/XI1/MM6_d
+ N_XI0/XI0/XI1/NET36_XI0/XI0/XI1/MM6_g N_VSS_XI0/XI0/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI1/MM7 N_XI0/XI0/XI1/NET36_XI0/XI0/XI1/MM7_d
+ N_XI0/XI0/XI1/NET35_XI0/XI0/XI1/MM7_g N_VSS_XI0/XI0/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI1/MM8 N_XI0/XI0/XI1/NET35_XI0/XI0/XI1/MM8_d N_WL<1>_XI0/XI0/XI1/MM8_g
+ N_BLN<14>_XI0/XI0/XI1/MM8_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI1/MM5 N_XI0/XI0/XI1/NET34_XI0/XI0/XI1/MM5_d
+ N_XI0/XI0/XI1/NET33_XI0/XI0/XI1/MM5_g N_VDD_XI0/XI0/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI1/MM4 N_XI0/XI0/XI1/NET33_XI0/XI0/XI1/MM4_d
+ N_XI0/XI0/XI1/NET34_XI0/XI0/XI1/MM4_g N_VDD_XI0/XI0/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI1/MM10 N_XI0/XI0/XI1/NET35_XI0/XI0/XI1/MM10_d
+ N_XI0/XI0/XI1/NET36_XI0/XI0/XI1/MM10_g N_VDD_XI0/XI0/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI1/MM11 N_XI0/XI0/XI1/NET36_XI0/XI0/XI1/MM11_d
+ N_XI0/XI0/XI1/NET35_XI0/XI0/XI1/MM11_g N_VDD_XI0/XI0/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI2/MM2 N_XI0/XI0/XI2/NET34_XI0/XI0/XI2/MM2_d
+ N_XI0/XI0/XI2/NET33_XI0/XI0/XI2/MM2_g N_VSS_XI0/XI0/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI2/MM3 N_XI0/XI0/XI2/NET33_XI0/XI0/XI2/MM3_d N_WL<0>_XI0/XI0/XI2/MM3_g
+ N_BLN<13>_XI0/XI0/XI2/MM3_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI2/MM0 N_XI0/XI0/XI2/NET34_XI0/XI0/XI2/MM0_d N_WL<0>_XI0/XI0/XI2/MM0_g
+ N_BL<13>_XI0/XI0/XI2/MM0_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI2/MM1 N_XI0/XI0/XI2/NET33_XI0/XI0/XI2/MM1_d
+ N_XI0/XI0/XI2/NET34_XI0/XI0/XI2/MM1_g N_VSS_XI0/XI0/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI2/MM9 N_XI0/XI0/XI2/NET36_XI0/XI0/XI2/MM9_d N_WL<1>_XI0/XI0/XI2/MM9_g
+ N_BL<13>_XI0/XI0/XI2/MM9_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI2/MM6 N_XI0/XI0/XI2/NET35_XI0/XI0/XI2/MM6_d
+ N_XI0/XI0/XI2/NET36_XI0/XI0/XI2/MM6_g N_VSS_XI0/XI0/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI2/MM7 N_XI0/XI0/XI2/NET36_XI0/XI0/XI2/MM7_d
+ N_XI0/XI0/XI2/NET35_XI0/XI0/XI2/MM7_g N_VSS_XI0/XI0/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI2/MM8 N_XI0/XI0/XI2/NET35_XI0/XI0/XI2/MM8_d N_WL<1>_XI0/XI0/XI2/MM8_g
+ N_BLN<13>_XI0/XI0/XI2/MM8_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI2/MM5 N_XI0/XI0/XI2/NET34_XI0/XI0/XI2/MM5_d
+ N_XI0/XI0/XI2/NET33_XI0/XI0/XI2/MM5_g N_VDD_XI0/XI0/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI2/MM4 N_XI0/XI0/XI2/NET33_XI0/XI0/XI2/MM4_d
+ N_XI0/XI0/XI2/NET34_XI0/XI0/XI2/MM4_g N_VDD_XI0/XI0/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI2/MM10 N_XI0/XI0/XI2/NET35_XI0/XI0/XI2/MM10_d
+ N_XI0/XI0/XI2/NET36_XI0/XI0/XI2/MM10_g N_VDD_XI0/XI0/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI2/MM11 N_XI0/XI0/XI2/NET36_XI0/XI0/XI2/MM11_d
+ N_XI0/XI0/XI2/NET35_XI0/XI0/XI2/MM11_g N_VDD_XI0/XI0/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI3/MM2 N_XI0/XI0/XI3/NET34_XI0/XI0/XI3/MM2_d
+ N_XI0/XI0/XI3/NET33_XI0/XI0/XI3/MM2_g N_VSS_XI0/XI0/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI3/MM3 N_XI0/XI0/XI3/NET33_XI0/XI0/XI3/MM3_d N_WL<0>_XI0/XI0/XI3/MM3_g
+ N_BLN<12>_XI0/XI0/XI3/MM3_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI3/MM0 N_XI0/XI0/XI3/NET34_XI0/XI0/XI3/MM0_d N_WL<0>_XI0/XI0/XI3/MM0_g
+ N_BL<12>_XI0/XI0/XI3/MM0_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI3/MM1 N_XI0/XI0/XI3/NET33_XI0/XI0/XI3/MM1_d
+ N_XI0/XI0/XI3/NET34_XI0/XI0/XI3/MM1_g N_VSS_XI0/XI0/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI3/MM9 N_XI0/XI0/XI3/NET36_XI0/XI0/XI3/MM9_d N_WL<1>_XI0/XI0/XI3/MM9_g
+ N_BL<12>_XI0/XI0/XI3/MM9_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI3/MM6 N_XI0/XI0/XI3/NET35_XI0/XI0/XI3/MM6_d
+ N_XI0/XI0/XI3/NET36_XI0/XI0/XI3/MM6_g N_VSS_XI0/XI0/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI3/MM7 N_XI0/XI0/XI3/NET36_XI0/XI0/XI3/MM7_d
+ N_XI0/XI0/XI3/NET35_XI0/XI0/XI3/MM7_g N_VSS_XI0/XI0/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI3/MM8 N_XI0/XI0/XI3/NET35_XI0/XI0/XI3/MM8_d N_WL<1>_XI0/XI0/XI3/MM8_g
+ N_BLN<12>_XI0/XI0/XI3/MM8_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI3/MM5 N_XI0/XI0/XI3/NET34_XI0/XI0/XI3/MM5_d
+ N_XI0/XI0/XI3/NET33_XI0/XI0/XI3/MM5_g N_VDD_XI0/XI0/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI3/MM4 N_XI0/XI0/XI3/NET33_XI0/XI0/XI3/MM4_d
+ N_XI0/XI0/XI3/NET34_XI0/XI0/XI3/MM4_g N_VDD_XI0/XI0/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI3/MM10 N_XI0/XI0/XI3/NET35_XI0/XI0/XI3/MM10_d
+ N_XI0/XI0/XI3/NET36_XI0/XI0/XI3/MM10_g N_VDD_XI0/XI0/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI3/MM11 N_XI0/XI0/XI3/NET36_XI0/XI0/XI3/MM11_d
+ N_XI0/XI0/XI3/NET35_XI0/XI0/XI3/MM11_g N_VDD_XI0/XI0/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI4/MM2 N_XI0/XI0/XI4/NET34_XI0/XI0/XI4/MM2_d
+ N_XI0/XI0/XI4/NET33_XI0/XI0/XI4/MM2_g N_VSS_XI0/XI0/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI4/MM3 N_XI0/XI0/XI4/NET33_XI0/XI0/XI4/MM3_d N_WL<0>_XI0/XI0/XI4/MM3_g
+ N_BLN<11>_XI0/XI0/XI4/MM3_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI4/MM0 N_XI0/XI0/XI4/NET34_XI0/XI0/XI4/MM0_d N_WL<0>_XI0/XI0/XI4/MM0_g
+ N_BL<11>_XI0/XI0/XI4/MM0_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI4/MM1 N_XI0/XI0/XI4/NET33_XI0/XI0/XI4/MM1_d
+ N_XI0/XI0/XI4/NET34_XI0/XI0/XI4/MM1_g N_VSS_XI0/XI0/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI4/MM9 N_XI0/XI0/XI4/NET36_XI0/XI0/XI4/MM9_d N_WL<1>_XI0/XI0/XI4/MM9_g
+ N_BL<11>_XI0/XI0/XI4/MM9_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI4/MM6 N_XI0/XI0/XI4/NET35_XI0/XI0/XI4/MM6_d
+ N_XI0/XI0/XI4/NET36_XI0/XI0/XI4/MM6_g N_VSS_XI0/XI0/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI4/MM7 N_XI0/XI0/XI4/NET36_XI0/XI0/XI4/MM7_d
+ N_XI0/XI0/XI4/NET35_XI0/XI0/XI4/MM7_g N_VSS_XI0/XI0/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI4/MM8 N_XI0/XI0/XI4/NET35_XI0/XI0/XI4/MM8_d N_WL<1>_XI0/XI0/XI4/MM8_g
+ N_BLN<11>_XI0/XI0/XI4/MM8_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI4/MM5 N_XI0/XI0/XI4/NET34_XI0/XI0/XI4/MM5_d
+ N_XI0/XI0/XI4/NET33_XI0/XI0/XI4/MM5_g N_VDD_XI0/XI0/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI4/MM4 N_XI0/XI0/XI4/NET33_XI0/XI0/XI4/MM4_d
+ N_XI0/XI0/XI4/NET34_XI0/XI0/XI4/MM4_g N_VDD_XI0/XI0/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI4/MM10 N_XI0/XI0/XI4/NET35_XI0/XI0/XI4/MM10_d
+ N_XI0/XI0/XI4/NET36_XI0/XI0/XI4/MM10_g N_VDD_XI0/XI0/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI4/MM11 N_XI0/XI0/XI4/NET36_XI0/XI0/XI4/MM11_d
+ N_XI0/XI0/XI4/NET35_XI0/XI0/XI4/MM11_g N_VDD_XI0/XI0/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI5/MM2 N_XI0/XI0/XI5/NET34_XI0/XI0/XI5/MM2_d
+ N_XI0/XI0/XI5/NET33_XI0/XI0/XI5/MM2_g N_VSS_XI0/XI0/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI5/MM3 N_XI0/XI0/XI5/NET33_XI0/XI0/XI5/MM3_d N_WL<0>_XI0/XI0/XI5/MM3_g
+ N_BLN<10>_XI0/XI0/XI5/MM3_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI5/MM0 N_XI0/XI0/XI5/NET34_XI0/XI0/XI5/MM0_d N_WL<0>_XI0/XI0/XI5/MM0_g
+ N_BL<10>_XI0/XI0/XI5/MM0_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI5/MM1 N_XI0/XI0/XI5/NET33_XI0/XI0/XI5/MM1_d
+ N_XI0/XI0/XI5/NET34_XI0/XI0/XI5/MM1_g N_VSS_XI0/XI0/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI5/MM9 N_XI0/XI0/XI5/NET36_XI0/XI0/XI5/MM9_d N_WL<1>_XI0/XI0/XI5/MM9_g
+ N_BL<10>_XI0/XI0/XI5/MM9_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI5/MM6 N_XI0/XI0/XI5/NET35_XI0/XI0/XI5/MM6_d
+ N_XI0/XI0/XI5/NET36_XI0/XI0/XI5/MM6_g N_VSS_XI0/XI0/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI5/MM7 N_XI0/XI0/XI5/NET36_XI0/XI0/XI5/MM7_d
+ N_XI0/XI0/XI5/NET35_XI0/XI0/XI5/MM7_g N_VSS_XI0/XI0/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI5/MM8 N_XI0/XI0/XI5/NET35_XI0/XI0/XI5/MM8_d N_WL<1>_XI0/XI0/XI5/MM8_g
+ N_BLN<10>_XI0/XI0/XI5/MM8_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI5/MM5 N_XI0/XI0/XI5/NET34_XI0/XI0/XI5/MM5_d
+ N_XI0/XI0/XI5/NET33_XI0/XI0/XI5/MM5_g N_VDD_XI0/XI0/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI5/MM4 N_XI0/XI0/XI5/NET33_XI0/XI0/XI5/MM4_d
+ N_XI0/XI0/XI5/NET34_XI0/XI0/XI5/MM4_g N_VDD_XI0/XI0/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI5/MM10 N_XI0/XI0/XI5/NET35_XI0/XI0/XI5/MM10_d
+ N_XI0/XI0/XI5/NET36_XI0/XI0/XI5/MM10_g N_VDD_XI0/XI0/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI5/MM11 N_XI0/XI0/XI5/NET36_XI0/XI0/XI5/MM11_d
+ N_XI0/XI0/XI5/NET35_XI0/XI0/XI5/MM11_g N_VDD_XI0/XI0/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI6/MM2 N_XI0/XI0/XI6/NET34_XI0/XI0/XI6/MM2_d
+ N_XI0/XI0/XI6/NET33_XI0/XI0/XI6/MM2_g N_VSS_XI0/XI0/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI6/MM3 N_XI0/XI0/XI6/NET33_XI0/XI0/XI6/MM3_d N_WL<0>_XI0/XI0/XI6/MM3_g
+ N_BLN<9>_XI0/XI0/XI6/MM3_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI6/MM0 N_XI0/XI0/XI6/NET34_XI0/XI0/XI6/MM0_d N_WL<0>_XI0/XI0/XI6/MM0_g
+ N_BL<9>_XI0/XI0/XI6/MM0_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI6/MM1 N_XI0/XI0/XI6/NET33_XI0/XI0/XI6/MM1_d
+ N_XI0/XI0/XI6/NET34_XI0/XI0/XI6/MM1_g N_VSS_XI0/XI0/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI6/MM9 N_XI0/XI0/XI6/NET36_XI0/XI0/XI6/MM9_d N_WL<1>_XI0/XI0/XI6/MM9_g
+ N_BL<9>_XI0/XI0/XI6/MM9_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI6/MM6 N_XI0/XI0/XI6/NET35_XI0/XI0/XI6/MM6_d
+ N_XI0/XI0/XI6/NET36_XI0/XI0/XI6/MM6_g N_VSS_XI0/XI0/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI6/MM7 N_XI0/XI0/XI6/NET36_XI0/XI0/XI6/MM7_d
+ N_XI0/XI0/XI6/NET35_XI0/XI0/XI6/MM7_g N_VSS_XI0/XI0/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI6/MM8 N_XI0/XI0/XI6/NET35_XI0/XI0/XI6/MM8_d N_WL<1>_XI0/XI0/XI6/MM8_g
+ N_BLN<9>_XI0/XI0/XI6/MM8_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI6/MM5 N_XI0/XI0/XI6/NET34_XI0/XI0/XI6/MM5_d
+ N_XI0/XI0/XI6/NET33_XI0/XI0/XI6/MM5_g N_VDD_XI0/XI0/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI6/MM4 N_XI0/XI0/XI6/NET33_XI0/XI0/XI6/MM4_d
+ N_XI0/XI0/XI6/NET34_XI0/XI0/XI6/MM4_g N_VDD_XI0/XI0/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI6/MM10 N_XI0/XI0/XI6/NET35_XI0/XI0/XI6/MM10_d
+ N_XI0/XI0/XI6/NET36_XI0/XI0/XI6/MM10_g N_VDD_XI0/XI0/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI6/MM11 N_XI0/XI0/XI6/NET36_XI0/XI0/XI6/MM11_d
+ N_XI0/XI0/XI6/NET35_XI0/XI0/XI6/MM11_g N_VDD_XI0/XI0/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI7/MM2 N_XI0/XI0/XI7/NET34_XI0/XI0/XI7/MM2_d
+ N_XI0/XI0/XI7/NET33_XI0/XI0/XI7/MM2_g N_VSS_XI0/XI0/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI7/MM3 N_XI0/XI0/XI7/NET33_XI0/XI0/XI7/MM3_d N_WL<0>_XI0/XI0/XI7/MM3_g
+ N_BLN<8>_XI0/XI0/XI7/MM3_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI7/MM0 N_XI0/XI0/XI7/NET34_XI0/XI0/XI7/MM0_d N_WL<0>_XI0/XI0/XI7/MM0_g
+ N_BL<8>_XI0/XI0/XI7/MM0_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI7/MM1 N_XI0/XI0/XI7/NET33_XI0/XI0/XI7/MM1_d
+ N_XI0/XI0/XI7/NET34_XI0/XI0/XI7/MM1_g N_VSS_XI0/XI0/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI7/MM9 N_XI0/XI0/XI7/NET36_XI0/XI0/XI7/MM9_d N_WL<1>_XI0/XI0/XI7/MM9_g
+ N_BL<8>_XI0/XI0/XI7/MM9_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI7/MM6 N_XI0/XI0/XI7/NET35_XI0/XI0/XI7/MM6_d
+ N_XI0/XI0/XI7/NET36_XI0/XI0/XI7/MM6_g N_VSS_XI0/XI0/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI7/MM7 N_XI0/XI0/XI7/NET36_XI0/XI0/XI7/MM7_d
+ N_XI0/XI0/XI7/NET35_XI0/XI0/XI7/MM7_g N_VSS_XI0/XI0/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI7/MM8 N_XI0/XI0/XI7/NET35_XI0/XI0/XI7/MM8_d N_WL<1>_XI0/XI0/XI7/MM8_g
+ N_BLN<8>_XI0/XI0/XI7/MM8_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI7/MM5 N_XI0/XI0/XI7/NET34_XI0/XI0/XI7/MM5_d
+ N_XI0/XI0/XI7/NET33_XI0/XI0/XI7/MM5_g N_VDD_XI0/XI0/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI7/MM4 N_XI0/XI0/XI7/NET33_XI0/XI0/XI7/MM4_d
+ N_XI0/XI0/XI7/NET34_XI0/XI0/XI7/MM4_g N_VDD_XI0/XI0/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI7/MM10 N_XI0/XI0/XI7/NET35_XI0/XI0/XI7/MM10_d
+ N_XI0/XI0/XI7/NET36_XI0/XI0/XI7/MM10_g N_VDD_XI0/XI0/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI7/MM11 N_XI0/XI0/XI7/NET36_XI0/XI0/XI7/MM11_d
+ N_XI0/XI0/XI7/NET35_XI0/XI0/XI7/MM11_g N_VDD_XI0/XI0/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI8/MM2 N_XI0/XI0/XI8/NET34_XI0/XI0/XI8/MM2_d
+ N_XI0/XI0/XI8/NET33_XI0/XI0/XI8/MM2_g N_VSS_XI0/XI0/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI8/MM3 N_XI0/XI0/XI8/NET33_XI0/XI0/XI8/MM3_d N_WL<0>_XI0/XI0/XI8/MM3_g
+ N_BLN<7>_XI0/XI0/XI8/MM3_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI8/MM0 N_XI0/XI0/XI8/NET34_XI0/XI0/XI8/MM0_d N_WL<0>_XI0/XI0/XI8/MM0_g
+ N_BL<7>_XI0/XI0/XI8/MM0_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI8/MM1 N_XI0/XI0/XI8/NET33_XI0/XI0/XI8/MM1_d
+ N_XI0/XI0/XI8/NET34_XI0/XI0/XI8/MM1_g N_VSS_XI0/XI0/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI8/MM9 N_XI0/XI0/XI8/NET36_XI0/XI0/XI8/MM9_d N_WL<1>_XI0/XI0/XI8/MM9_g
+ N_BL<7>_XI0/XI0/XI8/MM9_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI8/MM6 N_XI0/XI0/XI8/NET35_XI0/XI0/XI8/MM6_d
+ N_XI0/XI0/XI8/NET36_XI0/XI0/XI8/MM6_g N_VSS_XI0/XI0/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI8/MM7 N_XI0/XI0/XI8/NET36_XI0/XI0/XI8/MM7_d
+ N_XI0/XI0/XI8/NET35_XI0/XI0/XI8/MM7_g N_VSS_XI0/XI0/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI8/MM8 N_XI0/XI0/XI8/NET35_XI0/XI0/XI8/MM8_d N_WL<1>_XI0/XI0/XI8/MM8_g
+ N_BLN<7>_XI0/XI0/XI8/MM8_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI8/MM5 N_XI0/XI0/XI8/NET34_XI0/XI0/XI8/MM5_d
+ N_XI0/XI0/XI8/NET33_XI0/XI0/XI8/MM5_g N_VDD_XI0/XI0/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI8/MM4 N_XI0/XI0/XI8/NET33_XI0/XI0/XI8/MM4_d
+ N_XI0/XI0/XI8/NET34_XI0/XI0/XI8/MM4_g N_VDD_XI0/XI0/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI8/MM10 N_XI0/XI0/XI8/NET35_XI0/XI0/XI8/MM10_d
+ N_XI0/XI0/XI8/NET36_XI0/XI0/XI8/MM10_g N_VDD_XI0/XI0/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI8/MM11 N_XI0/XI0/XI8/NET36_XI0/XI0/XI8/MM11_d
+ N_XI0/XI0/XI8/NET35_XI0/XI0/XI8/MM11_g N_VDD_XI0/XI0/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI9/MM2 N_XI0/XI0/XI9/NET34_XI0/XI0/XI9/MM2_d
+ N_XI0/XI0/XI9/NET33_XI0/XI0/XI9/MM2_g N_VSS_XI0/XI0/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI9/MM3 N_XI0/XI0/XI9/NET33_XI0/XI0/XI9/MM3_d N_WL<0>_XI0/XI0/XI9/MM3_g
+ N_BLN<6>_XI0/XI0/XI9/MM3_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI9/MM0 N_XI0/XI0/XI9/NET34_XI0/XI0/XI9/MM0_d N_WL<0>_XI0/XI0/XI9/MM0_g
+ N_BL<6>_XI0/XI0/XI9/MM0_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI9/MM1 N_XI0/XI0/XI9/NET33_XI0/XI0/XI9/MM1_d
+ N_XI0/XI0/XI9/NET34_XI0/XI0/XI9/MM1_g N_VSS_XI0/XI0/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI9/MM9 N_XI0/XI0/XI9/NET36_XI0/XI0/XI9/MM9_d N_WL<1>_XI0/XI0/XI9/MM9_g
+ N_BL<6>_XI0/XI0/XI9/MM9_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI9/MM6 N_XI0/XI0/XI9/NET35_XI0/XI0/XI9/MM6_d
+ N_XI0/XI0/XI9/NET36_XI0/XI0/XI9/MM6_g N_VSS_XI0/XI0/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI9/MM7 N_XI0/XI0/XI9/NET36_XI0/XI0/XI9/MM7_d
+ N_XI0/XI0/XI9/NET35_XI0/XI0/XI9/MM7_g N_VSS_XI0/XI0/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI9/MM8 N_XI0/XI0/XI9/NET35_XI0/XI0/XI9/MM8_d N_WL<1>_XI0/XI0/XI9/MM8_g
+ N_BLN<6>_XI0/XI0/XI9/MM8_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI0/XI9/MM5 N_XI0/XI0/XI9/NET34_XI0/XI0/XI9/MM5_d
+ N_XI0/XI0/XI9/NET33_XI0/XI0/XI9/MM5_g N_VDD_XI0/XI0/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI9/MM4 N_XI0/XI0/XI9/NET33_XI0/XI0/XI9/MM4_d
+ N_XI0/XI0/XI9/NET34_XI0/XI0/XI9/MM4_g N_VDD_XI0/XI0/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI9/MM10 N_XI0/XI0/XI9/NET35_XI0/XI0/XI9/MM10_d
+ N_XI0/XI0/XI9/NET36_XI0/XI0/XI9/MM10_g N_VDD_XI0/XI0/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI9/MM11 N_XI0/XI0/XI9/NET36_XI0/XI0/XI9/MM11_d
+ N_XI0/XI0/XI9/NET35_XI0/XI0/XI9/MM11_g N_VDD_XI0/XI0/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI10/MM2 N_XI0/XI0/XI10/NET34_XI0/XI0/XI10/MM2_d
+ N_XI0/XI0/XI10/NET33_XI0/XI0/XI10/MM2_g N_VSS_XI0/XI0/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM3 N_XI0/XI0/XI10/NET33_XI0/XI0/XI10/MM3_d
+ N_WL<0>_XI0/XI0/XI10/MM3_g N_BLN<5>_XI0/XI0/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM0 N_XI0/XI0/XI10/NET34_XI0/XI0/XI10/MM0_d
+ N_WL<0>_XI0/XI0/XI10/MM0_g N_BL<5>_XI0/XI0/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM1 N_XI0/XI0/XI10/NET33_XI0/XI0/XI10/MM1_d
+ N_XI0/XI0/XI10/NET34_XI0/XI0/XI10/MM1_g N_VSS_XI0/XI0/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM9 N_XI0/XI0/XI10/NET36_XI0/XI0/XI10/MM9_d
+ N_WL<1>_XI0/XI0/XI10/MM9_g N_BL<5>_XI0/XI0/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM6 N_XI0/XI0/XI10/NET35_XI0/XI0/XI10/MM6_d
+ N_XI0/XI0/XI10/NET36_XI0/XI0/XI10/MM6_g N_VSS_XI0/XI0/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM7 N_XI0/XI0/XI10/NET36_XI0/XI0/XI10/MM7_d
+ N_XI0/XI0/XI10/NET35_XI0/XI0/XI10/MM7_g N_VSS_XI0/XI0/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM8 N_XI0/XI0/XI10/NET35_XI0/XI0/XI10/MM8_d
+ N_WL<1>_XI0/XI0/XI10/MM8_g N_BLN<5>_XI0/XI0/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI10/MM5 N_XI0/XI0/XI10/NET34_XI0/XI0/XI10/MM5_d
+ N_XI0/XI0/XI10/NET33_XI0/XI0/XI10/MM5_g N_VDD_XI0/XI0/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI10/MM4 N_XI0/XI0/XI10/NET33_XI0/XI0/XI10/MM4_d
+ N_XI0/XI0/XI10/NET34_XI0/XI0/XI10/MM4_g N_VDD_XI0/XI0/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI10/MM10 N_XI0/XI0/XI10/NET35_XI0/XI0/XI10/MM10_d
+ N_XI0/XI0/XI10/NET36_XI0/XI0/XI10/MM10_g N_VDD_XI0/XI0/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI10/MM11 N_XI0/XI0/XI10/NET36_XI0/XI0/XI10/MM11_d
+ N_XI0/XI0/XI10/NET35_XI0/XI0/XI10/MM11_g N_VDD_XI0/XI0/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI11/MM2 N_XI0/XI0/XI11/NET34_XI0/XI0/XI11/MM2_d
+ N_XI0/XI0/XI11/NET33_XI0/XI0/XI11/MM2_g N_VSS_XI0/XI0/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM3 N_XI0/XI0/XI11/NET33_XI0/XI0/XI11/MM3_d
+ N_WL<0>_XI0/XI0/XI11/MM3_g N_BLN<4>_XI0/XI0/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM0 N_XI0/XI0/XI11/NET34_XI0/XI0/XI11/MM0_d
+ N_WL<0>_XI0/XI0/XI11/MM0_g N_BL<4>_XI0/XI0/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM1 N_XI0/XI0/XI11/NET33_XI0/XI0/XI11/MM1_d
+ N_XI0/XI0/XI11/NET34_XI0/XI0/XI11/MM1_g N_VSS_XI0/XI0/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM9 N_XI0/XI0/XI11/NET36_XI0/XI0/XI11/MM9_d
+ N_WL<1>_XI0/XI0/XI11/MM9_g N_BL<4>_XI0/XI0/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM6 N_XI0/XI0/XI11/NET35_XI0/XI0/XI11/MM6_d
+ N_XI0/XI0/XI11/NET36_XI0/XI0/XI11/MM6_g N_VSS_XI0/XI0/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM7 N_XI0/XI0/XI11/NET36_XI0/XI0/XI11/MM7_d
+ N_XI0/XI0/XI11/NET35_XI0/XI0/XI11/MM7_g N_VSS_XI0/XI0/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM8 N_XI0/XI0/XI11/NET35_XI0/XI0/XI11/MM8_d
+ N_WL<1>_XI0/XI0/XI11/MM8_g N_BLN<4>_XI0/XI0/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI11/MM5 N_XI0/XI0/XI11/NET34_XI0/XI0/XI11/MM5_d
+ N_XI0/XI0/XI11/NET33_XI0/XI0/XI11/MM5_g N_VDD_XI0/XI0/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI11/MM4 N_XI0/XI0/XI11/NET33_XI0/XI0/XI11/MM4_d
+ N_XI0/XI0/XI11/NET34_XI0/XI0/XI11/MM4_g N_VDD_XI0/XI0/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI11/MM10 N_XI0/XI0/XI11/NET35_XI0/XI0/XI11/MM10_d
+ N_XI0/XI0/XI11/NET36_XI0/XI0/XI11/MM10_g N_VDD_XI0/XI0/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI11/MM11 N_XI0/XI0/XI11/NET36_XI0/XI0/XI11/MM11_d
+ N_XI0/XI0/XI11/NET35_XI0/XI0/XI11/MM11_g N_VDD_XI0/XI0/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI12/MM2 N_XI0/XI0/XI12/NET34_XI0/XI0/XI12/MM2_d
+ N_XI0/XI0/XI12/NET33_XI0/XI0/XI12/MM2_g N_VSS_XI0/XI0/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM3 N_XI0/XI0/XI12/NET33_XI0/XI0/XI12/MM3_d
+ N_WL<0>_XI0/XI0/XI12/MM3_g N_BLN<3>_XI0/XI0/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM0 N_XI0/XI0/XI12/NET34_XI0/XI0/XI12/MM0_d
+ N_WL<0>_XI0/XI0/XI12/MM0_g N_BL<3>_XI0/XI0/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM1 N_XI0/XI0/XI12/NET33_XI0/XI0/XI12/MM1_d
+ N_XI0/XI0/XI12/NET34_XI0/XI0/XI12/MM1_g N_VSS_XI0/XI0/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM9 N_XI0/XI0/XI12/NET36_XI0/XI0/XI12/MM9_d
+ N_WL<1>_XI0/XI0/XI12/MM9_g N_BL<3>_XI0/XI0/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM6 N_XI0/XI0/XI12/NET35_XI0/XI0/XI12/MM6_d
+ N_XI0/XI0/XI12/NET36_XI0/XI0/XI12/MM6_g N_VSS_XI0/XI0/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM7 N_XI0/XI0/XI12/NET36_XI0/XI0/XI12/MM7_d
+ N_XI0/XI0/XI12/NET35_XI0/XI0/XI12/MM7_g N_VSS_XI0/XI0/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM8 N_XI0/XI0/XI12/NET35_XI0/XI0/XI12/MM8_d
+ N_WL<1>_XI0/XI0/XI12/MM8_g N_BLN<3>_XI0/XI0/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI12/MM5 N_XI0/XI0/XI12/NET34_XI0/XI0/XI12/MM5_d
+ N_XI0/XI0/XI12/NET33_XI0/XI0/XI12/MM5_g N_VDD_XI0/XI0/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI12/MM4 N_XI0/XI0/XI12/NET33_XI0/XI0/XI12/MM4_d
+ N_XI0/XI0/XI12/NET34_XI0/XI0/XI12/MM4_g N_VDD_XI0/XI0/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI12/MM10 N_XI0/XI0/XI12/NET35_XI0/XI0/XI12/MM10_d
+ N_XI0/XI0/XI12/NET36_XI0/XI0/XI12/MM10_g N_VDD_XI0/XI0/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI12/MM11 N_XI0/XI0/XI12/NET36_XI0/XI0/XI12/MM11_d
+ N_XI0/XI0/XI12/NET35_XI0/XI0/XI12/MM11_g N_VDD_XI0/XI0/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI13/MM2 N_XI0/XI0/XI13/NET34_XI0/XI0/XI13/MM2_d
+ N_XI0/XI0/XI13/NET33_XI0/XI0/XI13/MM2_g N_VSS_XI0/XI0/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM3 N_XI0/XI0/XI13/NET33_XI0/XI0/XI13/MM3_d
+ N_WL<0>_XI0/XI0/XI13/MM3_g N_BLN<2>_XI0/XI0/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM0 N_XI0/XI0/XI13/NET34_XI0/XI0/XI13/MM0_d
+ N_WL<0>_XI0/XI0/XI13/MM0_g N_BL<2>_XI0/XI0/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM1 N_XI0/XI0/XI13/NET33_XI0/XI0/XI13/MM1_d
+ N_XI0/XI0/XI13/NET34_XI0/XI0/XI13/MM1_g N_VSS_XI0/XI0/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM9 N_XI0/XI0/XI13/NET36_XI0/XI0/XI13/MM9_d
+ N_WL<1>_XI0/XI0/XI13/MM9_g N_BL<2>_XI0/XI0/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM6 N_XI0/XI0/XI13/NET35_XI0/XI0/XI13/MM6_d
+ N_XI0/XI0/XI13/NET36_XI0/XI0/XI13/MM6_g N_VSS_XI0/XI0/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM7 N_XI0/XI0/XI13/NET36_XI0/XI0/XI13/MM7_d
+ N_XI0/XI0/XI13/NET35_XI0/XI0/XI13/MM7_g N_VSS_XI0/XI0/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM8 N_XI0/XI0/XI13/NET35_XI0/XI0/XI13/MM8_d
+ N_WL<1>_XI0/XI0/XI13/MM8_g N_BLN<2>_XI0/XI0/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI13/MM5 N_XI0/XI0/XI13/NET34_XI0/XI0/XI13/MM5_d
+ N_XI0/XI0/XI13/NET33_XI0/XI0/XI13/MM5_g N_VDD_XI0/XI0/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI13/MM4 N_XI0/XI0/XI13/NET33_XI0/XI0/XI13/MM4_d
+ N_XI0/XI0/XI13/NET34_XI0/XI0/XI13/MM4_g N_VDD_XI0/XI0/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI13/MM10 N_XI0/XI0/XI13/NET35_XI0/XI0/XI13/MM10_d
+ N_XI0/XI0/XI13/NET36_XI0/XI0/XI13/MM10_g N_VDD_XI0/XI0/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI13/MM11 N_XI0/XI0/XI13/NET36_XI0/XI0/XI13/MM11_d
+ N_XI0/XI0/XI13/NET35_XI0/XI0/XI13/MM11_g N_VDD_XI0/XI0/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI14/MM2 N_XI0/XI0/XI14/NET34_XI0/XI0/XI14/MM2_d
+ N_XI0/XI0/XI14/NET33_XI0/XI0/XI14/MM2_g N_VSS_XI0/XI0/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM3 N_XI0/XI0/XI14/NET33_XI0/XI0/XI14/MM3_d
+ N_WL<0>_XI0/XI0/XI14/MM3_g N_BLN<1>_XI0/XI0/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM0 N_XI0/XI0/XI14/NET34_XI0/XI0/XI14/MM0_d
+ N_WL<0>_XI0/XI0/XI14/MM0_g N_BL<1>_XI0/XI0/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM1 N_XI0/XI0/XI14/NET33_XI0/XI0/XI14/MM1_d
+ N_XI0/XI0/XI14/NET34_XI0/XI0/XI14/MM1_g N_VSS_XI0/XI0/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM9 N_XI0/XI0/XI14/NET36_XI0/XI0/XI14/MM9_d
+ N_WL<1>_XI0/XI0/XI14/MM9_g N_BL<1>_XI0/XI0/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM6 N_XI0/XI0/XI14/NET35_XI0/XI0/XI14/MM6_d
+ N_XI0/XI0/XI14/NET36_XI0/XI0/XI14/MM6_g N_VSS_XI0/XI0/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM7 N_XI0/XI0/XI14/NET36_XI0/XI0/XI14/MM7_d
+ N_XI0/XI0/XI14/NET35_XI0/XI0/XI14/MM7_g N_VSS_XI0/XI0/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM8 N_XI0/XI0/XI14/NET35_XI0/XI0/XI14/MM8_d
+ N_WL<1>_XI0/XI0/XI14/MM8_g N_BLN<1>_XI0/XI0/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI14/MM5 N_XI0/XI0/XI14/NET34_XI0/XI0/XI14/MM5_d
+ N_XI0/XI0/XI14/NET33_XI0/XI0/XI14/MM5_g N_VDD_XI0/XI0/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI14/MM4 N_XI0/XI0/XI14/NET33_XI0/XI0/XI14/MM4_d
+ N_XI0/XI0/XI14/NET34_XI0/XI0/XI14/MM4_g N_VDD_XI0/XI0/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI14/MM10 N_XI0/XI0/XI14/NET35_XI0/XI0/XI14/MM10_d
+ N_XI0/XI0/XI14/NET36_XI0/XI0/XI14/MM10_g N_VDD_XI0/XI0/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI14/MM11 N_XI0/XI0/XI14/NET36_XI0/XI0/XI14/MM11_d
+ N_XI0/XI0/XI14/NET35_XI0/XI0/XI14/MM11_g N_VDD_XI0/XI0/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI15/MM2 N_XI0/XI0/XI15/NET34_XI0/XI0/XI15/MM2_d
+ N_XI0/XI0/XI15/NET33_XI0/XI0/XI15/MM2_g N_VSS_XI0/XI0/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM3 N_XI0/XI0/XI15/NET33_XI0/XI0/XI15/MM3_d
+ N_WL<0>_XI0/XI0/XI15/MM3_g N_BLN<0>_XI0/XI0/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM0 N_XI0/XI0/XI15/NET34_XI0/XI0/XI15/MM0_d
+ N_WL<0>_XI0/XI0/XI15/MM0_g N_BL<0>_XI0/XI0/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM1 N_XI0/XI0/XI15/NET33_XI0/XI0/XI15/MM1_d
+ N_XI0/XI0/XI15/NET34_XI0/XI0/XI15/MM1_g N_VSS_XI0/XI0/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM9 N_XI0/XI0/XI15/NET36_XI0/XI0/XI15/MM9_d
+ N_WL<1>_XI0/XI0/XI15/MM9_g N_BL<0>_XI0/XI0/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM6 N_XI0/XI0/XI15/NET35_XI0/XI0/XI15/MM6_d
+ N_XI0/XI0/XI15/NET36_XI0/XI0/XI15/MM6_g N_VSS_XI0/XI0/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM7 N_XI0/XI0/XI15/NET36_XI0/XI0/XI15/MM7_d
+ N_XI0/XI0/XI15/NET35_XI0/XI0/XI15/MM7_g N_VSS_XI0/XI0/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM8 N_XI0/XI0/XI15/NET35_XI0/XI0/XI15/MM8_d
+ N_WL<1>_XI0/XI0/XI15/MM8_g N_BLN<0>_XI0/XI0/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/XI15/MM5 N_XI0/XI0/XI15/NET34_XI0/XI0/XI15/MM5_d
+ N_XI0/XI0/XI15/NET33_XI0/XI0/XI15/MM5_g N_VDD_XI0/XI0/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI15/MM4 N_XI0/XI0/XI15/NET33_XI0/XI0/XI15/MM4_d
+ N_XI0/XI0/XI15/NET34_XI0/XI0/XI15/MM4_g N_VDD_XI0/XI0/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI15/MM10 N_XI0/XI0/XI15/NET35_XI0/XI0/XI15/MM10_d
+ N_XI0/XI0/XI15/NET36_XI0/XI0/XI15/MM10_g N_VDD_XI0/XI0/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/XI15/MM11 N_XI0/XI0/XI15/NET36_XI0/XI0/XI15/MM11_d
+ N_XI0/XI0/XI15/NET35_XI0/XI0/XI15/MM11_g N_VDD_XI0/XI0/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI0/MM2 N_XI0/XI1/XI0/NET34_XI0/XI1/XI0/MM2_d
+ N_XI0/XI1/XI0/NET33_XI0/XI1/XI0/MM2_g N_VSS_XI0/XI1/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI0/MM3 N_XI0/XI1/XI0/NET33_XI0/XI1/XI0/MM3_d N_WL<2>_XI0/XI1/XI0/MM3_g
+ N_BLN<15>_XI0/XI1/XI0/MM3_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI0/MM0 N_XI0/XI1/XI0/NET34_XI0/XI1/XI0/MM0_d N_WL<2>_XI0/XI1/XI0/MM0_g
+ N_BL<15>_XI0/XI1/XI0/MM0_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI0/MM1 N_XI0/XI1/XI0/NET33_XI0/XI1/XI0/MM1_d
+ N_XI0/XI1/XI0/NET34_XI0/XI1/XI0/MM1_g N_VSS_XI0/XI1/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI0/MM9 N_XI0/XI1/XI0/NET36_XI0/XI1/XI0/MM9_d N_WL<3>_XI0/XI1/XI0/MM9_g
+ N_BL<15>_XI0/XI1/XI0/MM9_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI0/MM6 N_XI0/XI1/XI0/NET35_XI0/XI1/XI0/MM6_d
+ N_XI0/XI1/XI0/NET36_XI0/XI1/XI0/MM6_g N_VSS_XI0/XI1/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI0/MM7 N_XI0/XI1/XI0/NET36_XI0/XI1/XI0/MM7_d
+ N_XI0/XI1/XI0/NET35_XI0/XI1/XI0/MM7_g N_VSS_XI0/XI1/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI0/MM8 N_XI0/XI1/XI0/NET35_XI0/XI1/XI0/MM8_d N_WL<3>_XI0/XI1/XI0/MM8_g
+ N_BLN<15>_XI0/XI1/XI0/MM8_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI0/MM5 N_XI0/XI1/XI0/NET34_XI0/XI1/XI0/MM5_d
+ N_XI0/XI1/XI0/NET33_XI0/XI1/XI0/MM5_g N_VDD_XI0/XI1/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI0/MM4 N_XI0/XI1/XI0/NET33_XI0/XI1/XI0/MM4_d
+ N_XI0/XI1/XI0/NET34_XI0/XI1/XI0/MM4_g N_VDD_XI0/XI1/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI0/MM10 N_XI0/XI1/XI0/NET35_XI0/XI1/XI0/MM10_d
+ N_XI0/XI1/XI0/NET36_XI0/XI1/XI0/MM10_g N_VDD_XI0/XI1/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI0/MM11 N_XI0/XI1/XI0/NET36_XI0/XI1/XI0/MM11_d
+ N_XI0/XI1/XI0/NET35_XI0/XI1/XI0/MM11_g N_VDD_XI0/XI1/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI1/MM2 N_XI0/XI1/XI1/NET34_XI0/XI1/XI1/MM2_d
+ N_XI0/XI1/XI1/NET33_XI0/XI1/XI1/MM2_g N_VSS_XI0/XI1/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI1/MM3 N_XI0/XI1/XI1/NET33_XI0/XI1/XI1/MM3_d N_WL<2>_XI0/XI1/XI1/MM3_g
+ N_BLN<14>_XI0/XI1/XI1/MM3_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI1/MM0 N_XI0/XI1/XI1/NET34_XI0/XI1/XI1/MM0_d N_WL<2>_XI0/XI1/XI1/MM0_g
+ N_BL<14>_XI0/XI1/XI1/MM0_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI1/MM1 N_XI0/XI1/XI1/NET33_XI0/XI1/XI1/MM1_d
+ N_XI0/XI1/XI1/NET34_XI0/XI1/XI1/MM1_g N_VSS_XI0/XI1/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI1/MM9 N_XI0/XI1/XI1/NET36_XI0/XI1/XI1/MM9_d N_WL<3>_XI0/XI1/XI1/MM9_g
+ N_BL<14>_XI0/XI1/XI1/MM9_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI1/MM6 N_XI0/XI1/XI1/NET35_XI0/XI1/XI1/MM6_d
+ N_XI0/XI1/XI1/NET36_XI0/XI1/XI1/MM6_g N_VSS_XI0/XI1/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI1/MM7 N_XI0/XI1/XI1/NET36_XI0/XI1/XI1/MM7_d
+ N_XI0/XI1/XI1/NET35_XI0/XI1/XI1/MM7_g N_VSS_XI0/XI1/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI1/MM8 N_XI0/XI1/XI1/NET35_XI0/XI1/XI1/MM8_d N_WL<3>_XI0/XI1/XI1/MM8_g
+ N_BLN<14>_XI0/XI1/XI1/MM8_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI1/MM5 N_XI0/XI1/XI1/NET34_XI0/XI1/XI1/MM5_d
+ N_XI0/XI1/XI1/NET33_XI0/XI1/XI1/MM5_g N_VDD_XI0/XI1/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI1/MM4 N_XI0/XI1/XI1/NET33_XI0/XI1/XI1/MM4_d
+ N_XI0/XI1/XI1/NET34_XI0/XI1/XI1/MM4_g N_VDD_XI0/XI1/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI1/MM10 N_XI0/XI1/XI1/NET35_XI0/XI1/XI1/MM10_d
+ N_XI0/XI1/XI1/NET36_XI0/XI1/XI1/MM10_g N_VDD_XI0/XI1/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI1/MM11 N_XI0/XI1/XI1/NET36_XI0/XI1/XI1/MM11_d
+ N_XI0/XI1/XI1/NET35_XI0/XI1/XI1/MM11_g N_VDD_XI0/XI1/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI2/MM2 N_XI0/XI1/XI2/NET34_XI0/XI1/XI2/MM2_d
+ N_XI0/XI1/XI2/NET33_XI0/XI1/XI2/MM2_g N_VSS_XI0/XI1/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI2/MM3 N_XI0/XI1/XI2/NET33_XI0/XI1/XI2/MM3_d N_WL<2>_XI0/XI1/XI2/MM3_g
+ N_BLN<13>_XI0/XI1/XI2/MM3_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI2/MM0 N_XI0/XI1/XI2/NET34_XI0/XI1/XI2/MM0_d N_WL<2>_XI0/XI1/XI2/MM0_g
+ N_BL<13>_XI0/XI1/XI2/MM0_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI2/MM1 N_XI0/XI1/XI2/NET33_XI0/XI1/XI2/MM1_d
+ N_XI0/XI1/XI2/NET34_XI0/XI1/XI2/MM1_g N_VSS_XI0/XI1/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI2/MM9 N_XI0/XI1/XI2/NET36_XI0/XI1/XI2/MM9_d N_WL<3>_XI0/XI1/XI2/MM9_g
+ N_BL<13>_XI0/XI1/XI2/MM9_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI2/MM6 N_XI0/XI1/XI2/NET35_XI0/XI1/XI2/MM6_d
+ N_XI0/XI1/XI2/NET36_XI0/XI1/XI2/MM6_g N_VSS_XI0/XI1/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI2/MM7 N_XI0/XI1/XI2/NET36_XI0/XI1/XI2/MM7_d
+ N_XI0/XI1/XI2/NET35_XI0/XI1/XI2/MM7_g N_VSS_XI0/XI1/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI2/MM8 N_XI0/XI1/XI2/NET35_XI0/XI1/XI2/MM8_d N_WL<3>_XI0/XI1/XI2/MM8_g
+ N_BLN<13>_XI0/XI1/XI2/MM8_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI2/MM5 N_XI0/XI1/XI2/NET34_XI0/XI1/XI2/MM5_d
+ N_XI0/XI1/XI2/NET33_XI0/XI1/XI2/MM5_g N_VDD_XI0/XI1/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI2/MM4 N_XI0/XI1/XI2/NET33_XI0/XI1/XI2/MM4_d
+ N_XI0/XI1/XI2/NET34_XI0/XI1/XI2/MM4_g N_VDD_XI0/XI1/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI2/MM10 N_XI0/XI1/XI2/NET35_XI0/XI1/XI2/MM10_d
+ N_XI0/XI1/XI2/NET36_XI0/XI1/XI2/MM10_g N_VDD_XI0/XI1/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI2/MM11 N_XI0/XI1/XI2/NET36_XI0/XI1/XI2/MM11_d
+ N_XI0/XI1/XI2/NET35_XI0/XI1/XI2/MM11_g N_VDD_XI0/XI1/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI3/MM2 N_XI0/XI1/XI3/NET34_XI0/XI1/XI3/MM2_d
+ N_XI0/XI1/XI3/NET33_XI0/XI1/XI3/MM2_g N_VSS_XI0/XI1/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI3/MM3 N_XI0/XI1/XI3/NET33_XI0/XI1/XI3/MM3_d N_WL<2>_XI0/XI1/XI3/MM3_g
+ N_BLN<12>_XI0/XI1/XI3/MM3_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI3/MM0 N_XI0/XI1/XI3/NET34_XI0/XI1/XI3/MM0_d N_WL<2>_XI0/XI1/XI3/MM0_g
+ N_BL<12>_XI0/XI1/XI3/MM0_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI3/MM1 N_XI0/XI1/XI3/NET33_XI0/XI1/XI3/MM1_d
+ N_XI0/XI1/XI3/NET34_XI0/XI1/XI3/MM1_g N_VSS_XI0/XI1/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI3/MM9 N_XI0/XI1/XI3/NET36_XI0/XI1/XI3/MM9_d N_WL<3>_XI0/XI1/XI3/MM9_g
+ N_BL<12>_XI0/XI1/XI3/MM9_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI3/MM6 N_XI0/XI1/XI3/NET35_XI0/XI1/XI3/MM6_d
+ N_XI0/XI1/XI3/NET36_XI0/XI1/XI3/MM6_g N_VSS_XI0/XI1/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI3/MM7 N_XI0/XI1/XI3/NET36_XI0/XI1/XI3/MM7_d
+ N_XI0/XI1/XI3/NET35_XI0/XI1/XI3/MM7_g N_VSS_XI0/XI1/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI3/MM8 N_XI0/XI1/XI3/NET35_XI0/XI1/XI3/MM8_d N_WL<3>_XI0/XI1/XI3/MM8_g
+ N_BLN<12>_XI0/XI1/XI3/MM8_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI3/MM5 N_XI0/XI1/XI3/NET34_XI0/XI1/XI3/MM5_d
+ N_XI0/XI1/XI3/NET33_XI0/XI1/XI3/MM5_g N_VDD_XI0/XI1/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI3/MM4 N_XI0/XI1/XI3/NET33_XI0/XI1/XI3/MM4_d
+ N_XI0/XI1/XI3/NET34_XI0/XI1/XI3/MM4_g N_VDD_XI0/XI1/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI3/MM10 N_XI0/XI1/XI3/NET35_XI0/XI1/XI3/MM10_d
+ N_XI0/XI1/XI3/NET36_XI0/XI1/XI3/MM10_g N_VDD_XI0/XI1/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI3/MM11 N_XI0/XI1/XI3/NET36_XI0/XI1/XI3/MM11_d
+ N_XI0/XI1/XI3/NET35_XI0/XI1/XI3/MM11_g N_VDD_XI0/XI1/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI4/MM2 N_XI0/XI1/XI4/NET34_XI0/XI1/XI4/MM2_d
+ N_XI0/XI1/XI4/NET33_XI0/XI1/XI4/MM2_g N_VSS_XI0/XI1/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI4/MM3 N_XI0/XI1/XI4/NET33_XI0/XI1/XI4/MM3_d N_WL<2>_XI0/XI1/XI4/MM3_g
+ N_BLN<11>_XI0/XI1/XI4/MM3_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI4/MM0 N_XI0/XI1/XI4/NET34_XI0/XI1/XI4/MM0_d N_WL<2>_XI0/XI1/XI4/MM0_g
+ N_BL<11>_XI0/XI1/XI4/MM0_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI4/MM1 N_XI0/XI1/XI4/NET33_XI0/XI1/XI4/MM1_d
+ N_XI0/XI1/XI4/NET34_XI0/XI1/XI4/MM1_g N_VSS_XI0/XI1/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI4/MM9 N_XI0/XI1/XI4/NET36_XI0/XI1/XI4/MM9_d N_WL<3>_XI0/XI1/XI4/MM9_g
+ N_BL<11>_XI0/XI1/XI4/MM9_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI4/MM6 N_XI0/XI1/XI4/NET35_XI0/XI1/XI4/MM6_d
+ N_XI0/XI1/XI4/NET36_XI0/XI1/XI4/MM6_g N_VSS_XI0/XI1/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI4/MM7 N_XI0/XI1/XI4/NET36_XI0/XI1/XI4/MM7_d
+ N_XI0/XI1/XI4/NET35_XI0/XI1/XI4/MM7_g N_VSS_XI0/XI1/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI4/MM8 N_XI0/XI1/XI4/NET35_XI0/XI1/XI4/MM8_d N_WL<3>_XI0/XI1/XI4/MM8_g
+ N_BLN<11>_XI0/XI1/XI4/MM8_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI4/MM5 N_XI0/XI1/XI4/NET34_XI0/XI1/XI4/MM5_d
+ N_XI0/XI1/XI4/NET33_XI0/XI1/XI4/MM5_g N_VDD_XI0/XI1/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI4/MM4 N_XI0/XI1/XI4/NET33_XI0/XI1/XI4/MM4_d
+ N_XI0/XI1/XI4/NET34_XI0/XI1/XI4/MM4_g N_VDD_XI0/XI1/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI4/MM10 N_XI0/XI1/XI4/NET35_XI0/XI1/XI4/MM10_d
+ N_XI0/XI1/XI4/NET36_XI0/XI1/XI4/MM10_g N_VDD_XI0/XI1/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI4/MM11 N_XI0/XI1/XI4/NET36_XI0/XI1/XI4/MM11_d
+ N_XI0/XI1/XI4/NET35_XI0/XI1/XI4/MM11_g N_VDD_XI0/XI1/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI5/MM2 N_XI0/XI1/XI5/NET34_XI0/XI1/XI5/MM2_d
+ N_XI0/XI1/XI5/NET33_XI0/XI1/XI5/MM2_g N_VSS_XI0/XI1/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI5/MM3 N_XI0/XI1/XI5/NET33_XI0/XI1/XI5/MM3_d N_WL<2>_XI0/XI1/XI5/MM3_g
+ N_BLN<10>_XI0/XI1/XI5/MM3_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI5/MM0 N_XI0/XI1/XI5/NET34_XI0/XI1/XI5/MM0_d N_WL<2>_XI0/XI1/XI5/MM0_g
+ N_BL<10>_XI0/XI1/XI5/MM0_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI5/MM1 N_XI0/XI1/XI5/NET33_XI0/XI1/XI5/MM1_d
+ N_XI0/XI1/XI5/NET34_XI0/XI1/XI5/MM1_g N_VSS_XI0/XI1/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI5/MM9 N_XI0/XI1/XI5/NET36_XI0/XI1/XI5/MM9_d N_WL<3>_XI0/XI1/XI5/MM9_g
+ N_BL<10>_XI0/XI1/XI5/MM9_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI5/MM6 N_XI0/XI1/XI5/NET35_XI0/XI1/XI5/MM6_d
+ N_XI0/XI1/XI5/NET36_XI0/XI1/XI5/MM6_g N_VSS_XI0/XI1/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI5/MM7 N_XI0/XI1/XI5/NET36_XI0/XI1/XI5/MM7_d
+ N_XI0/XI1/XI5/NET35_XI0/XI1/XI5/MM7_g N_VSS_XI0/XI1/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI5/MM8 N_XI0/XI1/XI5/NET35_XI0/XI1/XI5/MM8_d N_WL<3>_XI0/XI1/XI5/MM8_g
+ N_BLN<10>_XI0/XI1/XI5/MM8_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI5/MM5 N_XI0/XI1/XI5/NET34_XI0/XI1/XI5/MM5_d
+ N_XI0/XI1/XI5/NET33_XI0/XI1/XI5/MM5_g N_VDD_XI0/XI1/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI5/MM4 N_XI0/XI1/XI5/NET33_XI0/XI1/XI5/MM4_d
+ N_XI0/XI1/XI5/NET34_XI0/XI1/XI5/MM4_g N_VDD_XI0/XI1/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI5/MM10 N_XI0/XI1/XI5/NET35_XI0/XI1/XI5/MM10_d
+ N_XI0/XI1/XI5/NET36_XI0/XI1/XI5/MM10_g N_VDD_XI0/XI1/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI5/MM11 N_XI0/XI1/XI5/NET36_XI0/XI1/XI5/MM11_d
+ N_XI0/XI1/XI5/NET35_XI0/XI1/XI5/MM11_g N_VDD_XI0/XI1/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI6/MM2 N_XI0/XI1/XI6/NET34_XI0/XI1/XI6/MM2_d
+ N_XI0/XI1/XI6/NET33_XI0/XI1/XI6/MM2_g N_VSS_XI0/XI1/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI6/MM3 N_XI0/XI1/XI6/NET33_XI0/XI1/XI6/MM3_d N_WL<2>_XI0/XI1/XI6/MM3_g
+ N_BLN<9>_XI0/XI1/XI6/MM3_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI6/MM0 N_XI0/XI1/XI6/NET34_XI0/XI1/XI6/MM0_d N_WL<2>_XI0/XI1/XI6/MM0_g
+ N_BL<9>_XI0/XI1/XI6/MM0_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI6/MM1 N_XI0/XI1/XI6/NET33_XI0/XI1/XI6/MM1_d
+ N_XI0/XI1/XI6/NET34_XI0/XI1/XI6/MM1_g N_VSS_XI0/XI1/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI6/MM9 N_XI0/XI1/XI6/NET36_XI0/XI1/XI6/MM9_d N_WL<3>_XI0/XI1/XI6/MM9_g
+ N_BL<9>_XI0/XI1/XI6/MM9_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI6/MM6 N_XI0/XI1/XI6/NET35_XI0/XI1/XI6/MM6_d
+ N_XI0/XI1/XI6/NET36_XI0/XI1/XI6/MM6_g N_VSS_XI0/XI1/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI6/MM7 N_XI0/XI1/XI6/NET36_XI0/XI1/XI6/MM7_d
+ N_XI0/XI1/XI6/NET35_XI0/XI1/XI6/MM7_g N_VSS_XI0/XI1/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI6/MM8 N_XI0/XI1/XI6/NET35_XI0/XI1/XI6/MM8_d N_WL<3>_XI0/XI1/XI6/MM8_g
+ N_BLN<9>_XI0/XI1/XI6/MM8_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI6/MM5 N_XI0/XI1/XI6/NET34_XI0/XI1/XI6/MM5_d
+ N_XI0/XI1/XI6/NET33_XI0/XI1/XI6/MM5_g N_VDD_XI0/XI1/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI6/MM4 N_XI0/XI1/XI6/NET33_XI0/XI1/XI6/MM4_d
+ N_XI0/XI1/XI6/NET34_XI0/XI1/XI6/MM4_g N_VDD_XI0/XI1/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI6/MM10 N_XI0/XI1/XI6/NET35_XI0/XI1/XI6/MM10_d
+ N_XI0/XI1/XI6/NET36_XI0/XI1/XI6/MM10_g N_VDD_XI0/XI1/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI6/MM11 N_XI0/XI1/XI6/NET36_XI0/XI1/XI6/MM11_d
+ N_XI0/XI1/XI6/NET35_XI0/XI1/XI6/MM11_g N_VDD_XI0/XI1/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI7/MM2 N_XI0/XI1/XI7/NET34_XI0/XI1/XI7/MM2_d
+ N_XI0/XI1/XI7/NET33_XI0/XI1/XI7/MM2_g N_VSS_XI0/XI1/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI7/MM3 N_XI0/XI1/XI7/NET33_XI0/XI1/XI7/MM3_d N_WL<2>_XI0/XI1/XI7/MM3_g
+ N_BLN<8>_XI0/XI1/XI7/MM3_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI7/MM0 N_XI0/XI1/XI7/NET34_XI0/XI1/XI7/MM0_d N_WL<2>_XI0/XI1/XI7/MM0_g
+ N_BL<8>_XI0/XI1/XI7/MM0_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI7/MM1 N_XI0/XI1/XI7/NET33_XI0/XI1/XI7/MM1_d
+ N_XI0/XI1/XI7/NET34_XI0/XI1/XI7/MM1_g N_VSS_XI0/XI1/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI7/MM9 N_XI0/XI1/XI7/NET36_XI0/XI1/XI7/MM9_d N_WL<3>_XI0/XI1/XI7/MM9_g
+ N_BL<8>_XI0/XI1/XI7/MM9_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI7/MM6 N_XI0/XI1/XI7/NET35_XI0/XI1/XI7/MM6_d
+ N_XI0/XI1/XI7/NET36_XI0/XI1/XI7/MM6_g N_VSS_XI0/XI1/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI7/MM7 N_XI0/XI1/XI7/NET36_XI0/XI1/XI7/MM7_d
+ N_XI0/XI1/XI7/NET35_XI0/XI1/XI7/MM7_g N_VSS_XI0/XI1/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI7/MM8 N_XI0/XI1/XI7/NET35_XI0/XI1/XI7/MM8_d N_WL<3>_XI0/XI1/XI7/MM8_g
+ N_BLN<8>_XI0/XI1/XI7/MM8_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI7/MM5 N_XI0/XI1/XI7/NET34_XI0/XI1/XI7/MM5_d
+ N_XI0/XI1/XI7/NET33_XI0/XI1/XI7/MM5_g N_VDD_XI0/XI1/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI7/MM4 N_XI0/XI1/XI7/NET33_XI0/XI1/XI7/MM4_d
+ N_XI0/XI1/XI7/NET34_XI0/XI1/XI7/MM4_g N_VDD_XI0/XI1/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI7/MM10 N_XI0/XI1/XI7/NET35_XI0/XI1/XI7/MM10_d
+ N_XI0/XI1/XI7/NET36_XI0/XI1/XI7/MM10_g N_VDD_XI0/XI1/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI7/MM11 N_XI0/XI1/XI7/NET36_XI0/XI1/XI7/MM11_d
+ N_XI0/XI1/XI7/NET35_XI0/XI1/XI7/MM11_g N_VDD_XI0/XI1/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI8/MM2 N_XI0/XI1/XI8/NET34_XI0/XI1/XI8/MM2_d
+ N_XI0/XI1/XI8/NET33_XI0/XI1/XI8/MM2_g N_VSS_XI0/XI1/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI8/MM3 N_XI0/XI1/XI8/NET33_XI0/XI1/XI8/MM3_d N_WL<2>_XI0/XI1/XI8/MM3_g
+ N_BLN<7>_XI0/XI1/XI8/MM3_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI8/MM0 N_XI0/XI1/XI8/NET34_XI0/XI1/XI8/MM0_d N_WL<2>_XI0/XI1/XI8/MM0_g
+ N_BL<7>_XI0/XI1/XI8/MM0_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI8/MM1 N_XI0/XI1/XI8/NET33_XI0/XI1/XI8/MM1_d
+ N_XI0/XI1/XI8/NET34_XI0/XI1/XI8/MM1_g N_VSS_XI0/XI1/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI8/MM9 N_XI0/XI1/XI8/NET36_XI0/XI1/XI8/MM9_d N_WL<3>_XI0/XI1/XI8/MM9_g
+ N_BL<7>_XI0/XI1/XI8/MM9_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI8/MM6 N_XI0/XI1/XI8/NET35_XI0/XI1/XI8/MM6_d
+ N_XI0/XI1/XI8/NET36_XI0/XI1/XI8/MM6_g N_VSS_XI0/XI1/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI8/MM7 N_XI0/XI1/XI8/NET36_XI0/XI1/XI8/MM7_d
+ N_XI0/XI1/XI8/NET35_XI0/XI1/XI8/MM7_g N_VSS_XI0/XI1/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI8/MM8 N_XI0/XI1/XI8/NET35_XI0/XI1/XI8/MM8_d N_WL<3>_XI0/XI1/XI8/MM8_g
+ N_BLN<7>_XI0/XI1/XI8/MM8_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI8/MM5 N_XI0/XI1/XI8/NET34_XI0/XI1/XI8/MM5_d
+ N_XI0/XI1/XI8/NET33_XI0/XI1/XI8/MM5_g N_VDD_XI0/XI1/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI8/MM4 N_XI0/XI1/XI8/NET33_XI0/XI1/XI8/MM4_d
+ N_XI0/XI1/XI8/NET34_XI0/XI1/XI8/MM4_g N_VDD_XI0/XI1/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI8/MM10 N_XI0/XI1/XI8/NET35_XI0/XI1/XI8/MM10_d
+ N_XI0/XI1/XI8/NET36_XI0/XI1/XI8/MM10_g N_VDD_XI0/XI1/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI8/MM11 N_XI0/XI1/XI8/NET36_XI0/XI1/XI8/MM11_d
+ N_XI0/XI1/XI8/NET35_XI0/XI1/XI8/MM11_g N_VDD_XI0/XI1/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI9/MM2 N_XI0/XI1/XI9/NET34_XI0/XI1/XI9/MM2_d
+ N_XI0/XI1/XI9/NET33_XI0/XI1/XI9/MM2_g N_VSS_XI0/XI1/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI9/MM3 N_XI0/XI1/XI9/NET33_XI0/XI1/XI9/MM3_d N_WL<2>_XI0/XI1/XI9/MM3_g
+ N_BLN<6>_XI0/XI1/XI9/MM3_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI9/MM0 N_XI0/XI1/XI9/NET34_XI0/XI1/XI9/MM0_d N_WL<2>_XI0/XI1/XI9/MM0_g
+ N_BL<6>_XI0/XI1/XI9/MM0_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI9/MM1 N_XI0/XI1/XI9/NET33_XI0/XI1/XI9/MM1_d
+ N_XI0/XI1/XI9/NET34_XI0/XI1/XI9/MM1_g N_VSS_XI0/XI1/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI9/MM9 N_XI0/XI1/XI9/NET36_XI0/XI1/XI9/MM9_d N_WL<3>_XI0/XI1/XI9/MM9_g
+ N_BL<6>_XI0/XI1/XI9/MM9_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI9/MM6 N_XI0/XI1/XI9/NET35_XI0/XI1/XI9/MM6_d
+ N_XI0/XI1/XI9/NET36_XI0/XI1/XI9/MM6_g N_VSS_XI0/XI1/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI9/MM7 N_XI0/XI1/XI9/NET36_XI0/XI1/XI9/MM7_d
+ N_XI0/XI1/XI9/NET35_XI0/XI1/XI9/MM7_g N_VSS_XI0/XI1/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI9/MM8 N_XI0/XI1/XI9/NET35_XI0/XI1/XI9/MM8_d N_WL<3>_XI0/XI1/XI9/MM8_g
+ N_BLN<6>_XI0/XI1/XI9/MM8_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI1/XI9/MM5 N_XI0/XI1/XI9/NET34_XI0/XI1/XI9/MM5_d
+ N_XI0/XI1/XI9/NET33_XI0/XI1/XI9/MM5_g N_VDD_XI0/XI1/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI9/MM4 N_XI0/XI1/XI9/NET33_XI0/XI1/XI9/MM4_d
+ N_XI0/XI1/XI9/NET34_XI0/XI1/XI9/MM4_g N_VDD_XI0/XI1/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI9/MM10 N_XI0/XI1/XI9/NET35_XI0/XI1/XI9/MM10_d
+ N_XI0/XI1/XI9/NET36_XI0/XI1/XI9/MM10_g N_VDD_XI0/XI1/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI9/MM11 N_XI0/XI1/XI9/NET36_XI0/XI1/XI9/MM11_d
+ N_XI0/XI1/XI9/NET35_XI0/XI1/XI9/MM11_g N_VDD_XI0/XI1/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI10/MM2 N_XI0/XI1/XI10/NET34_XI0/XI1/XI10/MM2_d
+ N_XI0/XI1/XI10/NET33_XI0/XI1/XI10/MM2_g N_VSS_XI0/XI1/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM3 N_XI0/XI1/XI10/NET33_XI0/XI1/XI10/MM3_d
+ N_WL<2>_XI0/XI1/XI10/MM3_g N_BLN<5>_XI0/XI1/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM0 N_XI0/XI1/XI10/NET34_XI0/XI1/XI10/MM0_d
+ N_WL<2>_XI0/XI1/XI10/MM0_g N_BL<5>_XI0/XI1/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM1 N_XI0/XI1/XI10/NET33_XI0/XI1/XI10/MM1_d
+ N_XI0/XI1/XI10/NET34_XI0/XI1/XI10/MM1_g N_VSS_XI0/XI1/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM9 N_XI0/XI1/XI10/NET36_XI0/XI1/XI10/MM9_d
+ N_WL<3>_XI0/XI1/XI10/MM9_g N_BL<5>_XI0/XI1/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM6 N_XI0/XI1/XI10/NET35_XI0/XI1/XI10/MM6_d
+ N_XI0/XI1/XI10/NET36_XI0/XI1/XI10/MM6_g N_VSS_XI0/XI1/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM7 N_XI0/XI1/XI10/NET36_XI0/XI1/XI10/MM7_d
+ N_XI0/XI1/XI10/NET35_XI0/XI1/XI10/MM7_g N_VSS_XI0/XI1/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM8 N_XI0/XI1/XI10/NET35_XI0/XI1/XI10/MM8_d
+ N_WL<3>_XI0/XI1/XI10/MM8_g N_BLN<5>_XI0/XI1/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI10/MM5 N_XI0/XI1/XI10/NET34_XI0/XI1/XI10/MM5_d
+ N_XI0/XI1/XI10/NET33_XI0/XI1/XI10/MM5_g N_VDD_XI0/XI1/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI10/MM4 N_XI0/XI1/XI10/NET33_XI0/XI1/XI10/MM4_d
+ N_XI0/XI1/XI10/NET34_XI0/XI1/XI10/MM4_g N_VDD_XI0/XI1/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI10/MM10 N_XI0/XI1/XI10/NET35_XI0/XI1/XI10/MM10_d
+ N_XI0/XI1/XI10/NET36_XI0/XI1/XI10/MM10_g N_VDD_XI0/XI1/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI10/MM11 N_XI0/XI1/XI10/NET36_XI0/XI1/XI10/MM11_d
+ N_XI0/XI1/XI10/NET35_XI0/XI1/XI10/MM11_g N_VDD_XI0/XI1/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI11/MM2 N_XI0/XI1/XI11/NET34_XI0/XI1/XI11/MM2_d
+ N_XI0/XI1/XI11/NET33_XI0/XI1/XI11/MM2_g N_VSS_XI0/XI1/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM3 N_XI0/XI1/XI11/NET33_XI0/XI1/XI11/MM3_d
+ N_WL<2>_XI0/XI1/XI11/MM3_g N_BLN<4>_XI0/XI1/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM0 N_XI0/XI1/XI11/NET34_XI0/XI1/XI11/MM0_d
+ N_WL<2>_XI0/XI1/XI11/MM0_g N_BL<4>_XI0/XI1/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM1 N_XI0/XI1/XI11/NET33_XI0/XI1/XI11/MM1_d
+ N_XI0/XI1/XI11/NET34_XI0/XI1/XI11/MM1_g N_VSS_XI0/XI1/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM9 N_XI0/XI1/XI11/NET36_XI0/XI1/XI11/MM9_d
+ N_WL<3>_XI0/XI1/XI11/MM9_g N_BL<4>_XI0/XI1/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM6 N_XI0/XI1/XI11/NET35_XI0/XI1/XI11/MM6_d
+ N_XI0/XI1/XI11/NET36_XI0/XI1/XI11/MM6_g N_VSS_XI0/XI1/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM7 N_XI0/XI1/XI11/NET36_XI0/XI1/XI11/MM7_d
+ N_XI0/XI1/XI11/NET35_XI0/XI1/XI11/MM7_g N_VSS_XI0/XI1/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM8 N_XI0/XI1/XI11/NET35_XI0/XI1/XI11/MM8_d
+ N_WL<3>_XI0/XI1/XI11/MM8_g N_BLN<4>_XI0/XI1/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI11/MM5 N_XI0/XI1/XI11/NET34_XI0/XI1/XI11/MM5_d
+ N_XI0/XI1/XI11/NET33_XI0/XI1/XI11/MM5_g N_VDD_XI0/XI1/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI11/MM4 N_XI0/XI1/XI11/NET33_XI0/XI1/XI11/MM4_d
+ N_XI0/XI1/XI11/NET34_XI0/XI1/XI11/MM4_g N_VDD_XI0/XI1/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI11/MM10 N_XI0/XI1/XI11/NET35_XI0/XI1/XI11/MM10_d
+ N_XI0/XI1/XI11/NET36_XI0/XI1/XI11/MM10_g N_VDD_XI0/XI1/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI11/MM11 N_XI0/XI1/XI11/NET36_XI0/XI1/XI11/MM11_d
+ N_XI0/XI1/XI11/NET35_XI0/XI1/XI11/MM11_g N_VDD_XI0/XI1/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI12/MM2 N_XI0/XI1/XI12/NET34_XI0/XI1/XI12/MM2_d
+ N_XI0/XI1/XI12/NET33_XI0/XI1/XI12/MM2_g N_VSS_XI0/XI1/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM3 N_XI0/XI1/XI12/NET33_XI0/XI1/XI12/MM3_d
+ N_WL<2>_XI0/XI1/XI12/MM3_g N_BLN<3>_XI0/XI1/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM0 N_XI0/XI1/XI12/NET34_XI0/XI1/XI12/MM0_d
+ N_WL<2>_XI0/XI1/XI12/MM0_g N_BL<3>_XI0/XI1/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM1 N_XI0/XI1/XI12/NET33_XI0/XI1/XI12/MM1_d
+ N_XI0/XI1/XI12/NET34_XI0/XI1/XI12/MM1_g N_VSS_XI0/XI1/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM9 N_XI0/XI1/XI12/NET36_XI0/XI1/XI12/MM9_d
+ N_WL<3>_XI0/XI1/XI12/MM9_g N_BL<3>_XI0/XI1/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM6 N_XI0/XI1/XI12/NET35_XI0/XI1/XI12/MM6_d
+ N_XI0/XI1/XI12/NET36_XI0/XI1/XI12/MM6_g N_VSS_XI0/XI1/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM7 N_XI0/XI1/XI12/NET36_XI0/XI1/XI12/MM7_d
+ N_XI0/XI1/XI12/NET35_XI0/XI1/XI12/MM7_g N_VSS_XI0/XI1/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM8 N_XI0/XI1/XI12/NET35_XI0/XI1/XI12/MM8_d
+ N_WL<3>_XI0/XI1/XI12/MM8_g N_BLN<3>_XI0/XI1/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI12/MM5 N_XI0/XI1/XI12/NET34_XI0/XI1/XI12/MM5_d
+ N_XI0/XI1/XI12/NET33_XI0/XI1/XI12/MM5_g N_VDD_XI0/XI1/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI12/MM4 N_XI0/XI1/XI12/NET33_XI0/XI1/XI12/MM4_d
+ N_XI0/XI1/XI12/NET34_XI0/XI1/XI12/MM4_g N_VDD_XI0/XI1/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI12/MM10 N_XI0/XI1/XI12/NET35_XI0/XI1/XI12/MM10_d
+ N_XI0/XI1/XI12/NET36_XI0/XI1/XI12/MM10_g N_VDD_XI0/XI1/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI12/MM11 N_XI0/XI1/XI12/NET36_XI0/XI1/XI12/MM11_d
+ N_XI0/XI1/XI12/NET35_XI0/XI1/XI12/MM11_g N_VDD_XI0/XI1/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI13/MM2 N_XI0/XI1/XI13/NET34_XI0/XI1/XI13/MM2_d
+ N_XI0/XI1/XI13/NET33_XI0/XI1/XI13/MM2_g N_VSS_XI0/XI1/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM3 N_XI0/XI1/XI13/NET33_XI0/XI1/XI13/MM3_d
+ N_WL<2>_XI0/XI1/XI13/MM3_g N_BLN<2>_XI0/XI1/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM0 N_XI0/XI1/XI13/NET34_XI0/XI1/XI13/MM0_d
+ N_WL<2>_XI0/XI1/XI13/MM0_g N_BL<2>_XI0/XI1/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM1 N_XI0/XI1/XI13/NET33_XI0/XI1/XI13/MM1_d
+ N_XI0/XI1/XI13/NET34_XI0/XI1/XI13/MM1_g N_VSS_XI0/XI1/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM9 N_XI0/XI1/XI13/NET36_XI0/XI1/XI13/MM9_d
+ N_WL<3>_XI0/XI1/XI13/MM9_g N_BL<2>_XI0/XI1/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM6 N_XI0/XI1/XI13/NET35_XI0/XI1/XI13/MM6_d
+ N_XI0/XI1/XI13/NET36_XI0/XI1/XI13/MM6_g N_VSS_XI0/XI1/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM7 N_XI0/XI1/XI13/NET36_XI0/XI1/XI13/MM7_d
+ N_XI0/XI1/XI13/NET35_XI0/XI1/XI13/MM7_g N_VSS_XI0/XI1/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM8 N_XI0/XI1/XI13/NET35_XI0/XI1/XI13/MM8_d
+ N_WL<3>_XI0/XI1/XI13/MM8_g N_BLN<2>_XI0/XI1/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI13/MM5 N_XI0/XI1/XI13/NET34_XI0/XI1/XI13/MM5_d
+ N_XI0/XI1/XI13/NET33_XI0/XI1/XI13/MM5_g N_VDD_XI0/XI1/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI13/MM4 N_XI0/XI1/XI13/NET33_XI0/XI1/XI13/MM4_d
+ N_XI0/XI1/XI13/NET34_XI0/XI1/XI13/MM4_g N_VDD_XI0/XI1/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI13/MM10 N_XI0/XI1/XI13/NET35_XI0/XI1/XI13/MM10_d
+ N_XI0/XI1/XI13/NET36_XI0/XI1/XI13/MM10_g N_VDD_XI0/XI1/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI13/MM11 N_XI0/XI1/XI13/NET36_XI0/XI1/XI13/MM11_d
+ N_XI0/XI1/XI13/NET35_XI0/XI1/XI13/MM11_g N_VDD_XI0/XI1/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI14/MM2 N_XI0/XI1/XI14/NET34_XI0/XI1/XI14/MM2_d
+ N_XI0/XI1/XI14/NET33_XI0/XI1/XI14/MM2_g N_VSS_XI0/XI1/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM3 N_XI0/XI1/XI14/NET33_XI0/XI1/XI14/MM3_d
+ N_WL<2>_XI0/XI1/XI14/MM3_g N_BLN<1>_XI0/XI1/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM0 N_XI0/XI1/XI14/NET34_XI0/XI1/XI14/MM0_d
+ N_WL<2>_XI0/XI1/XI14/MM0_g N_BL<1>_XI0/XI1/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM1 N_XI0/XI1/XI14/NET33_XI0/XI1/XI14/MM1_d
+ N_XI0/XI1/XI14/NET34_XI0/XI1/XI14/MM1_g N_VSS_XI0/XI1/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM9 N_XI0/XI1/XI14/NET36_XI0/XI1/XI14/MM9_d
+ N_WL<3>_XI0/XI1/XI14/MM9_g N_BL<1>_XI0/XI1/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM6 N_XI0/XI1/XI14/NET35_XI0/XI1/XI14/MM6_d
+ N_XI0/XI1/XI14/NET36_XI0/XI1/XI14/MM6_g N_VSS_XI0/XI1/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM7 N_XI0/XI1/XI14/NET36_XI0/XI1/XI14/MM7_d
+ N_XI0/XI1/XI14/NET35_XI0/XI1/XI14/MM7_g N_VSS_XI0/XI1/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM8 N_XI0/XI1/XI14/NET35_XI0/XI1/XI14/MM8_d
+ N_WL<3>_XI0/XI1/XI14/MM8_g N_BLN<1>_XI0/XI1/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI14/MM5 N_XI0/XI1/XI14/NET34_XI0/XI1/XI14/MM5_d
+ N_XI0/XI1/XI14/NET33_XI0/XI1/XI14/MM5_g N_VDD_XI0/XI1/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI14/MM4 N_XI0/XI1/XI14/NET33_XI0/XI1/XI14/MM4_d
+ N_XI0/XI1/XI14/NET34_XI0/XI1/XI14/MM4_g N_VDD_XI0/XI1/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI14/MM10 N_XI0/XI1/XI14/NET35_XI0/XI1/XI14/MM10_d
+ N_XI0/XI1/XI14/NET36_XI0/XI1/XI14/MM10_g N_VDD_XI0/XI1/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI14/MM11 N_XI0/XI1/XI14/NET36_XI0/XI1/XI14/MM11_d
+ N_XI0/XI1/XI14/NET35_XI0/XI1/XI14/MM11_g N_VDD_XI0/XI1/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI15/MM2 N_XI0/XI1/XI15/NET34_XI0/XI1/XI15/MM2_d
+ N_XI0/XI1/XI15/NET33_XI0/XI1/XI15/MM2_g N_VSS_XI0/XI1/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM3 N_XI0/XI1/XI15/NET33_XI0/XI1/XI15/MM3_d
+ N_WL<2>_XI0/XI1/XI15/MM3_g N_BLN<0>_XI0/XI1/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM0 N_XI0/XI1/XI15/NET34_XI0/XI1/XI15/MM0_d
+ N_WL<2>_XI0/XI1/XI15/MM0_g N_BL<0>_XI0/XI1/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM1 N_XI0/XI1/XI15/NET33_XI0/XI1/XI15/MM1_d
+ N_XI0/XI1/XI15/NET34_XI0/XI1/XI15/MM1_g N_VSS_XI0/XI1/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM9 N_XI0/XI1/XI15/NET36_XI0/XI1/XI15/MM9_d
+ N_WL<3>_XI0/XI1/XI15/MM9_g N_BL<0>_XI0/XI1/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM6 N_XI0/XI1/XI15/NET35_XI0/XI1/XI15/MM6_d
+ N_XI0/XI1/XI15/NET36_XI0/XI1/XI15/MM6_g N_VSS_XI0/XI1/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM7 N_XI0/XI1/XI15/NET36_XI0/XI1/XI15/MM7_d
+ N_XI0/XI1/XI15/NET35_XI0/XI1/XI15/MM7_g N_VSS_XI0/XI1/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM8 N_XI0/XI1/XI15/NET35_XI0/XI1/XI15/MM8_d
+ N_WL<3>_XI0/XI1/XI15/MM8_g N_BLN<0>_XI0/XI1/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/XI15/MM5 N_XI0/XI1/XI15/NET34_XI0/XI1/XI15/MM5_d
+ N_XI0/XI1/XI15/NET33_XI0/XI1/XI15/MM5_g N_VDD_XI0/XI1/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI15/MM4 N_XI0/XI1/XI15/NET33_XI0/XI1/XI15/MM4_d
+ N_XI0/XI1/XI15/NET34_XI0/XI1/XI15/MM4_g N_VDD_XI0/XI1/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI15/MM10 N_XI0/XI1/XI15/NET35_XI0/XI1/XI15/MM10_d
+ N_XI0/XI1/XI15/NET36_XI0/XI1/XI15/MM10_g N_VDD_XI0/XI1/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/XI15/MM11 N_XI0/XI1/XI15/NET36_XI0/XI1/XI15/MM11_d
+ N_XI0/XI1/XI15/NET35_XI0/XI1/XI15/MM11_g N_VDD_XI0/XI1/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI0/MM2 N_XI0/XI4/XI0/NET34_XI0/XI4/XI0/MM2_d
+ N_XI0/XI4/XI0/NET33_XI0/XI4/XI0/MM2_g N_VSS_XI0/XI4/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI0/MM3 N_XI0/XI4/XI0/NET33_XI0/XI4/XI0/MM3_d N_WL<4>_XI0/XI4/XI0/MM3_g
+ N_BLN<15>_XI0/XI4/XI0/MM3_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI0/MM0 N_XI0/XI4/XI0/NET34_XI0/XI4/XI0/MM0_d N_WL<4>_XI0/XI4/XI0/MM0_g
+ N_BL<15>_XI0/XI4/XI0/MM0_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI0/MM1 N_XI0/XI4/XI0/NET33_XI0/XI4/XI0/MM1_d
+ N_XI0/XI4/XI0/NET34_XI0/XI4/XI0/MM1_g N_VSS_XI0/XI4/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI0/MM9 N_XI0/XI4/XI0/NET36_XI0/XI4/XI0/MM9_d N_WL<5>_XI0/XI4/XI0/MM9_g
+ N_BL<15>_XI0/XI4/XI0/MM9_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI0/MM6 N_XI0/XI4/XI0/NET35_XI0/XI4/XI0/MM6_d
+ N_XI0/XI4/XI0/NET36_XI0/XI4/XI0/MM6_g N_VSS_XI0/XI4/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI0/MM7 N_XI0/XI4/XI0/NET36_XI0/XI4/XI0/MM7_d
+ N_XI0/XI4/XI0/NET35_XI0/XI4/XI0/MM7_g N_VSS_XI0/XI4/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI0/MM8 N_XI0/XI4/XI0/NET35_XI0/XI4/XI0/MM8_d N_WL<5>_XI0/XI4/XI0/MM8_g
+ N_BLN<15>_XI0/XI4/XI0/MM8_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI0/MM5 N_XI0/XI4/XI0/NET34_XI0/XI4/XI0/MM5_d
+ N_XI0/XI4/XI0/NET33_XI0/XI4/XI0/MM5_g N_VDD_XI0/XI4/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI0/MM4 N_XI0/XI4/XI0/NET33_XI0/XI4/XI0/MM4_d
+ N_XI0/XI4/XI0/NET34_XI0/XI4/XI0/MM4_g N_VDD_XI0/XI4/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI0/MM10 N_XI0/XI4/XI0/NET35_XI0/XI4/XI0/MM10_d
+ N_XI0/XI4/XI0/NET36_XI0/XI4/XI0/MM10_g N_VDD_XI0/XI4/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI0/MM11 N_XI0/XI4/XI0/NET36_XI0/XI4/XI0/MM11_d
+ N_XI0/XI4/XI0/NET35_XI0/XI4/XI0/MM11_g N_VDD_XI0/XI4/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI1/MM2 N_XI0/XI4/XI1/NET34_XI0/XI4/XI1/MM2_d
+ N_XI0/XI4/XI1/NET33_XI0/XI4/XI1/MM2_g N_VSS_XI0/XI4/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI1/MM3 N_XI0/XI4/XI1/NET33_XI0/XI4/XI1/MM3_d N_WL<4>_XI0/XI4/XI1/MM3_g
+ N_BLN<14>_XI0/XI4/XI1/MM3_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI1/MM0 N_XI0/XI4/XI1/NET34_XI0/XI4/XI1/MM0_d N_WL<4>_XI0/XI4/XI1/MM0_g
+ N_BL<14>_XI0/XI4/XI1/MM0_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI1/MM1 N_XI0/XI4/XI1/NET33_XI0/XI4/XI1/MM1_d
+ N_XI0/XI4/XI1/NET34_XI0/XI4/XI1/MM1_g N_VSS_XI0/XI4/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI1/MM9 N_XI0/XI4/XI1/NET36_XI0/XI4/XI1/MM9_d N_WL<5>_XI0/XI4/XI1/MM9_g
+ N_BL<14>_XI0/XI4/XI1/MM9_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI1/MM6 N_XI0/XI4/XI1/NET35_XI0/XI4/XI1/MM6_d
+ N_XI0/XI4/XI1/NET36_XI0/XI4/XI1/MM6_g N_VSS_XI0/XI4/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI1/MM7 N_XI0/XI4/XI1/NET36_XI0/XI4/XI1/MM7_d
+ N_XI0/XI4/XI1/NET35_XI0/XI4/XI1/MM7_g N_VSS_XI0/XI4/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI1/MM8 N_XI0/XI4/XI1/NET35_XI0/XI4/XI1/MM8_d N_WL<5>_XI0/XI4/XI1/MM8_g
+ N_BLN<14>_XI0/XI4/XI1/MM8_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI1/MM5 N_XI0/XI4/XI1/NET34_XI0/XI4/XI1/MM5_d
+ N_XI0/XI4/XI1/NET33_XI0/XI4/XI1/MM5_g N_VDD_XI0/XI4/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI1/MM4 N_XI0/XI4/XI1/NET33_XI0/XI4/XI1/MM4_d
+ N_XI0/XI4/XI1/NET34_XI0/XI4/XI1/MM4_g N_VDD_XI0/XI4/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI1/MM10 N_XI0/XI4/XI1/NET35_XI0/XI4/XI1/MM10_d
+ N_XI0/XI4/XI1/NET36_XI0/XI4/XI1/MM10_g N_VDD_XI0/XI4/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI1/MM11 N_XI0/XI4/XI1/NET36_XI0/XI4/XI1/MM11_d
+ N_XI0/XI4/XI1/NET35_XI0/XI4/XI1/MM11_g N_VDD_XI0/XI4/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI2/MM2 N_XI0/XI4/XI2/NET34_XI0/XI4/XI2/MM2_d
+ N_XI0/XI4/XI2/NET33_XI0/XI4/XI2/MM2_g N_VSS_XI0/XI4/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI2/MM3 N_XI0/XI4/XI2/NET33_XI0/XI4/XI2/MM3_d N_WL<4>_XI0/XI4/XI2/MM3_g
+ N_BLN<13>_XI0/XI4/XI2/MM3_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI2/MM0 N_XI0/XI4/XI2/NET34_XI0/XI4/XI2/MM0_d N_WL<4>_XI0/XI4/XI2/MM0_g
+ N_BL<13>_XI0/XI4/XI2/MM0_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI2/MM1 N_XI0/XI4/XI2/NET33_XI0/XI4/XI2/MM1_d
+ N_XI0/XI4/XI2/NET34_XI0/XI4/XI2/MM1_g N_VSS_XI0/XI4/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI2/MM9 N_XI0/XI4/XI2/NET36_XI0/XI4/XI2/MM9_d N_WL<5>_XI0/XI4/XI2/MM9_g
+ N_BL<13>_XI0/XI4/XI2/MM9_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI2/MM6 N_XI0/XI4/XI2/NET35_XI0/XI4/XI2/MM6_d
+ N_XI0/XI4/XI2/NET36_XI0/XI4/XI2/MM6_g N_VSS_XI0/XI4/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI2/MM7 N_XI0/XI4/XI2/NET36_XI0/XI4/XI2/MM7_d
+ N_XI0/XI4/XI2/NET35_XI0/XI4/XI2/MM7_g N_VSS_XI0/XI4/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI2/MM8 N_XI0/XI4/XI2/NET35_XI0/XI4/XI2/MM8_d N_WL<5>_XI0/XI4/XI2/MM8_g
+ N_BLN<13>_XI0/XI4/XI2/MM8_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI2/MM5 N_XI0/XI4/XI2/NET34_XI0/XI4/XI2/MM5_d
+ N_XI0/XI4/XI2/NET33_XI0/XI4/XI2/MM5_g N_VDD_XI0/XI4/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI2/MM4 N_XI0/XI4/XI2/NET33_XI0/XI4/XI2/MM4_d
+ N_XI0/XI4/XI2/NET34_XI0/XI4/XI2/MM4_g N_VDD_XI0/XI4/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI2/MM10 N_XI0/XI4/XI2/NET35_XI0/XI4/XI2/MM10_d
+ N_XI0/XI4/XI2/NET36_XI0/XI4/XI2/MM10_g N_VDD_XI0/XI4/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI2/MM11 N_XI0/XI4/XI2/NET36_XI0/XI4/XI2/MM11_d
+ N_XI0/XI4/XI2/NET35_XI0/XI4/XI2/MM11_g N_VDD_XI0/XI4/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI3/MM2 N_XI0/XI4/XI3/NET34_XI0/XI4/XI3/MM2_d
+ N_XI0/XI4/XI3/NET33_XI0/XI4/XI3/MM2_g N_VSS_XI0/XI4/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI3/MM3 N_XI0/XI4/XI3/NET33_XI0/XI4/XI3/MM3_d N_WL<4>_XI0/XI4/XI3/MM3_g
+ N_BLN<12>_XI0/XI4/XI3/MM3_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI3/MM0 N_XI0/XI4/XI3/NET34_XI0/XI4/XI3/MM0_d N_WL<4>_XI0/XI4/XI3/MM0_g
+ N_BL<12>_XI0/XI4/XI3/MM0_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI3/MM1 N_XI0/XI4/XI3/NET33_XI0/XI4/XI3/MM1_d
+ N_XI0/XI4/XI3/NET34_XI0/XI4/XI3/MM1_g N_VSS_XI0/XI4/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI3/MM9 N_XI0/XI4/XI3/NET36_XI0/XI4/XI3/MM9_d N_WL<5>_XI0/XI4/XI3/MM9_g
+ N_BL<12>_XI0/XI4/XI3/MM9_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI3/MM6 N_XI0/XI4/XI3/NET35_XI0/XI4/XI3/MM6_d
+ N_XI0/XI4/XI3/NET36_XI0/XI4/XI3/MM6_g N_VSS_XI0/XI4/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI3/MM7 N_XI0/XI4/XI3/NET36_XI0/XI4/XI3/MM7_d
+ N_XI0/XI4/XI3/NET35_XI0/XI4/XI3/MM7_g N_VSS_XI0/XI4/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI3/MM8 N_XI0/XI4/XI3/NET35_XI0/XI4/XI3/MM8_d N_WL<5>_XI0/XI4/XI3/MM8_g
+ N_BLN<12>_XI0/XI4/XI3/MM8_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI3/MM5 N_XI0/XI4/XI3/NET34_XI0/XI4/XI3/MM5_d
+ N_XI0/XI4/XI3/NET33_XI0/XI4/XI3/MM5_g N_VDD_XI0/XI4/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI3/MM4 N_XI0/XI4/XI3/NET33_XI0/XI4/XI3/MM4_d
+ N_XI0/XI4/XI3/NET34_XI0/XI4/XI3/MM4_g N_VDD_XI0/XI4/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI3/MM10 N_XI0/XI4/XI3/NET35_XI0/XI4/XI3/MM10_d
+ N_XI0/XI4/XI3/NET36_XI0/XI4/XI3/MM10_g N_VDD_XI0/XI4/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI3/MM11 N_XI0/XI4/XI3/NET36_XI0/XI4/XI3/MM11_d
+ N_XI0/XI4/XI3/NET35_XI0/XI4/XI3/MM11_g N_VDD_XI0/XI4/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI4/MM2 N_XI0/XI4/XI4/NET34_XI0/XI4/XI4/MM2_d
+ N_XI0/XI4/XI4/NET33_XI0/XI4/XI4/MM2_g N_VSS_XI0/XI4/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI4/MM3 N_XI0/XI4/XI4/NET33_XI0/XI4/XI4/MM3_d N_WL<4>_XI0/XI4/XI4/MM3_g
+ N_BLN<11>_XI0/XI4/XI4/MM3_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI4/MM0 N_XI0/XI4/XI4/NET34_XI0/XI4/XI4/MM0_d N_WL<4>_XI0/XI4/XI4/MM0_g
+ N_BL<11>_XI0/XI4/XI4/MM0_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI4/MM1 N_XI0/XI4/XI4/NET33_XI0/XI4/XI4/MM1_d
+ N_XI0/XI4/XI4/NET34_XI0/XI4/XI4/MM1_g N_VSS_XI0/XI4/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI4/MM9 N_XI0/XI4/XI4/NET36_XI0/XI4/XI4/MM9_d N_WL<5>_XI0/XI4/XI4/MM9_g
+ N_BL<11>_XI0/XI4/XI4/MM9_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI4/MM6 N_XI0/XI4/XI4/NET35_XI0/XI4/XI4/MM6_d
+ N_XI0/XI4/XI4/NET36_XI0/XI4/XI4/MM6_g N_VSS_XI0/XI4/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI4/MM7 N_XI0/XI4/XI4/NET36_XI0/XI4/XI4/MM7_d
+ N_XI0/XI4/XI4/NET35_XI0/XI4/XI4/MM7_g N_VSS_XI0/XI4/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI4/MM8 N_XI0/XI4/XI4/NET35_XI0/XI4/XI4/MM8_d N_WL<5>_XI0/XI4/XI4/MM8_g
+ N_BLN<11>_XI0/XI4/XI4/MM8_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI4/MM5 N_XI0/XI4/XI4/NET34_XI0/XI4/XI4/MM5_d
+ N_XI0/XI4/XI4/NET33_XI0/XI4/XI4/MM5_g N_VDD_XI0/XI4/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI4/MM4 N_XI0/XI4/XI4/NET33_XI0/XI4/XI4/MM4_d
+ N_XI0/XI4/XI4/NET34_XI0/XI4/XI4/MM4_g N_VDD_XI0/XI4/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI4/MM10 N_XI0/XI4/XI4/NET35_XI0/XI4/XI4/MM10_d
+ N_XI0/XI4/XI4/NET36_XI0/XI4/XI4/MM10_g N_VDD_XI0/XI4/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI4/MM11 N_XI0/XI4/XI4/NET36_XI0/XI4/XI4/MM11_d
+ N_XI0/XI4/XI4/NET35_XI0/XI4/XI4/MM11_g N_VDD_XI0/XI4/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI5/MM2 N_XI0/XI4/XI5/NET34_XI0/XI4/XI5/MM2_d
+ N_XI0/XI4/XI5/NET33_XI0/XI4/XI5/MM2_g N_VSS_XI0/XI4/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI5/MM3 N_XI0/XI4/XI5/NET33_XI0/XI4/XI5/MM3_d N_WL<4>_XI0/XI4/XI5/MM3_g
+ N_BLN<10>_XI0/XI4/XI5/MM3_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI5/MM0 N_XI0/XI4/XI5/NET34_XI0/XI4/XI5/MM0_d N_WL<4>_XI0/XI4/XI5/MM0_g
+ N_BL<10>_XI0/XI4/XI5/MM0_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI5/MM1 N_XI0/XI4/XI5/NET33_XI0/XI4/XI5/MM1_d
+ N_XI0/XI4/XI5/NET34_XI0/XI4/XI5/MM1_g N_VSS_XI0/XI4/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI5/MM9 N_XI0/XI4/XI5/NET36_XI0/XI4/XI5/MM9_d N_WL<5>_XI0/XI4/XI5/MM9_g
+ N_BL<10>_XI0/XI4/XI5/MM9_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI5/MM6 N_XI0/XI4/XI5/NET35_XI0/XI4/XI5/MM6_d
+ N_XI0/XI4/XI5/NET36_XI0/XI4/XI5/MM6_g N_VSS_XI0/XI4/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI5/MM7 N_XI0/XI4/XI5/NET36_XI0/XI4/XI5/MM7_d
+ N_XI0/XI4/XI5/NET35_XI0/XI4/XI5/MM7_g N_VSS_XI0/XI4/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI5/MM8 N_XI0/XI4/XI5/NET35_XI0/XI4/XI5/MM8_d N_WL<5>_XI0/XI4/XI5/MM8_g
+ N_BLN<10>_XI0/XI4/XI5/MM8_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI5/MM5 N_XI0/XI4/XI5/NET34_XI0/XI4/XI5/MM5_d
+ N_XI0/XI4/XI5/NET33_XI0/XI4/XI5/MM5_g N_VDD_XI0/XI4/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI5/MM4 N_XI0/XI4/XI5/NET33_XI0/XI4/XI5/MM4_d
+ N_XI0/XI4/XI5/NET34_XI0/XI4/XI5/MM4_g N_VDD_XI0/XI4/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI5/MM10 N_XI0/XI4/XI5/NET35_XI0/XI4/XI5/MM10_d
+ N_XI0/XI4/XI5/NET36_XI0/XI4/XI5/MM10_g N_VDD_XI0/XI4/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI5/MM11 N_XI0/XI4/XI5/NET36_XI0/XI4/XI5/MM11_d
+ N_XI0/XI4/XI5/NET35_XI0/XI4/XI5/MM11_g N_VDD_XI0/XI4/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI6/MM2 N_XI0/XI4/XI6/NET34_XI0/XI4/XI6/MM2_d
+ N_XI0/XI4/XI6/NET33_XI0/XI4/XI6/MM2_g N_VSS_XI0/XI4/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI6/MM3 N_XI0/XI4/XI6/NET33_XI0/XI4/XI6/MM3_d N_WL<4>_XI0/XI4/XI6/MM3_g
+ N_BLN<9>_XI0/XI4/XI6/MM3_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI6/MM0 N_XI0/XI4/XI6/NET34_XI0/XI4/XI6/MM0_d N_WL<4>_XI0/XI4/XI6/MM0_g
+ N_BL<9>_XI0/XI4/XI6/MM0_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI6/MM1 N_XI0/XI4/XI6/NET33_XI0/XI4/XI6/MM1_d
+ N_XI0/XI4/XI6/NET34_XI0/XI4/XI6/MM1_g N_VSS_XI0/XI4/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI6/MM9 N_XI0/XI4/XI6/NET36_XI0/XI4/XI6/MM9_d N_WL<5>_XI0/XI4/XI6/MM9_g
+ N_BL<9>_XI0/XI4/XI6/MM9_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI6/MM6 N_XI0/XI4/XI6/NET35_XI0/XI4/XI6/MM6_d
+ N_XI0/XI4/XI6/NET36_XI0/XI4/XI6/MM6_g N_VSS_XI0/XI4/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI6/MM7 N_XI0/XI4/XI6/NET36_XI0/XI4/XI6/MM7_d
+ N_XI0/XI4/XI6/NET35_XI0/XI4/XI6/MM7_g N_VSS_XI0/XI4/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI6/MM8 N_XI0/XI4/XI6/NET35_XI0/XI4/XI6/MM8_d N_WL<5>_XI0/XI4/XI6/MM8_g
+ N_BLN<9>_XI0/XI4/XI6/MM8_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI6/MM5 N_XI0/XI4/XI6/NET34_XI0/XI4/XI6/MM5_d
+ N_XI0/XI4/XI6/NET33_XI0/XI4/XI6/MM5_g N_VDD_XI0/XI4/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI6/MM4 N_XI0/XI4/XI6/NET33_XI0/XI4/XI6/MM4_d
+ N_XI0/XI4/XI6/NET34_XI0/XI4/XI6/MM4_g N_VDD_XI0/XI4/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI6/MM10 N_XI0/XI4/XI6/NET35_XI0/XI4/XI6/MM10_d
+ N_XI0/XI4/XI6/NET36_XI0/XI4/XI6/MM10_g N_VDD_XI0/XI4/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI6/MM11 N_XI0/XI4/XI6/NET36_XI0/XI4/XI6/MM11_d
+ N_XI0/XI4/XI6/NET35_XI0/XI4/XI6/MM11_g N_VDD_XI0/XI4/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI7/MM2 N_XI0/XI4/XI7/NET34_XI0/XI4/XI7/MM2_d
+ N_XI0/XI4/XI7/NET33_XI0/XI4/XI7/MM2_g N_VSS_XI0/XI4/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI7/MM3 N_XI0/XI4/XI7/NET33_XI0/XI4/XI7/MM3_d N_WL<4>_XI0/XI4/XI7/MM3_g
+ N_BLN<8>_XI0/XI4/XI7/MM3_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI7/MM0 N_XI0/XI4/XI7/NET34_XI0/XI4/XI7/MM0_d N_WL<4>_XI0/XI4/XI7/MM0_g
+ N_BL<8>_XI0/XI4/XI7/MM0_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI7/MM1 N_XI0/XI4/XI7/NET33_XI0/XI4/XI7/MM1_d
+ N_XI0/XI4/XI7/NET34_XI0/XI4/XI7/MM1_g N_VSS_XI0/XI4/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI7/MM9 N_XI0/XI4/XI7/NET36_XI0/XI4/XI7/MM9_d N_WL<5>_XI0/XI4/XI7/MM9_g
+ N_BL<8>_XI0/XI4/XI7/MM9_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI7/MM6 N_XI0/XI4/XI7/NET35_XI0/XI4/XI7/MM6_d
+ N_XI0/XI4/XI7/NET36_XI0/XI4/XI7/MM6_g N_VSS_XI0/XI4/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI7/MM7 N_XI0/XI4/XI7/NET36_XI0/XI4/XI7/MM7_d
+ N_XI0/XI4/XI7/NET35_XI0/XI4/XI7/MM7_g N_VSS_XI0/XI4/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI7/MM8 N_XI0/XI4/XI7/NET35_XI0/XI4/XI7/MM8_d N_WL<5>_XI0/XI4/XI7/MM8_g
+ N_BLN<8>_XI0/XI4/XI7/MM8_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI7/MM5 N_XI0/XI4/XI7/NET34_XI0/XI4/XI7/MM5_d
+ N_XI0/XI4/XI7/NET33_XI0/XI4/XI7/MM5_g N_VDD_XI0/XI4/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI7/MM4 N_XI0/XI4/XI7/NET33_XI0/XI4/XI7/MM4_d
+ N_XI0/XI4/XI7/NET34_XI0/XI4/XI7/MM4_g N_VDD_XI0/XI4/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI7/MM10 N_XI0/XI4/XI7/NET35_XI0/XI4/XI7/MM10_d
+ N_XI0/XI4/XI7/NET36_XI0/XI4/XI7/MM10_g N_VDD_XI0/XI4/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI7/MM11 N_XI0/XI4/XI7/NET36_XI0/XI4/XI7/MM11_d
+ N_XI0/XI4/XI7/NET35_XI0/XI4/XI7/MM11_g N_VDD_XI0/XI4/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI8/MM2 N_XI0/XI4/XI8/NET34_XI0/XI4/XI8/MM2_d
+ N_XI0/XI4/XI8/NET33_XI0/XI4/XI8/MM2_g N_VSS_XI0/XI4/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI8/MM3 N_XI0/XI4/XI8/NET33_XI0/XI4/XI8/MM3_d N_WL<4>_XI0/XI4/XI8/MM3_g
+ N_BLN<7>_XI0/XI4/XI8/MM3_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI8/MM0 N_XI0/XI4/XI8/NET34_XI0/XI4/XI8/MM0_d N_WL<4>_XI0/XI4/XI8/MM0_g
+ N_BL<7>_XI0/XI4/XI8/MM0_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI8/MM1 N_XI0/XI4/XI8/NET33_XI0/XI4/XI8/MM1_d
+ N_XI0/XI4/XI8/NET34_XI0/XI4/XI8/MM1_g N_VSS_XI0/XI4/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI8/MM9 N_XI0/XI4/XI8/NET36_XI0/XI4/XI8/MM9_d N_WL<5>_XI0/XI4/XI8/MM9_g
+ N_BL<7>_XI0/XI4/XI8/MM9_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI8/MM6 N_XI0/XI4/XI8/NET35_XI0/XI4/XI8/MM6_d
+ N_XI0/XI4/XI8/NET36_XI0/XI4/XI8/MM6_g N_VSS_XI0/XI4/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI8/MM7 N_XI0/XI4/XI8/NET36_XI0/XI4/XI8/MM7_d
+ N_XI0/XI4/XI8/NET35_XI0/XI4/XI8/MM7_g N_VSS_XI0/XI4/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI8/MM8 N_XI0/XI4/XI8/NET35_XI0/XI4/XI8/MM8_d N_WL<5>_XI0/XI4/XI8/MM8_g
+ N_BLN<7>_XI0/XI4/XI8/MM8_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI8/MM5 N_XI0/XI4/XI8/NET34_XI0/XI4/XI8/MM5_d
+ N_XI0/XI4/XI8/NET33_XI0/XI4/XI8/MM5_g N_VDD_XI0/XI4/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI8/MM4 N_XI0/XI4/XI8/NET33_XI0/XI4/XI8/MM4_d
+ N_XI0/XI4/XI8/NET34_XI0/XI4/XI8/MM4_g N_VDD_XI0/XI4/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI8/MM10 N_XI0/XI4/XI8/NET35_XI0/XI4/XI8/MM10_d
+ N_XI0/XI4/XI8/NET36_XI0/XI4/XI8/MM10_g N_VDD_XI0/XI4/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI8/MM11 N_XI0/XI4/XI8/NET36_XI0/XI4/XI8/MM11_d
+ N_XI0/XI4/XI8/NET35_XI0/XI4/XI8/MM11_g N_VDD_XI0/XI4/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI9/MM2 N_XI0/XI4/XI9/NET34_XI0/XI4/XI9/MM2_d
+ N_XI0/XI4/XI9/NET33_XI0/XI4/XI9/MM2_g N_VSS_XI0/XI4/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI9/MM3 N_XI0/XI4/XI9/NET33_XI0/XI4/XI9/MM3_d N_WL<4>_XI0/XI4/XI9/MM3_g
+ N_BLN<6>_XI0/XI4/XI9/MM3_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI9/MM0 N_XI0/XI4/XI9/NET34_XI0/XI4/XI9/MM0_d N_WL<4>_XI0/XI4/XI9/MM0_g
+ N_BL<6>_XI0/XI4/XI9/MM0_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI9/MM1 N_XI0/XI4/XI9/NET33_XI0/XI4/XI9/MM1_d
+ N_XI0/XI4/XI9/NET34_XI0/XI4/XI9/MM1_g N_VSS_XI0/XI4/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI9/MM9 N_XI0/XI4/XI9/NET36_XI0/XI4/XI9/MM9_d N_WL<5>_XI0/XI4/XI9/MM9_g
+ N_BL<6>_XI0/XI4/XI9/MM9_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI9/MM6 N_XI0/XI4/XI9/NET35_XI0/XI4/XI9/MM6_d
+ N_XI0/XI4/XI9/NET36_XI0/XI4/XI9/MM6_g N_VSS_XI0/XI4/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI9/MM7 N_XI0/XI4/XI9/NET36_XI0/XI4/XI9/MM7_d
+ N_XI0/XI4/XI9/NET35_XI0/XI4/XI9/MM7_g N_VSS_XI0/XI4/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI9/MM8 N_XI0/XI4/XI9/NET35_XI0/XI4/XI9/MM8_d N_WL<5>_XI0/XI4/XI9/MM8_g
+ N_BLN<6>_XI0/XI4/XI9/MM8_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI4/XI9/MM5 N_XI0/XI4/XI9/NET34_XI0/XI4/XI9/MM5_d
+ N_XI0/XI4/XI9/NET33_XI0/XI4/XI9/MM5_g N_VDD_XI0/XI4/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI9/MM4 N_XI0/XI4/XI9/NET33_XI0/XI4/XI9/MM4_d
+ N_XI0/XI4/XI9/NET34_XI0/XI4/XI9/MM4_g N_VDD_XI0/XI4/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI9/MM10 N_XI0/XI4/XI9/NET35_XI0/XI4/XI9/MM10_d
+ N_XI0/XI4/XI9/NET36_XI0/XI4/XI9/MM10_g N_VDD_XI0/XI4/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI9/MM11 N_XI0/XI4/XI9/NET36_XI0/XI4/XI9/MM11_d
+ N_XI0/XI4/XI9/NET35_XI0/XI4/XI9/MM11_g N_VDD_XI0/XI4/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI10/MM2 N_XI0/XI4/XI10/NET34_XI0/XI4/XI10/MM2_d
+ N_XI0/XI4/XI10/NET33_XI0/XI4/XI10/MM2_g N_VSS_XI0/XI4/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM3 N_XI0/XI4/XI10/NET33_XI0/XI4/XI10/MM3_d
+ N_WL<4>_XI0/XI4/XI10/MM3_g N_BLN<5>_XI0/XI4/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM0 N_XI0/XI4/XI10/NET34_XI0/XI4/XI10/MM0_d
+ N_WL<4>_XI0/XI4/XI10/MM0_g N_BL<5>_XI0/XI4/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM1 N_XI0/XI4/XI10/NET33_XI0/XI4/XI10/MM1_d
+ N_XI0/XI4/XI10/NET34_XI0/XI4/XI10/MM1_g N_VSS_XI0/XI4/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM9 N_XI0/XI4/XI10/NET36_XI0/XI4/XI10/MM9_d
+ N_WL<5>_XI0/XI4/XI10/MM9_g N_BL<5>_XI0/XI4/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM6 N_XI0/XI4/XI10/NET35_XI0/XI4/XI10/MM6_d
+ N_XI0/XI4/XI10/NET36_XI0/XI4/XI10/MM6_g N_VSS_XI0/XI4/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM7 N_XI0/XI4/XI10/NET36_XI0/XI4/XI10/MM7_d
+ N_XI0/XI4/XI10/NET35_XI0/XI4/XI10/MM7_g N_VSS_XI0/XI4/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM8 N_XI0/XI4/XI10/NET35_XI0/XI4/XI10/MM8_d
+ N_WL<5>_XI0/XI4/XI10/MM8_g N_BLN<5>_XI0/XI4/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI10/MM5 N_XI0/XI4/XI10/NET34_XI0/XI4/XI10/MM5_d
+ N_XI0/XI4/XI10/NET33_XI0/XI4/XI10/MM5_g N_VDD_XI0/XI4/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI10/MM4 N_XI0/XI4/XI10/NET33_XI0/XI4/XI10/MM4_d
+ N_XI0/XI4/XI10/NET34_XI0/XI4/XI10/MM4_g N_VDD_XI0/XI4/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI10/MM10 N_XI0/XI4/XI10/NET35_XI0/XI4/XI10/MM10_d
+ N_XI0/XI4/XI10/NET36_XI0/XI4/XI10/MM10_g N_VDD_XI0/XI4/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI10/MM11 N_XI0/XI4/XI10/NET36_XI0/XI4/XI10/MM11_d
+ N_XI0/XI4/XI10/NET35_XI0/XI4/XI10/MM11_g N_VDD_XI0/XI4/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI11/MM2 N_XI0/XI4/XI11/NET34_XI0/XI4/XI11/MM2_d
+ N_XI0/XI4/XI11/NET33_XI0/XI4/XI11/MM2_g N_VSS_XI0/XI4/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM3 N_XI0/XI4/XI11/NET33_XI0/XI4/XI11/MM3_d
+ N_WL<4>_XI0/XI4/XI11/MM3_g N_BLN<4>_XI0/XI4/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM0 N_XI0/XI4/XI11/NET34_XI0/XI4/XI11/MM0_d
+ N_WL<4>_XI0/XI4/XI11/MM0_g N_BL<4>_XI0/XI4/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM1 N_XI0/XI4/XI11/NET33_XI0/XI4/XI11/MM1_d
+ N_XI0/XI4/XI11/NET34_XI0/XI4/XI11/MM1_g N_VSS_XI0/XI4/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM9 N_XI0/XI4/XI11/NET36_XI0/XI4/XI11/MM9_d
+ N_WL<5>_XI0/XI4/XI11/MM9_g N_BL<4>_XI0/XI4/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM6 N_XI0/XI4/XI11/NET35_XI0/XI4/XI11/MM6_d
+ N_XI0/XI4/XI11/NET36_XI0/XI4/XI11/MM6_g N_VSS_XI0/XI4/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM7 N_XI0/XI4/XI11/NET36_XI0/XI4/XI11/MM7_d
+ N_XI0/XI4/XI11/NET35_XI0/XI4/XI11/MM7_g N_VSS_XI0/XI4/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM8 N_XI0/XI4/XI11/NET35_XI0/XI4/XI11/MM8_d
+ N_WL<5>_XI0/XI4/XI11/MM8_g N_BLN<4>_XI0/XI4/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI11/MM5 N_XI0/XI4/XI11/NET34_XI0/XI4/XI11/MM5_d
+ N_XI0/XI4/XI11/NET33_XI0/XI4/XI11/MM5_g N_VDD_XI0/XI4/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI11/MM4 N_XI0/XI4/XI11/NET33_XI0/XI4/XI11/MM4_d
+ N_XI0/XI4/XI11/NET34_XI0/XI4/XI11/MM4_g N_VDD_XI0/XI4/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI11/MM10 N_XI0/XI4/XI11/NET35_XI0/XI4/XI11/MM10_d
+ N_XI0/XI4/XI11/NET36_XI0/XI4/XI11/MM10_g N_VDD_XI0/XI4/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI11/MM11 N_XI0/XI4/XI11/NET36_XI0/XI4/XI11/MM11_d
+ N_XI0/XI4/XI11/NET35_XI0/XI4/XI11/MM11_g N_VDD_XI0/XI4/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI12/MM2 N_XI0/XI4/XI12/NET34_XI0/XI4/XI12/MM2_d
+ N_XI0/XI4/XI12/NET33_XI0/XI4/XI12/MM2_g N_VSS_XI0/XI4/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM3 N_XI0/XI4/XI12/NET33_XI0/XI4/XI12/MM3_d
+ N_WL<4>_XI0/XI4/XI12/MM3_g N_BLN<3>_XI0/XI4/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM0 N_XI0/XI4/XI12/NET34_XI0/XI4/XI12/MM0_d
+ N_WL<4>_XI0/XI4/XI12/MM0_g N_BL<3>_XI0/XI4/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM1 N_XI0/XI4/XI12/NET33_XI0/XI4/XI12/MM1_d
+ N_XI0/XI4/XI12/NET34_XI0/XI4/XI12/MM1_g N_VSS_XI0/XI4/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM9 N_XI0/XI4/XI12/NET36_XI0/XI4/XI12/MM9_d
+ N_WL<5>_XI0/XI4/XI12/MM9_g N_BL<3>_XI0/XI4/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM6 N_XI0/XI4/XI12/NET35_XI0/XI4/XI12/MM6_d
+ N_XI0/XI4/XI12/NET36_XI0/XI4/XI12/MM6_g N_VSS_XI0/XI4/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM7 N_XI0/XI4/XI12/NET36_XI0/XI4/XI12/MM7_d
+ N_XI0/XI4/XI12/NET35_XI0/XI4/XI12/MM7_g N_VSS_XI0/XI4/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM8 N_XI0/XI4/XI12/NET35_XI0/XI4/XI12/MM8_d
+ N_WL<5>_XI0/XI4/XI12/MM8_g N_BLN<3>_XI0/XI4/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI12/MM5 N_XI0/XI4/XI12/NET34_XI0/XI4/XI12/MM5_d
+ N_XI0/XI4/XI12/NET33_XI0/XI4/XI12/MM5_g N_VDD_XI0/XI4/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI12/MM4 N_XI0/XI4/XI12/NET33_XI0/XI4/XI12/MM4_d
+ N_XI0/XI4/XI12/NET34_XI0/XI4/XI12/MM4_g N_VDD_XI0/XI4/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI12/MM10 N_XI0/XI4/XI12/NET35_XI0/XI4/XI12/MM10_d
+ N_XI0/XI4/XI12/NET36_XI0/XI4/XI12/MM10_g N_VDD_XI0/XI4/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI12/MM11 N_XI0/XI4/XI12/NET36_XI0/XI4/XI12/MM11_d
+ N_XI0/XI4/XI12/NET35_XI0/XI4/XI12/MM11_g N_VDD_XI0/XI4/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI13/MM2 N_XI0/XI4/XI13/NET34_XI0/XI4/XI13/MM2_d
+ N_XI0/XI4/XI13/NET33_XI0/XI4/XI13/MM2_g N_VSS_XI0/XI4/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM3 N_XI0/XI4/XI13/NET33_XI0/XI4/XI13/MM3_d
+ N_WL<4>_XI0/XI4/XI13/MM3_g N_BLN<2>_XI0/XI4/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM0 N_XI0/XI4/XI13/NET34_XI0/XI4/XI13/MM0_d
+ N_WL<4>_XI0/XI4/XI13/MM0_g N_BL<2>_XI0/XI4/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM1 N_XI0/XI4/XI13/NET33_XI0/XI4/XI13/MM1_d
+ N_XI0/XI4/XI13/NET34_XI0/XI4/XI13/MM1_g N_VSS_XI0/XI4/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM9 N_XI0/XI4/XI13/NET36_XI0/XI4/XI13/MM9_d
+ N_WL<5>_XI0/XI4/XI13/MM9_g N_BL<2>_XI0/XI4/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM6 N_XI0/XI4/XI13/NET35_XI0/XI4/XI13/MM6_d
+ N_XI0/XI4/XI13/NET36_XI0/XI4/XI13/MM6_g N_VSS_XI0/XI4/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM7 N_XI0/XI4/XI13/NET36_XI0/XI4/XI13/MM7_d
+ N_XI0/XI4/XI13/NET35_XI0/XI4/XI13/MM7_g N_VSS_XI0/XI4/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM8 N_XI0/XI4/XI13/NET35_XI0/XI4/XI13/MM8_d
+ N_WL<5>_XI0/XI4/XI13/MM8_g N_BLN<2>_XI0/XI4/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI13/MM5 N_XI0/XI4/XI13/NET34_XI0/XI4/XI13/MM5_d
+ N_XI0/XI4/XI13/NET33_XI0/XI4/XI13/MM5_g N_VDD_XI0/XI4/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI13/MM4 N_XI0/XI4/XI13/NET33_XI0/XI4/XI13/MM4_d
+ N_XI0/XI4/XI13/NET34_XI0/XI4/XI13/MM4_g N_VDD_XI0/XI4/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI13/MM10 N_XI0/XI4/XI13/NET35_XI0/XI4/XI13/MM10_d
+ N_XI0/XI4/XI13/NET36_XI0/XI4/XI13/MM10_g N_VDD_XI0/XI4/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI13/MM11 N_XI0/XI4/XI13/NET36_XI0/XI4/XI13/MM11_d
+ N_XI0/XI4/XI13/NET35_XI0/XI4/XI13/MM11_g N_VDD_XI0/XI4/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI14/MM2 N_XI0/XI4/XI14/NET34_XI0/XI4/XI14/MM2_d
+ N_XI0/XI4/XI14/NET33_XI0/XI4/XI14/MM2_g N_VSS_XI0/XI4/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM3 N_XI0/XI4/XI14/NET33_XI0/XI4/XI14/MM3_d
+ N_WL<4>_XI0/XI4/XI14/MM3_g N_BLN<1>_XI0/XI4/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM0 N_XI0/XI4/XI14/NET34_XI0/XI4/XI14/MM0_d
+ N_WL<4>_XI0/XI4/XI14/MM0_g N_BL<1>_XI0/XI4/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM1 N_XI0/XI4/XI14/NET33_XI0/XI4/XI14/MM1_d
+ N_XI0/XI4/XI14/NET34_XI0/XI4/XI14/MM1_g N_VSS_XI0/XI4/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM9 N_XI0/XI4/XI14/NET36_XI0/XI4/XI14/MM9_d
+ N_WL<5>_XI0/XI4/XI14/MM9_g N_BL<1>_XI0/XI4/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM6 N_XI0/XI4/XI14/NET35_XI0/XI4/XI14/MM6_d
+ N_XI0/XI4/XI14/NET36_XI0/XI4/XI14/MM6_g N_VSS_XI0/XI4/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM7 N_XI0/XI4/XI14/NET36_XI0/XI4/XI14/MM7_d
+ N_XI0/XI4/XI14/NET35_XI0/XI4/XI14/MM7_g N_VSS_XI0/XI4/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM8 N_XI0/XI4/XI14/NET35_XI0/XI4/XI14/MM8_d
+ N_WL<5>_XI0/XI4/XI14/MM8_g N_BLN<1>_XI0/XI4/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI14/MM5 N_XI0/XI4/XI14/NET34_XI0/XI4/XI14/MM5_d
+ N_XI0/XI4/XI14/NET33_XI0/XI4/XI14/MM5_g N_VDD_XI0/XI4/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI14/MM4 N_XI0/XI4/XI14/NET33_XI0/XI4/XI14/MM4_d
+ N_XI0/XI4/XI14/NET34_XI0/XI4/XI14/MM4_g N_VDD_XI0/XI4/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI14/MM10 N_XI0/XI4/XI14/NET35_XI0/XI4/XI14/MM10_d
+ N_XI0/XI4/XI14/NET36_XI0/XI4/XI14/MM10_g N_VDD_XI0/XI4/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI14/MM11 N_XI0/XI4/XI14/NET36_XI0/XI4/XI14/MM11_d
+ N_XI0/XI4/XI14/NET35_XI0/XI4/XI14/MM11_g N_VDD_XI0/XI4/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI15/MM2 N_XI0/XI4/XI15/NET34_XI0/XI4/XI15/MM2_d
+ N_XI0/XI4/XI15/NET33_XI0/XI4/XI15/MM2_g N_VSS_XI0/XI4/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM3 N_XI0/XI4/XI15/NET33_XI0/XI4/XI15/MM3_d
+ N_WL<4>_XI0/XI4/XI15/MM3_g N_BLN<0>_XI0/XI4/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM0 N_XI0/XI4/XI15/NET34_XI0/XI4/XI15/MM0_d
+ N_WL<4>_XI0/XI4/XI15/MM0_g N_BL<0>_XI0/XI4/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM1 N_XI0/XI4/XI15/NET33_XI0/XI4/XI15/MM1_d
+ N_XI0/XI4/XI15/NET34_XI0/XI4/XI15/MM1_g N_VSS_XI0/XI4/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM9 N_XI0/XI4/XI15/NET36_XI0/XI4/XI15/MM9_d
+ N_WL<5>_XI0/XI4/XI15/MM9_g N_BL<0>_XI0/XI4/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM6 N_XI0/XI4/XI15/NET35_XI0/XI4/XI15/MM6_d
+ N_XI0/XI4/XI15/NET36_XI0/XI4/XI15/MM6_g N_VSS_XI0/XI4/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM7 N_XI0/XI4/XI15/NET36_XI0/XI4/XI15/MM7_d
+ N_XI0/XI4/XI15/NET35_XI0/XI4/XI15/MM7_g N_VSS_XI0/XI4/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM8 N_XI0/XI4/XI15/NET35_XI0/XI4/XI15/MM8_d
+ N_WL<5>_XI0/XI4/XI15/MM8_g N_BLN<0>_XI0/XI4/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/XI15/MM5 N_XI0/XI4/XI15/NET34_XI0/XI4/XI15/MM5_d
+ N_XI0/XI4/XI15/NET33_XI0/XI4/XI15/MM5_g N_VDD_XI0/XI4/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI15/MM4 N_XI0/XI4/XI15/NET33_XI0/XI4/XI15/MM4_d
+ N_XI0/XI4/XI15/NET34_XI0/XI4/XI15/MM4_g N_VDD_XI0/XI4/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI15/MM10 N_XI0/XI4/XI15/NET35_XI0/XI4/XI15/MM10_d
+ N_XI0/XI4/XI15/NET36_XI0/XI4/XI15/MM10_g N_VDD_XI0/XI4/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/XI15/MM11 N_XI0/XI4/XI15/NET36_XI0/XI4/XI15/MM11_d
+ N_XI0/XI4/XI15/NET35_XI0/XI4/XI15/MM11_g N_VDD_XI0/XI4/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI0/MM2 N_XI0/XI5/XI0/NET34_XI0/XI5/XI0/MM2_d
+ N_XI0/XI5/XI0/NET33_XI0/XI5/XI0/MM2_g N_VSS_XI0/XI5/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI0/MM3 N_XI0/XI5/XI0/NET33_XI0/XI5/XI0/MM3_d N_WL<6>_XI0/XI5/XI0/MM3_g
+ N_BLN<15>_XI0/XI5/XI0/MM3_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI0/MM0 N_XI0/XI5/XI0/NET34_XI0/XI5/XI0/MM0_d N_WL<6>_XI0/XI5/XI0/MM0_g
+ N_BL<15>_XI0/XI5/XI0/MM0_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI0/MM1 N_XI0/XI5/XI0/NET33_XI0/XI5/XI0/MM1_d
+ N_XI0/XI5/XI0/NET34_XI0/XI5/XI0/MM1_g N_VSS_XI0/XI5/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI0/MM9 N_XI0/XI5/XI0/NET36_XI0/XI5/XI0/MM9_d N_WL<7>_XI0/XI5/XI0/MM9_g
+ N_BL<15>_XI0/XI5/XI0/MM9_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI0/MM6 N_XI0/XI5/XI0/NET35_XI0/XI5/XI0/MM6_d
+ N_XI0/XI5/XI0/NET36_XI0/XI5/XI0/MM6_g N_VSS_XI0/XI5/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI0/MM7 N_XI0/XI5/XI0/NET36_XI0/XI5/XI0/MM7_d
+ N_XI0/XI5/XI0/NET35_XI0/XI5/XI0/MM7_g N_VSS_XI0/XI5/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI0/MM8 N_XI0/XI5/XI0/NET35_XI0/XI5/XI0/MM8_d N_WL<7>_XI0/XI5/XI0/MM8_g
+ N_BLN<15>_XI0/XI5/XI0/MM8_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI0/MM5 N_XI0/XI5/XI0/NET34_XI0/XI5/XI0/MM5_d
+ N_XI0/XI5/XI0/NET33_XI0/XI5/XI0/MM5_g N_VDD_XI0/XI5/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI0/MM4 N_XI0/XI5/XI0/NET33_XI0/XI5/XI0/MM4_d
+ N_XI0/XI5/XI0/NET34_XI0/XI5/XI0/MM4_g N_VDD_XI0/XI5/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI0/MM10 N_XI0/XI5/XI0/NET35_XI0/XI5/XI0/MM10_d
+ N_XI0/XI5/XI0/NET36_XI0/XI5/XI0/MM10_g N_VDD_XI0/XI5/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI0/MM11 N_XI0/XI5/XI0/NET36_XI0/XI5/XI0/MM11_d
+ N_XI0/XI5/XI0/NET35_XI0/XI5/XI0/MM11_g N_VDD_XI0/XI5/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI1/MM2 N_XI0/XI5/XI1/NET34_XI0/XI5/XI1/MM2_d
+ N_XI0/XI5/XI1/NET33_XI0/XI5/XI1/MM2_g N_VSS_XI0/XI5/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI1/MM3 N_XI0/XI5/XI1/NET33_XI0/XI5/XI1/MM3_d N_WL<6>_XI0/XI5/XI1/MM3_g
+ N_BLN<14>_XI0/XI5/XI1/MM3_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI1/MM0 N_XI0/XI5/XI1/NET34_XI0/XI5/XI1/MM0_d N_WL<6>_XI0/XI5/XI1/MM0_g
+ N_BL<14>_XI0/XI5/XI1/MM0_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI1/MM1 N_XI0/XI5/XI1/NET33_XI0/XI5/XI1/MM1_d
+ N_XI0/XI5/XI1/NET34_XI0/XI5/XI1/MM1_g N_VSS_XI0/XI5/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI1/MM9 N_XI0/XI5/XI1/NET36_XI0/XI5/XI1/MM9_d N_WL<7>_XI0/XI5/XI1/MM9_g
+ N_BL<14>_XI0/XI5/XI1/MM9_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI1/MM6 N_XI0/XI5/XI1/NET35_XI0/XI5/XI1/MM6_d
+ N_XI0/XI5/XI1/NET36_XI0/XI5/XI1/MM6_g N_VSS_XI0/XI5/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI1/MM7 N_XI0/XI5/XI1/NET36_XI0/XI5/XI1/MM7_d
+ N_XI0/XI5/XI1/NET35_XI0/XI5/XI1/MM7_g N_VSS_XI0/XI5/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI1/MM8 N_XI0/XI5/XI1/NET35_XI0/XI5/XI1/MM8_d N_WL<7>_XI0/XI5/XI1/MM8_g
+ N_BLN<14>_XI0/XI5/XI1/MM8_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI1/MM5 N_XI0/XI5/XI1/NET34_XI0/XI5/XI1/MM5_d
+ N_XI0/XI5/XI1/NET33_XI0/XI5/XI1/MM5_g N_VDD_XI0/XI5/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI1/MM4 N_XI0/XI5/XI1/NET33_XI0/XI5/XI1/MM4_d
+ N_XI0/XI5/XI1/NET34_XI0/XI5/XI1/MM4_g N_VDD_XI0/XI5/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI1/MM10 N_XI0/XI5/XI1/NET35_XI0/XI5/XI1/MM10_d
+ N_XI0/XI5/XI1/NET36_XI0/XI5/XI1/MM10_g N_VDD_XI0/XI5/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI1/MM11 N_XI0/XI5/XI1/NET36_XI0/XI5/XI1/MM11_d
+ N_XI0/XI5/XI1/NET35_XI0/XI5/XI1/MM11_g N_VDD_XI0/XI5/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI2/MM2 N_XI0/XI5/XI2/NET34_XI0/XI5/XI2/MM2_d
+ N_XI0/XI5/XI2/NET33_XI0/XI5/XI2/MM2_g N_VSS_XI0/XI5/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI2/MM3 N_XI0/XI5/XI2/NET33_XI0/XI5/XI2/MM3_d N_WL<6>_XI0/XI5/XI2/MM3_g
+ N_BLN<13>_XI0/XI5/XI2/MM3_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI2/MM0 N_XI0/XI5/XI2/NET34_XI0/XI5/XI2/MM0_d N_WL<6>_XI0/XI5/XI2/MM0_g
+ N_BL<13>_XI0/XI5/XI2/MM0_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI2/MM1 N_XI0/XI5/XI2/NET33_XI0/XI5/XI2/MM1_d
+ N_XI0/XI5/XI2/NET34_XI0/XI5/XI2/MM1_g N_VSS_XI0/XI5/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI2/MM9 N_XI0/XI5/XI2/NET36_XI0/XI5/XI2/MM9_d N_WL<7>_XI0/XI5/XI2/MM9_g
+ N_BL<13>_XI0/XI5/XI2/MM9_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI2/MM6 N_XI0/XI5/XI2/NET35_XI0/XI5/XI2/MM6_d
+ N_XI0/XI5/XI2/NET36_XI0/XI5/XI2/MM6_g N_VSS_XI0/XI5/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI2/MM7 N_XI0/XI5/XI2/NET36_XI0/XI5/XI2/MM7_d
+ N_XI0/XI5/XI2/NET35_XI0/XI5/XI2/MM7_g N_VSS_XI0/XI5/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI2/MM8 N_XI0/XI5/XI2/NET35_XI0/XI5/XI2/MM8_d N_WL<7>_XI0/XI5/XI2/MM8_g
+ N_BLN<13>_XI0/XI5/XI2/MM8_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI2/MM5 N_XI0/XI5/XI2/NET34_XI0/XI5/XI2/MM5_d
+ N_XI0/XI5/XI2/NET33_XI0/XI5/XI2/MM5_g N_VDD_XI0/XI5/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI2/MM4 N_XI0/XI5/XI2/NET33_XI0/XI5/XI2/MM4_d
+ N_XI0/XI5/XI2/NET34_XI0/XI5/XI2/MM4_g N_VDD_XI0/XI5/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI2/MM10 N_XI0/XI5/XI2/NET35_XI0/XI5/XI2/MM10_d
+ N_XI0/XI5/XI2/NET36_XI0/XI5/XI2/MM10_g N_VDD_XI0/XI5/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI2/MM11 N_XI0/XI5/XI2/NET36_XI0/XI5/XI2/MM11_d
+ N_XI0/XI5/XI2/NET35_XI0/XI5/XI2/MM11_g N_VDD_XI0/XI5/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI3/MM2 N_XI0/XI5/XI3/NET34_XI0/XI5/XI3/MM2_d
+ N_XI0/XI5/XI3/NET33_XI0/XI5/XI3/MM2_g N_VSS_XI0/XI5/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI3/MM3 N_XI0/XI5/XI3/NET33_XI0/XI5/XI3/MM3_d N_WL<6>_XI0/XI5/XI3/MM3_g
+ N_BLN<12>_XI0/XI5/XI3/MM3_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI3/MM0 N_XI0/XI5/XI3/NET34_XI0/XI5/XI3/MM0_d N_WL<6>_XI0/XI5/XI3/MM0_g
+ N_BL<12>_XI0/XI5/XI3/MM0_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI3/MM1 N_XI0/XI5/XI3/NET33_XI0/XI5/XI3/MM1_d
+ N_XI0/XI5/XI3/NET34_XI0/XI5/XI3/MM1_g N_VSS_XI0/XI5/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI3/MM9 N_XI0/XI5/XI3/NET36_XI0/XI5/XI3/MM9_d N_WL<7>_XI0/XI5/XI3/MM9_g
+ N_BL<12>_XI0/XI5/XI3/MM9_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI3/MM6 N_XI0/XI5/XI3/NET35_XI0/XI5/XI3/MM6_d
+ N_XI0/XI5/XI3/NET36_XI0/XI5/XI3/MM6_g N_VSS_XI0/XI5/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI3/MM7 N_XI0/XI5/XI3/NET36_XI0/XI5/XI3/MM7_d
+ N_XI0/XI5/XI3/NET35_XI0/XI5/XI3/MM7_g N_VSS_XI0/XI5/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI3/MM8 N_XI0/XI5/XI3/NET35_XI0/XI5/XI3/MM8_d N_WL<7>_XI0/XI5/XI3/MM8_g
+ N_BLN<12>_XI0/XI5/XI3/MM8_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI3/MM5 N_XI0/XI5/XI3/NET34_XI0/XI5/XI3/MM5_d
+ N_XI0/XI5/XI3/NET33_XI0/XI5/XI3/MM5_g N_VDD_XI0/XI5/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI3/MM4 N_XI0/XI5/XI3/NET33_XI0/XI5/XI3/MM4_d
+ N_XI0/XI5/XI3/NET34_XI0/XI5/XI3/MM4_g N_VDD_XI0/XI5/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI3/MM10 N_XI0/XI5/XI3/NET35_XI0/XI5/XI3/MM10_d
+ N_XI0/XI5/XI3/NET36_XI0/XI5/XI3/MM10_g N_VDD_XI0/XI5/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI3/MM11 N_XI0/XI5/XI3/NET36_XI0/XI5/XI3/MM11_d
+ N_XI0/XI5/XI3/NET35_XI0/XI5/XI3/MM11_g N_VDD_XI0/XI5/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI4/MM2 N_XI0/XI5/XI4/NET34_XI0/XI5/XI4/MM2_d
+ N_XI0/XI5/XI4/NET33_XI0/XI5/XI4/MM2_g N_VSS_XI0/XI5/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI4/MM3 N_XI0/XI5/XI4/NET33_XI0/XI5/XI4/MM3_d N_WL<6>_XI0/XI5/XI4/MM3_g
+ N_BLN<11>_XI0/XI5/XI4/MM3_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI4/MM0 N_XI0/XI5/XI4/NET34_XI0/XI5/XI4/MM0_d N_WL<6>_XI0/XI5/XI4/MM0_g
+ N_BL<11>_XI0/XI5/XI4/MM0_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI4/MM1 N_XI0/XI5/XI4/NET33_XI0/XI5/XI4/MM1_d
+ N_XI0/XI5/XI4/NET34_XI0/XI5/XI4/MM1_g N_VSS_XI0/XI5/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI4/MM9 N_XI0/XI5/XI4/NET36_XI0/XI5/XI4/MM9_d N_WL<7>_XI0/XI5/XI4/MM9_g
+ N_BL<11>_XI0/XI5/XI4/MM9_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI4/MM6 N_XI0/XI5/XI4/NET35_XI0/XI5/XI4/MM6_d
+ N_XI0/XI5/XI4/NET36_XI0/XI5/XI4/MM6_g N_VSS_XI0/XI5/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI4/MM7 N_XI0/XI5/XI4/NET36_XI0/XI5/XI4/MM7_d
+ N_XI0/XI5/XI4/NET35_XI0/XI5/XI4/MM7_g N_VSS_XI0/XI5/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI4/MM8 N_XI0/XI5/XI4/NET35_XI0/XI5/XI4/MM8_d N_WL<7>_XI0/XI5/XI4/MM8_g
+ N_BLN<11>_XI0/XI5/XI4/MM8_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI4/MM5 N_XI0/XI5/XI4/NET34_XI0/XI5/XI4/MM5_d
+ N_XI0/XI5/XI4/NET33_XI0/XI5/XI4/MM5_g N_VDD_XI0/XI5/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI4/MM4 N_XI0/XI5/XI4/NET33_XI0/XI5/XI4/MM4_d
+ N_XI0/XI5/XI4/NET34_XI0/XI5/XI4/MM4_g N_VDD_XI0/XI5/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI4/MM10 N_XI0/XI5/XI4/NET35_XI0/XI5/XI4/MM10_d
+ N_XI0/XI5/XI4/NET36_XI0/XI5/XI4/MM10_g N_VDD_XI0/XI5/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI4/MM11 N_XI0/XI5/XI4/NET36_XI0/XI5/XI4/MM11_d
+ N_XI0/XI5/XI4/NET35_XI0/XI5/XI4/MM11_g N_VDD_XI0/XI5/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI5/MM2 N_XI0/XI5/XI5/NET34_XI0/XI5/XI5/MM2_d
+ N_XI0/XI5/XI5/NET33_XI0/XI5/XI5/MM2_g N_VSS_XI0/XI5/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI5/MM3 N_XI0/XI5/XI5/NET33_XI0/XI5/XI5/MM3_d N_WL<6>_XI0/XI5/XI5/MM3_g
+ N_BLN<10>_XI0/XI5/XI5/MM3_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI5/MM0 N_XI0/XI5/XI5/NET34_XI0/XI5/XI5/MM0_d N_WL<6>_XI0/XI5/XI5/MM0_g
+ N_BL<10>_XI0/XI5/XI5/MM0_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI5/MM1 N_XI0/XI5/XI5/NET33_XI0/XI5/XI5/MM1_d
+ N_XI0/XI5/XI5/NET34_XI0/XI5/XI5/MM1_g N_VSS_XI0/XI5/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI5/MM9 N_XI0/XI5/XI5/NET36_XI0/XI5/XI5/MM9_d N_WL<7>_XI0/XI5/XI5/MM9_g
+ N_BL<10>_XI0/XI5/XI5/MM9_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI5/MM6 N_XI0/XI5/XI5/NET35_XI0/XI5/XI5/MM6_d
+ N_XI0/XI5/XI5/NET36_XI0/XI5/XI5/MM6_g N_VSS_XI0/XI5/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI5/MM7 N_XI0/XI5/XI5/NET36_XI0/XI5/XI5/MM7_d
+ N_XI0/XI5/XI5/NET35_XI0/XI5/XI5/MM7_g N_VSS_XI0/XI5/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI5/MM8 N_XI0/XI5/XI5/NET35_XI0/XI5/XI5/MM8_d N_WL<7>_XI0/XI5/XI5/MM8_g
+ N_BLN<10>_XI0/XI5/XI5/MM8_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI5/MM5 N_XI0/XI5/XI5/NET34_XI0/XI5/XI5/MM5_d
+ N_XI0/XI5/XI5/NET33_XI0/XI5/XI5/MM5_g N_VDD_XI0/XI5/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI5/MM4 N_XI0/XI5/XI5/NET33_XI0/XI5/XI5/MM4_d
+ N_XI0/XI5/XI5/NET34_XI0/XI5/XI5/MM4_g N_VDD_XI0/XI5/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI5/MM10 N_XI0/XI5/XI5/NET35_XI0/XI5/XI5/MM10_d
+ N_XI0/XI5/XI5/NET36_XI0/XI5/XI5/MM10_g N_VDD_XI0/XI5/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI5/MM11 N_XI0/XI5/XI5/NET36_XI0/XI5/XI5/MM11_d
+ N_XI0/XI5/XI5/NET35_XI0/XI5/XI5/MM11_g N_VDD_XI0/XI5/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI6/MM2 N_XI0/XI5/XI6/NET34_XI0/XI5/XI6/MM2_d
+ N_XI0/XI5/XI6/NET33_XI0/XI5/XI6/MM2_g N_VSS_XI0/XI5/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI6/MM3 N_XI0/XI5/XI6/NET33_XI0/XI5/XI6/MM3_d N_WL<6>_XI0/XI5/XI6/MM3_g
+ N_BLN<9>_XI0/XI5/XI6/MM3_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI6/MM0 N_XI0/XI5/XI6/NET34_XI0/XI5/XI6/MM0_d N_WL<6>_XI0/XI5/XI6/MM0_g
+ N_BL<9>_XI0/XI5/XI6/MM0_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI6/MM1 N_XI0/XI5/XI6/NET33_XI0/XI5/XI6/MM1_d
+ N_XI0/XI5/XI6/NET34_XI0/XI5/XI6/MM1_g N_VSS_XI0/XI5/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI6/MM9 N_XI0/XI5/XI6/NET36_XI0/XI5/XI6/MM9_d N_WL<7>_XI0/XI5/XI6/MM9_g
+ N_BL<9>_XI0/XI5/XI6/MM9_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI6/MM6 N_XI0/XI5/XI6/NET35_XI0/XI5/XI6/MM6_d
+ N_XI0/XI5/XI6/NET36_XI0/XI5/XI6/MM6_g N_VSS_XI0/XI5/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI6/MM7 N_XI0/XI5/XI6/NET36_XI0/XI5/XI6/MM7_d
+ N_XI0/XI5/XI6/NET35_XI0/XI5/XI6/MM7_g N_VSS_XI0/XI5/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI6/MM8 N_XI0/XI5/XI6/NET35_XI0/XI5/XI6/MM8_d N_WL<7>_XI0/XI5/XI6/MM8_g
+ N_BLN<9>_XI0/XI5/XI6/MM8_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI6/MM5 N_XI0/XI5/XI6/NET34_XI0/XI5/XI6/MM5_d
+ N_XI0/XI5/XI6/NET33_XI0/XI5/XI6/MM5_g N_VDD_XI0/XI5/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI6/MM4 N_XI0/XI5/XI6/NET33_XI0/XI5/XI6/MM4_d
+ N_XI0/XI5/XI6/NET34_XI0/XI5/XI6/MM4_g N_VDD_XI0/XI5/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI6/MM10 N_XI0/XI5/XI6/NET35_XI0/XI5/XI6/MM10_d
+ N_XI0/XI5/XI6/NET36_XI0/XI5/XI6/MM10_g N_VDD_XI0/XI5/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI6/MM11 N_XI0/XI5/XI6/NET36_XI0/XI5/XI6/MM11_d
+ N_XI0/XI5/XI6/NET35_XI0/XI5/XI6/MM11_g N_VDD_XI0/XI5/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI7/MM2 N_XI0/XI5/XI7/NET34_XI0/XI5/XI7/MM2_d
+ N_XI0/XI5/XI7/NET33_XI0/XI5/XI7/MM2_g N_VSS_XI0/XI5/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI7/MM3 N_XI0/XI5/XI7/NET33_XI0/XI5/XI7/MM3_d N_WL<6>_XI0/XI5/XI7/MM3_g
+ N_BLN<8>_XI0/XI5/XI7/MM3_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI7/MM0 N_XI0/XI5/XI7/NET34_XI0/XI5/XI7/MM0_d N_WL<6>_XI0/XI5/XI7/MM0_g
+ N_BL<8>_XI0/XI5/XI7/MM0_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI7/MM1 N_XI0/XI5/XI7/NET33_XI0/XI5/XI7/MM1_d
+ N_XI0/XI5/XI7/NET34_XI0/XI5/XI7/MM1_g N_VSS_XI0/XI5/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI7/MM9 N_XI0/XI5/XI7/NET36_XI0/XI5/XI7/MM9_d N_WL<7>_XI0/XI5/XI7/MM9_g
+ N_BL<8>_XI0/XI5/XI7/MM9_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI7/MM6 N_XI0/XI5/XI7/NET35_XI0/XI5/XI7/MM6_d
+ N_XI0/XI5/XI7/NET36_XI0/XI5/XI7/MM6_g N_VSS_XI0/XI5/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI7/MM7 N_XI0/XI5/XI7/NET36_XI0/XI5/XI7/MM7_d
+ N_XI0/XI5/XI7/NET35_XI0/XI5/XI7/MM7_g N_VSS_XI0/XI5/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI7/MM8 N_XI0/XI5/XI7/NET35_XI0/XI5/XI7/MM8_d N_WL<7>_XI0/XI5/XI7/MM8_g
+ N_BLN<8>_XI0/XI5/XI7/MM8_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI7/MM5 N_XI0/XI5/XI7/NET34_XI0/XI5/XI7/MM5_d
+ N_XI0/XI5/XI7/NET33_XI0/XI5/XI7/MM5_g N_VDD_XI0/XI5/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI7/MM4 N_XI0/XI5/XI7/NET33_XI0/XI5/XI7/MM4_d
+ N_XI0/XI5/XI7/NET34_XI0/XI5/XI7/MM4_g N_VDD_XI0/XI5/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI7/MM10 N_XI0/XI5/XI7/NET35_XI0/XI5/XI7/MM10_d
+ N_XI0/XI5/XI7/NET36_XI0/XI5/XI7/MM10_g N_VDD_XI0/XI5/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI7/MM11 N_XI0/XI5/XI7/NET36_XI0/XI5/XI7/MM11_d
+ N_XI0/XI5/XI7/NET35_XI0/XI5/XI7/MM11_g N_VDD_XI0/XI5/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI8/MM2 N_XI0/XI5/XI8/NET34_XI0/XI5/XI8/MM2_d
+ N_XI0/XI5/XI8/NET33_XI0/XI5/XI8/MM2_g N_VSS_XI0/XI5/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI8/MM3 N_XI0/XI5/XI8/NET33_XI0/XI5/XI8/MM3_d N_WL<6>_XI0/XI5/XI8/MM3_g
+ N_BLN<7>_XI0/XI5/XI8/MM3_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI8/MM0 N_XI0/XI5/XI8/NET34_XI0/XI5/XI8/MM0_d N_WL<6>_XI0/XI5/XI8/MM0_g
+ N_BL<7>_XI0/XI5/XI8/MM0_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI8/MM1 N_XI0/XI5/XI8/NET33_XI0/XI5/XI8/MM1_d
+ N_XI0/XI5/XI8/NET34_XI0/XI5/XI8/MM1_g N_VSS_XI0/XI5/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI8/MM9 N_XI0/XI5/XI8/NET36_XI0/XI5/XI8/MM9_d N_WL<7>_XI0/XI5/XI8/MM9_g
+ N_BL<7>_XI0/XI5/XI8/MM9_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI8/MM6 N_XI0/XI5/XI8/NET35_XI0/XI5/XI8/MM6_d
+ N_XI0/XI5/XI8/NET36_XI0/XI5/XI8/MM6_g N_VSS_XI0/XI5/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI8/MM7 N_XI0/XI5/XI8/NET36_XI0/XI5/XI8/MM7_d
+ N_XI0/XI5/XI8/NET35_XI0/XI5/XI8/MM7_g N_VSS_XI0/XI5/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI8/MM8 N_XI0/XI5/XI8/NET35_XI0/XI5/XI8/MM8_d N_WL<7>_XI0/XI5/XI8/MM8_g
+ N_BLN<7>_XI0/XI5/XI8/MM8_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI8/MM5 N_XI0/XI5/XI8/NET34_XI0/XI5/XI8/MM5_d
+ N_XI0/XI5/XI8/NET33_XI0/XI5/XI8/MM5_g N_VDD_XI0/XI5/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI8/MM4 N_XI0/XI5/XI8/NET33_XI0/XI5/XI8/MM4_d
+ N_XI0/XI5/XI8/NET34_XI0/XI5/XI8/MM4_g N_VDD_XI0/XI5/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI8/MM10 N_XI0/XI5/XI8/NET35_XI0/XI5/XI8/MM10_d
+ N_XI0/XI5/XI8/NET36_XI0/XI5/XI8/MM10_g N_VDD_XI0/XI5/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI8/MM11 N_XI0/XI5/XI8/NET36_XI0/XI5/XI8/MM11_d
+ N_XI0/XI5/XI8/NET35_XI0/XI5/XI8/MM11_g N_VDD_XI0/XI5/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI9/MM2 N_XI0/XI5/XI9/NET34_XI0/XI5/XI9/MM2_d
+ N_XI0/XI5/XI9/NET33_XI0/XI5/XI9/MM2_g N_VSS_XI0/XI5/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI9/MM3 N_XI0/XI5/XI9/NET33_XI0/XI5/XI9/MM3_d N_WL<6>_XI0/XI5/XI9/MM3_g
+ N_BLN<6>_XI0/XI5/XI9/MM3_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI9/MM0 N_XI0/XI5/XI9/NET34_XI0/XI5/XI9/MM0_d N_WL<6>_XI0/XI5/XI9/MM0_g
+ N_BL<6>_XI0/XI5/XI9/MM0_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI9/MM1 N_XI0/XI5/XI9/NET33_XI0/XI5/XI9/MM1_d
+ N_XI0/XI5/XI9/NET34_XI0/XI5/XI9/MM1_g N_VSS_XI0/XI5/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI9/MM9 N_XI0/XI5/XI9/NET36_XI0/XI5/XI9/MM9_d N_WL<7>_XI0/XI5/XI9/MM9_g
+ N_BL<6>_XI0/XI5/XI9/MM9_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI9/MM6 N_XI0/XI5/XI9/NET35_XI0/XI5/XI9/MM6_d
+ N_XI0/XI5/XI9/NET36_XI0/XI5/XI9/MM6_g N_VSS_XI0/XI5/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI9/MM7 N_XI0/XI5/XI9/NET36_XI0/XI5/XI9/MM7_d
+ N_XI0/XI5/XI9/NET35_XI0/XI5/XI9/MM7_g N_VSS_XI0/XI5/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI9/MM8 N_XI0/XI5/XI9/NET35_XI0/XI5/XI9/MM8_d N_WL<7>_XI0/XI5/XI9/MM8_g
+ N_BLN<6>_XI0/XI5/XI9/MM8_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI5/XI9/MM5 N_XI0/XI5/XI9/NET34_XI0/XI5/XI9/MM5_d
+ N_XI0/XI5/XI9/NET33_XI0/XI5/XI9/MM5_g N_VDD_XI0/XI5/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI9/MM4 N_XI0/XI5/XI9/NET33_XI0/XI5/XI9/MM4_d
+ N_XI0/XI5/XI9/NET34_XI0/XI5/XI9/MM4_g N_VDD_XI0/XI5/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI9/MM10 N_XI0/XI5/XI9/NET35_XI0/XI5/XI9/MM10_d
+ N_XI0/XI5/XI9/NET36_XI0/XI5/XI9/MM10_g N_VDD_XI0/XI5/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI9/MM11 N_XI0/XI5/XI9/NET36_XI0/XI5/XI9/MM11_d
+ N_XI0/XI5/XI9/NET35_XI0/XI5/XI9/MM11_g N_VDD_XI0/XI5/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI10/MM2 N_XI0/XI5/XI10/NET34_XI0/XI5/XI10/MM2_d
+ N_XI0/XI5/XI10/NET33_XI0/XI5/XI10/MM2_g N_VSS_XI0/XI5/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM3 N_XI0/XI5/XI10/NET33_XI0/XI5/XI10/MM3_d
+ N_WL<6>_XI0/XI5/XI10/MM3_g N_BLN<5>_XI0/XI5/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM0 N_XI0/XI5/XI10/NET34_XI0/XI5/XI10/MM0_d
+ N_WL<6>_XI0/XI5/XI10/MM0_g N_BL<5>_XI0/XI5/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM1 N_XI0/XI5/XI10/NET33_XI0/XI5/XI10/MM1_d
+ N_XI0/XI5/XI10/NET34_XI0/XI5/XI10/MM1_g N_VSS_XI0/XI5/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM9 N_XI0/XI5/XI10/NET36_XI0/XI5/XI10/MM9_d
+ N_WL<7>_XI0/XI5/XI10/MM9_g N_BL<5>_XI0/XI5/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM6 N_XI0/XI5/XI10/NET35_XI0/XI5/XI10/MM6_d
+ N_XI0/XI5/XI10/NET36_XI0/XI5/XI10/MM6_g N_VSS_XI0/XI5/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM7 N_XI0/XI5/XI10/NET36_XI0/XI5/XI10/MM7_d
+ N_XI0/XI5/XI10/NET35_XI0/XI5/XI10/MM7_g N_VSS_XI0/XI5/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM8 N_XI0/XI5/XI10/NET35_XI0/XI5/XI10/MM8_d
+ N_WL<7>_XI0/XI5/XI10/MM8_g N_BLN<5>_XI0/XI5/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI10/MM5 N_XI0/XI5/XI10/NET34_XI0/XI5/XI10/MM5_d
+ N_XI0/XI5/XI10/NET33_XI0/XI5/XI10/MM5_g N_VDD_XI0/XI5/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI10/MM4 N_XI0/XI5/XI10/NET33_XI0/XI5/XI10/MM4_d
+ N_XI0/XI5/XI10/NET34_XI0/XI5/XI10/MM4_g N_VDD_XI0/XI5/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI10/MM10 N_XI0/XI5/XI10/NET35_XI0/XI5/XI10/MM10_d
+ N_XI0/XI5/XI10/NET36_XI0/XI5/XI10/MM10_g N_VDD_XI0/XI5/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI10/MM11 N_XI0/XI5/XI10/NET36_XI0/XI5/XI10/MM11_d
+ N_XI0/XI5/XI10/NET35_XI0/XI5/XI10/MM11_g N_VDD_XI0/XI5/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI11/MM2 N_XI0/XI5/XI11/NET34_XI0/XI5/XI11/MM2_d
+ N_XI0/XI5/XI11/NET33_XI0/XI5/XI11/MM2_g N_VSS_XI0/XI5/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM3 N_XI0/XI5/XI11/NET33_XI0/XI5/XI11/MM3_d
+ N_WL<6>_XI0/XI5/XI11/MM3_g N_BLN<4>_XI0/XI5/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM0 N_XI0/XI5/XI11/NET34_XI0/XI5/XI11/MM0_d
+ N_WL<6>_XI0/XI5/XI11/MM0_g N_BL<4>_XI0/XI5/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM1 N_XI0/XI5/XI11/NET33_XI0/XI5/XI11/MM1_d
+ N_XI0/XI5/XI11/NET34_XI0/XI5/XI11/MM1_g N_VSS_XI0/XI5/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM9 N_XI0/XI5/XI11/NET36_XI0/XI5/XI11/MM9_d
+ N_WL<7>_XI0/XI5/XI11/MM9_g N_BL<4>_XI0/XI5/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM6 N_XI0/XI5/XI11/NET35_XI0/XI5/XI11/MM6_d
+ N_XI0/XI5/XI11/NET36_XI0/XI5/XI11/MM6_g N_VSS_XI0/XI5/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM7 N_XI0/XI5/XI11/NET36_XI0/XI5/XI11/MM7_d
+ N_XI0/XI5/XI11/NET35_XI0/XI5/XI11/MM7_g N_VSS_XI0/XI5/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM8 N_XI0/XI5/XI11/NET35_XI0/XI5/XI11/MM8_d
+ N_WL<7>_XI0/XI5/XI11/MM8_g N_BLN<4>_XI0/XI5/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI11/MM5 N_XI0/XI5/XI11/NET34_XI0/XI5/XI11/MM5_d
+ N_XI0/XI5/XI11/NET33_XI0/XI5/XI11/MM5_g N_VDD_XI0/XI5/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI11/MM4 N_XI0/XI5/XI11/NET33_XI0/XI5/XI11/MM4_d
+ N_XI0/XI5/XI11/NET34_XI0/XI5/XI11/MM4_g N_VDD_XI0/XI5/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI11/MM10 N_XI0/XI5/XI11/NET35_XI0/XI5/XI11/MM10_d
+ N_XI0/XI5/XI11/NET36_XI0/XI5/XI11/MM10_g N_VDD_XI0/XI5/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI11/MM11 N_XI0/XI5/XI11/NET36_XI0/XI5/XI11/MM11_d
+ N_XI0/XI5/XI11/NET35_XI0/XI5/XI11/MM11_g N_VDD_XI0/XI5/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI12/MM2 N_XI0/XI5/XI12/NET34_XI0/XI5/XI12/MM2_d
+ N_XI0/XI5/XI12/NET33_XI0/XI5/XI12/MM2_g N_VSS_XI0/XI5/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM3 N_XI0/XI5/XI12/NET33_XI0/XI5/XI12/MM3_d
+ N_WL<6>_XI0/XI5/XI12/MM3_g N_BLN<3>_XI0/XI5/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM0 N_XI0/XI5/XI12/NET34_XI0/XI5/XI12/MM0_d
+ N_WL<6>_XI0/XI5/XI12/MM0_g N_BL<3>_XI0/XI5/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM1 N_XI0/XI5/XI12/NET33_XI0/XI5/XI12/MM1_d
+ N_XI0/XI5/XI12/NET34_XI0/XI5/XI12/MM1_g N_VSS_XI0/XI5/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM9 N_XI0/XI5/XI12/NET36_XI0/XI5/XI12/MM9_d
+ N_WL<7>_XI0/XI5/XI12/MM9_g N_BL<3>_XI0/XI5/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM6 N_XI0/XI5/XI12/NET35_XI0/XI5/XI12/MM6_d
+ N_XI0/XI5/XI12/NET36_XI0/XI5/XI12/MM6_g N_VSS_XI0/XI5/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM7 N_XI0/XI5/XI12/NET36_XI0/XI5/XI12/MM7_d
+ N_XI0/XI5/XI12/NET35_XI0/XI5/XI12/MM7_g N_VSS_XI0/XI5/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM8 N_XI0/XI5/XI12/NET35_XI0/XI5/XI12/MM8_d
+ N_WL<7>_XI0/XI5/XI12/MM8_g N_BLN<3>_XI0/XI5/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI12/MM5 N_XI0/XI5/XI12/NET34_XI0/XI5/XI12/MM5_d
+ N_XI0/XI5/XI12/NET33_XI0/XI5/XI12/MM5_g N_VDD_XI0/XI5/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI12/MM4 N_XI0/XI5/XI12/NET33_XI0/XI5/XI12/MM4_d
+ N_XI0/XI5/XI12/NET34_XI0/XI5/XI12/MM4_g N_VDD_XI0/XI5/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI12/MM10 N_XI0/XI5/XI12/NET35_XI0/XI5/XI12/MM10_d
+ N_XI0/XI5/XI12/NET36_XI0/XI5/XI12/MM10_g N_VDD_XI0/XI5/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI12/MM11 N_XI0/XI5/XI12/NET36_XI0/XI5/XI12/MM11_d
+ N_XI0/XI5/XI12/NET35_XI0/XI5/XI12/MM11_g N_VDD_XI0/XI5/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI13/MM2 N_XI0/XI5/XI13/NET34_XI0/XI5/XI13/MM2_d
+ N_XI0/XI5/XI13/NET33_XI0/XI5/XI13/MM2_g N_VSS_XI0/XI5/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM3 N_XI0/XI5/XI13/NET33_XI0/XI5/XI13/MM3_d
+ N_WL<6>_XI0/XI5/XI13/MM3_g N_BLN<2>_XI0/XI5/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM0 N_XI0/XI5/XI13/NET34_XI0/XI5/XI13/MM0_d
+ N_WL<6>_XI0/XI5/XI13/MM0_g N_BL<2>_XI0/XI5/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM1 N_XI0/XI5/XI13/NET33_XI0/XI5/XI13/MM1_d
+ N_XI0/XI5/XI13/NET34_XI0/XI5/XI13/MM1_g N_VSS_XI0/XI5/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM9 N_XI0/XI5/XI13/NET36_XI0/XI5/XI13/MM9_d
+ N_WL<7>_XI0/XI5/XI13/MM9_g N_BL<2>_XI0/XI5/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM6 N_XI0/XI5/XI13/NET35_XI0/XI5/XI13/MM6_d
+ N_XI0/XI5/XI13/NET36_XI0/XI5/XI13/MM6_g N_VSS_XI0/XI5/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM7 N_XI0/XI5/XI13/NET36_XI0/XI5/XI13/MM7_d
+ N_XI0/XI5/XI13/NET35_XI0/XI5/XI13/MM7_g N_VSS_XI0/XI5/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM8 N_XI0/XI5/XI13/NET35_XI0/XI5/XI13/MM8_d
+ N_WL<7>_XI0/XI5/XI13/MM8_g N_BLN<2>_XI0/XI5/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI13/MM5 N_XI0/XI5/XI13/NET34_XI0/XI5/XI13/MM5_d
+ N_XI0/XI5/XI13/NET33_XI0/XI5/XI13/MM5_g N_VDD_XI0/XI5/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI13/MM4 N_XI0/XI5/XI13/NET33_XI0/XI5/XI13/MM4_d
+ N_XI0/XI5/XI13/NET34_XI0/XI5/XI13/MM4_g N_VDD_XI0/XI5/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI13/MM10 N_XI0/XI5/XI13/NET35_XI0/XI5/XI13/MM10_d
+ N_XI0/XI5/XI13/NET36_XI0/XI5/XI13/MM10_g N_VDD_XI0/XI5/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI13/MM11 N_XI0/XI5/XI13/NET36_XI0/XI5/XI13/MM11_d
+ N_XI0/XI5/XI13/NET35_XI0/XI5/XI13/MM11_g N_VDD_XI0/XI5/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI14/MM2 N_XI0/XI5/XI14/NET34_XI0/XI5/XI14/MM2_d
+ N_XI0/XI5/XI14/NET33_XI0/XI5/XI14/MM2_g N_VSS_XI0/XI5/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM3 N_XI0/XI5/XI14/NET33_XI0/XI5/XI14/MM3_d
+ N_WL<6>_XI0/XI5/XI14/MM3_g N_BLN<1>_XI0/XI5/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM0 N_XI0/XI5/XI14/NET34_XI0/XI5/XI14/MM0_d
+ N_WL<6>_XI0/XI5/XI14/MM0_g N_BL<1>_XI0/XI5/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM1 N_XI0/XI5/XI14/NET33_XI0/XI5/XI14/MM1_d
+ N_XI0/XI5/XI14/NET34_XI0/XI5/XI14/MM1_g N_VSS_XI0/XI5/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM9 N_XI0/XI5/XI14/NET36_XI0/XI5/XI14/MM9_d
+ N_WL<7>_XI0/XI5/XI14/MM9_g N_BL<1>_XI0/XI5/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM6 N_XI0/XI5/XI14/NET35_XI0/XI5/XI14/MM6_d
+ N_XI0/XI5/XI14/NET36_XI0/XI5/XI14/MM6_g N_VSS_XI0/XI5/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM7 N_XI0/XI5/XI14/NET36_XI0/XI5/XI14/MM7_d
+ N_XI0/XI5/XI14/NET35_XI0/XI5/XI14/MM7_g N_VSS_XI0/XI5/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM8 N_XI0/XI5/XI14/NET35_XI0/XI5/XI14/MM8_d
+ N_WL<7>_XI0/XI5/XI14/MM8_g N_BLN<1>_XI0/XI5/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI14/MM5 N_XI0/XI5/XI14/NET34_XI0/XI5/XI14/MM5_d
+ N_XI0/XI5/XI14/NET33_XI0/XI5/XI14/MM5_g N_VDD_XI0/XI5/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI14/MM4 N_XI0/XI5/XI14/NET33_XI0/XI5/XI14/MM4_d
+ N_XI0/XI5/XI14/NET34_XI0/XI5/XI14/MM4_g N_VDD_XI0/XI5/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI14/MM10 N_XI0/XI5/XI14/NET35_XI0/XI5/XI14/MM10_d
+ N_XI0/XI5/XI14/NET36_XI0/XI5/XI14/MM10_g N_VDD_XI0/XI5/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI14/MM11 N_XI0/XI5/XI14/NET36_XI0/XI5/XI14/MM11_d
+ N_XI0/XI5/XI14/NET35_XI0/XI5/XI14/MM11_g N_VDD_XI0/XI5/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI15/MM2 N_XI0/XI5/XI15/NET34_XI0/XI5/XI15/MM2_d
+ N_XI0/XI5/XI15/NET33_XI0/XI5/XI15/MM2_g N_VSS_XI0/XI5/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM3 N_XI0/XI5/XI15/NET33_XI0/XI5/XI15/MM3_d
+ N_WL<6>_XI0/XI5/XI15/MM3_g N_BLN<0>_XI0/XI5/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM0 N_XI0/XI5/XI15/NET34_XI0/XI5/XI15/MM0_d
+ N_WL<6>_XI0/XI5/XI15/MM0_g N_BL<0>_XI0/XI5/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM1 N_XI0/XI5/XI15/NET33_XI0/XI5/XI15/MM1_d
+ N_XI0/XI5/XI15/NET34_XI0/XI5/XI15/MM1_g N_VSS_XI0/XI5/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM9 N_XI0/XI5/XI15/NET36_XI0/XI5/XI15/MM9_d
+ N_WL<7>_XI0/XI5/XI15/MM9_g N_BL<0>_XI0/XI5/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM6 N_XI0/XI5/XI15/NET35_XI0/XI5/XI15/MM6_d
+ N_XI0/XI5/XI15/NET36_XI0/XI5/XI15/MM6_g N_VSS_XI0/XI5/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM7 N_XI0/XI5/XI15/NET36_XI0/XI5/XI15/MM7_d
+ N_XI0/XI5/XI15/NET35_XI0/XI5/XI15/MM7_g N_VSS_XI0/XI5/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM8 N_XI0/XI5/XI15/NET35_XI0/XI5/XI15/MM8_d
+ N_WL<7>_XI0/XI5/XI15/MM8_g N_BLN<0>_XI0/XI5/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/XI15/MM5 N_XI0/XI5/XI15/NET34_XI0/XI5/XI15/MM5_d
+ N_XI0/XI5/XI15/NET33_XI0/XI5/XI15/MM5_g N_VDD_XI0/XI5/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI15/MM4 N_XI0/XI5/XI15/NET33_XI0/XI5/XI15/MM4_d
+ N_XI0/XI5/XI15/NET34_XI0/XI5/XI15/MM4_g N_VDD_XI0/XI5/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI15/MM10 N_XI0/XI5/XI15/NET35_XI0/XI5/XI15/MM10_d
+ N_XI0/XI5/XI15/NET36_XI0/XI5/XI15/MM10_g N_VDD_XI0/XI5/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/XI15/MM11 N_XI0/XI5/XI15/NET36_XI0/XI5/XI15/MM11_d
+ N_XI0/XI5/XI15/NET35_XI0/XI5/XI15/MM11_g N_VDD_XI0/XI5/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI0/MM2 N_XI0/XI6/XI0/NET34_XI0/XI6/XI0/MM2_d
+ N_XI0/XI6/XI0/NET33_XI0/XI6/XI0/MM2_g N_VSS_XI0/XI6/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI0/MM3 N_XI0/XI6/XI0/NET33_XI0/XI6/XI0/MM3_d N_WL<8>_XI0/XI6/XI0/MM3_g
+ N_BLN<15>_XI0/XI6/XI0/MM3_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI0/MM0 N_XI0/XI6/XI0/NET34_XI0/XI6/XI0/MM0_d N_WL<8>_XI0/XI6/XI0/MM0_g
+ N_BL<15>_XI0/XI6/XI0/MM0_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI0/MM1 N_XI0/XI6/XI0/NET33_XI0/XI6/XI0/MM1_d
+ N_XI0/XI6/XI0/NET34_XI0/XI6/XI0/MM1_g N_VSS_XI0/XI6/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI0/MM9 N_XI0/XI6/XI0/NET36_XI0/XI6/XI0/MM9_d N_WL<9>_XI0/XI6/XI0/MM9_g
+ N_BL<15>_XI0/XI6/XI0/MM9_s N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI0/MM6 N_XI0/XI6/XI0/NET35_XI0/XI6/XI0/MM6_d
+ N_XI0/XI6/XI0/NET36_XI0/XI6/XI0/MM6_g N_VSS_XI0/XI6/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI0/MM7 N_XI0/XI6/XI0/NET36_XI0/XI6/XI0/MM7_d
+ N_XI0/XI6/XI0/NET35_XI0/XI6/XI0/MM7_g N_VSS_XI0/XI6/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI0/MM8 N_XI0/XI6/XI0/NET35_XI0/XI6/XI0/MM8_d N_WL<9>_XI0/XI6/XI0/MM8_g
+ N_BLN<15>_XI0/XI6/XI0/MM8_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI0/MM5 N_XI0/XI6/XI0/NET34_XI0/XI6/XI0/MM5_d
+ N_XI0/XI6/XI0/NET33_XI0/XI6/XI0/MM5_g N_VDD_XI0/XI6/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI0/MM4 N_XI0/XI6/XI0/NET33_XI0/XI6/XI0/MM4_d
+ N_XI0/XI6/XI0/NET34_XI0/XI6/XI0/MM4_g N_VDD_XI0/XI6/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI0/MM10 N_XI0/XI6/XI0/NET35_XI0/XI6/XI0/MM10_d
+ N_XI0/XI6/XI0/NET36_XI0/XI6/XI0/MM10_g N_VDD_XI0/XI6/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI0/MM11 N_XI0/XI6/XI0/NET36_XI0/XI6/XI0/MM11_d
+ N_XI0/XI6/XI0/NET35_XI0/XI6/XI0/MM11_g N_VDD_XI0/XI6/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI1/MM2 N_XI0/XI6/XI1/NET34_XI0/XI6/XI1/MM2_d
+ N_XI0/XI6/XI1/NET33_XI0/XI6/XI1/MM2_g N_VSS_XI0/XI6/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI1/MM3 N_XI0/XI6/XI1/NET33_XI0/XI6/XI1/MM3_d N_WL<8>_XI0/XI6/XI1/MM3_g
+ N_BLN<14>_XI0/XI6/XI1/MM3_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI1/MM0 N_XI0/XI6/XI1/NET34_XI0/XI6/XI1/MM0_d N_WL<8>_XI0/XI6/XI1/MM0_g
+ N_BL<14>_XI0/XI6/XI1/MM0_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI1/MM1 N_XI0/XI6/XI1/NET33_XI0/XI6/XI1/MM1_d
+ N_XI0/XI6/XI1/NET34_XI0/XI6/XI1/MM1_g N_VSS_XI0/XI6/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI1/MM9 N_XI0/XI6/XI1/NET36_XI0/XI6/XI1/MM9_d N_WL<9>_XI0/XI6/XI1/MM9_g
+ N_BL<14>_XI0/XI6/XI1/MM9_s N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI1/MM6 N_XI0/XI6/XI1/NET35_XI0/XI6/XI1/MM6_d
+ N_XI0/XI6/XI1/NET36_XI0/XI6/XI1/MM6_g N_VSS_XI0/XI6/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI1/MM7 N_XI0/XI6/XI1/NET36_XI0/XI6/XI1/MM7_d
+ N_XI0/XI6/XI1/NET35_XI0/XI6/XI1/MM7_g N_VSS_XI0/XI6/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI1/MM8 N_XI0/XI6/XI1/NET35_XI0/XI6/XI1/MM8_d N_WL<9>_XI0/XI6/XI1/MM8_g
+ N_BLN<14>_XI0/XI6/XI1/MM8_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI1/MM5 N_XI0/XI6/XI1/NET34_XI0/XI6/XI1/MM5_d
+ N_XI0/XI6/XI1/NET33_XI0/XI6/XI1/MM5_g N_VDD_XI0/XI6/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI1/MM4 N_XI0/XI6/XI1/NET33_XI0/XI6/XI1/MM4_d
+ N_XI0/XI6/XI1/NET34_XI0/XI6/XI1/MM4_g N_VDD_XI0/XI6/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI1/MM10 N_XI0/XI6/XI1/NET35_XI0/XI6/XI1/MM10_d
+ N_XI0/XI6/XI1/NET36_XI0/XI6/XI1/MM10_g N_VDD_XI0/XI6/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI1/MM11 N_XI0/XI6/XI1/NET36_XI0/XI6/XI1/MM11_d
+ N_XI0/XI6/XI1/NET35_XI0/XI6/XI1/MM11_g N_VDD_XI0/XI6/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI2/MM2 N_XI0/XI6/XI2/NET34_XI0/XI6/XI2/MM2_d
+ N_XI0/XI6/XI2/NET33_XI0/XI6/XI2/MM2_g N_VSS_XI0/XI6/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI2/MM3 N_XI0/XI6/XI2/NET33_XI0/XI6/XI2/MM3_d N_WL<8>_XI0/XI6/XI2/MM3_g
+ N_BLN<13>_XI0/XI6/XI2/MM3_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI2/MM0 N_XI0/XI6/XI2/NET34_XI0/XI6/XI2/MM0_d N_WL<8>_XI0/XI6/XI2/MM0_g
+ N_BL<13>_XI0/XI6/XI2/MM0_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI2/MM1 N_XI0/XI6/XI2/NET33_XI0/XI6/XI2/MM1_d
+ N_XI0/XI6/XI2/NET34_XI0/XI6/XI2/MM1_g N_VSS_XI0/XI6/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI2/MM9 N_XI0/XI6/XI2/NET36_XI0/XI6/XI2/MM9_d N_WL<9>_XI0/XI6/XI2/MM9_g
+ N_BL<13>_XI0/XI6/XI2/MM9_s N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI2/MM6 N_XI0/XI6/XI2/NET35_XI0/XI6/XI2/MM6_d
+ N_XI0/XI6/XI2/NET36_XI0/XI6/XI2/MM6_g N_VSS_XI0/XI6/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI2/MM7 N_XI0/XI6/XI2/NET36_XI0/XI6/XI2/MM7_d
+ N_XI0/XI6/XI2/NET35_XI0/XI6/XI2/MM7_g N_VSS_XI0/XI6/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI2/MM8 N_XI0/XI6/XI2/NET35_XI0/XI6/XI2/MM8_d N_WL<9>_XI0/XI6/XI2/MM8_g
+ N_BLN<13>_XI0/XI6/XI2/MM8_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI2/MM5 N_XI0/XI6/XI2/NET34_XI0/XI6/XI2/MM5_d
+ N_XI0/XI6/XI2/NET33_XI0/XI6/XI2/MM5_g N_VDD_XI0/XI6/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI2/MM4 N_XI0/XI6/XI2/NET33_XI0/XI6/XI2/MM4_d
+ N_XI0/XI6/XI2/NET34_XI0/XI6/XI2/MM4_g N_VDD_XI0/XI6/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI2/MM10 N_XI0/XI6/XI2/NET35_XI0/XI6/XI2/MM10_d
+ N_XI0/XI6/XI2/NET36_XI0/XI6/XI2/MM10_g N_VDD_XI0/XI6/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI2/MM11 N_XI0/XI6/XI2/NET36_XI0/XI6/XI2/MM11_d
+ N_XI0/XI6/XI2/NET35_XI0/XI6/XI2/MM11_g N_VDD_XI0/XI6/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI3/MM2 N_XI0/XI6/XI3/NET34_XI0/XI6/XI3/MM2_d
+ N_XI0/XI6/XI3/NET33_XI0/XI6/XI3/MM2_g N_VSS_XI0/XI6/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI3/MM3 N_XI0/XI6/XI3/NET33_XI0/XI6/XI3/MM3_d N_WL<8>_XI0/XI6/XI3/MM3_g
+ N_BLN<12>_XI0/XI6/XI3/MM3_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI3/MM0 N_XI0/XI6/XI3/NET34_XI0/XI6/XI3/MM0_d N_WL<8>_XI0/XI6/XI3/MM0_g
+ N_BL<12>_XI0/XI6/XI3/MM0_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI3/MM1 N_XI0/XI6/XI3/NET33_XI0/XI6/XI3/MM1_d
+ N_XI0/XI6/XI3/NET34_XI0/XI6/XI3/MM1_g N_VSS_XI0/XI6/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI3/MM9 N_XI0/XI6/XI3/NET36_XI0/XI6/XI3/MM9_d N_WL<9>_XI0/XI6/XI3/MM9_g
+ N_BL<12>_XI0/XI6/XI3/MM9_s N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI3/MM6 N_XI0/XI6/XI3/NET35_XI0/XI6/XI3/MM6_d
+ N_XI0/XI6/XI3/NET36_XI0/XI6/XI3/MM6_g N_VSS_XI0/XI6/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI3/MM7 N_XI0/XI6/XI3/NET36_XI0/XI6/XI3/MM7_d
+ N_XI0/XI6/XI3/NET35_XI0/XI6/XI3/MM7_g N_VSS_XI0/XI6/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI3/MM8 N_XI0/XI6/XI3/NET35_XI0/XI6/XI3/MM8_d N_WL<9>_XI0/XI6/XI3/MM8_g
+ N_BLN<12>_XI0/XI6/XI3/MM8_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI3/MM5 N_XI0/XI6/XI3/NET34_XI0/XI6/XI3/MM5_d
+ N_XI0/XI6/XI3/NET33_XI0/XI6/XI3/MM5_g N_VDD_XI0/XI6/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI3/MM4 N_XI0/XI6/XI3/NET33_XI0/XI6/XI3/MM4_d
+ N_XI0/XI6/XI3/NET34_XI0/XI6/XI3/MM4_g N_VDD_XI0/XI6/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI3/MM10 N_XI0/XI6/XI3/NET35_XI0/XI6/XI3/MM10_d
+ N_XI0/XI6/XI3/NET36_XI0/XI6/XI3/MM10_g N_VDD_XI0/XI6/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI3/MM11 N_XI0/XI6/XI3/NET36_XI0/XI6/XI3/MM11_d
+ N_XI0/XI6/XI3/NET35_XI0/XI6/XI3/MM11_g N_VDD_XI0/XI6/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI4/MM2 N_XI0/XI6/XI4/NET34_XI0/XI6/XI4/MM2_d
+ N_XI0/XI6/XI4/NET33_XI0/XI6/XI4/MM2_g N_VSS_XI0/XI6/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI4/MM3 N_XI0/XI6/XI4/NET33_XI0/XI6/XI4/MM3_d N_WL<8>_XI0/XI6/XI4/MM3_g
+ N_BLN<11>_XI0/XI6/XI4/MM3_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI4/MM0 N_XI0/XI6/XI4/NET34_XI0/XI6/XI4/MM0_d N_WL<8>_XI0/XI6/XI4/MM0_g
+ N_BL<11>_XI0/XI6/XI4/MM0_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI4/MM1 N_XI0/XI6/XI4/NET33_XI0/XI6/XI4/MM1_d
+ N_XI0/XI6/XI4/NET34_XI0/XI6/XI4/MM1_g N_VSS_XI0/XI6/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI4/MM9 N_XI0/XI6/XI4/NET36_XI0/XI6/XI4/MM9_d N_WL<9>_XI0/XI6/XI4/MM9_g
+ N_BL<11>_XI0/XI6/XI4/MM9_s N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI4/MM6 N_XI0/XI6/XI4/NET35_XI0/XI6/XI4/MM6_d
+ N_XI0/XI6/XI4/NET36_XI0/XI6/XI4/MM6_g N_VSS_XI0/XI6/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI4/MM7 N_XI0/XI6/XI4/NET36_XI0/XI6/XI4/MM7_d
+ N_XI0/XI6/XI4/NET35_XI0/XI6/XI4/MM7_g N_VSS_XI0/XI6/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI4/MM8 N_XI0/XI6/XI4/NET35_XI0/XI6/XI4/MM8_d N_WL<9>_XI0/XI6/XI4/MM8_g
+ N_BLN<11>_XI0/XI6/XI4/MM8_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI4/MM5 N_XI0/XI6/XI4/NET34_XI0/XI6/XI4/MM5_d
+ N_XI0/XI6/XI4/NET33_XI0/XI6/XI4/MM5_g N_VDD_XI0/XI6/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI4/MM4 N_XI0/XI6/XI4/NET33_XI0/XI6/XI4/MM4_d
+ N_XI0/XI6/XI4/NET34_XI0/XI6/XI4/MM4_g N_VDD_XI0/XI6/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI4/MM10 N_XI0/XI6/XI4/NET35_XI0/XI6/XI4/MM10_d
+ N_XI0/XI6/XI4/NET36_XI0/XI6/XI4/MM10_g N_VDD_XI0/XI6/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI4/MM11 N_XI0/XI6/XI4/NET36_XI0/XI6/XI4/MM11_d
+ N_XI0/XI6/XI4/NET35_XI0/XI6/XI4/MM11_g N_VDD_XI0/XI6/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI5/MM2 N_XI0/XI6/XI5/NET34_XI0/XI6/XI5/MM2_d
+ N_XI0/XI6/XI5/NET33_XI0/XI6/XI5/MM2_g N_VSS_XI0/XI6/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI5/MM3 N_XI0/XI6/XI5/NET33_XI0/XI6/XI5/MM3_d N_WL<8>_XI0/XI6/XI5/MM3_g
+ N_BLN<10>_XI0/XI6/XI5/MM3_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI5/MM0 N_XI0/XI6/XI5/NET34_XI0/XI6/XI5/MM0_d N_WL<8>_XI0/XI6/XI5/MM0_g
+ N_BL<10>_XI0/XI6/XI5/MM0_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI5/MM1 N_XI0/XI6/XI5/NET33_XI0/XI6/XI5/MM1_d
+ N_XI0/XI6/XI5/NET34_XI0/XI6/XI5/MM1_g N_VSS_XI0/XI6/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI5/MM9 N_XI0/XI6/XI5/NET36_XI0/XI6/XI5/MM9_d N_WL<9>_XI0/XI6/XI5/MM9_g
+ N_BL<10>_XI0/XI6/XI5/MM9_s N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI5/MM6 N_XI0/XI6/XI5/NET35_XI0/XI6/XI5/MM6_d
+ N_XI0/XI6/XI5/NET36_XI0/XI6/XI5/MM6_g N_VSS_XI0/XI6/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI5/MM7 N_XI0/XI6/XI5/NET36_XI0/XI6/XI5/MM7_d
+ N_XI0/XI6/XI5/NET35_XI0/XI6/XI5/MM7_g N_VSS_XI0/XI6/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI5/MM8 N_XI0/XI6/XI5/NET35_XI0/XI6/XI5/MM8_d N_WL<9>_XI0/XI6/XI5/MM8_g
+ N_BLN<10>_XI0/XI6/XI5/MM8_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI5/MM5 N_XI0/XI6/XI5/NET34_XI0/XI6/XI5/MM5_d
+ N_XI0/XI6/XI5/NET33_XI0/XI6/XI5/MM5_g N_VDD_XI0/XI6/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI5/MM4 N_XI0/XI6/XI5/NET33_XI0/XI6/XI5/MM4_d
+ N_XI0/XI6/XI5/NET34_XI0/XI6/XI5/MM4_g N_VDD_XI0/XI6/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI5/MM10 N_XI0/XI6/XI5/NET35_XI0/XI6/XI5/MM10_d
+ N_XI0/XI6/XI5/NET36_XI0/XI6/XI5/MM10_g N_VDD_XI0/XI6/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI5/MM11 N_XI0/XI6/XI5/NET36_XI0/XI6/XI5/MM11_d
+ N_XI0/XI6/XI5/NET35_XI0/XI6/XI5/MM11_g N_VDD_XI0/XI6/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI6/MM2 N_XI0/XI6/XI6/NET34_XI0/XI6/XI6/MM2_d
+ N_XI0/XI6/XI6/NET33_XI0/XI6/XI6/MM2_g N_VSS_XI0/XI6/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI6/MM3 N_XI0/XI6/XI6/NET33_XI0/XI6/XI6/MM3_d N_WL<8>_XI0/XI6/XI6/MM3_g
+ N_BLN<9>_XI0/XI6/XI6/MM3_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI6/MM0 N_XI0/XI6/XI6/NET34_XI0/XI6/XI6/MM0_d N_WL<8>_XI0/XI6/XI6/MM0_g
+ N_BL<9>_XI0/XI6/XI6/MM0_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI6/MM1 N_XI0/XI6/XI6/NET33_XI0/XI6/XI6/MM1_d
+ N_XI0/XI6/XI6/NET34_XI0/XI6/XI6/MM1_g N_VSS_XI0/XI6/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI6/MM9 N_XI0/XI6/XI6/NET36_XI0/XI6/XI6/MM9_d N_WL<9>_XI0/XI6/XI6/MM9_g
+ N_BL<9>_XI0/XI6/XI6/MM9_s N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI6/MM6 N_XI0/XI6/XI6/NET35_XI0/XI6/XI6/MM6_d
+ N_XI0/XI6/XI6/NET36_XI0/XI6/XI6/MM6_g N_VSS_XI0/XI6/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI6/MM7 N_XI0/XI6/XI6/NET36_XI0/XI6/XI6/MM7_d
+ N_XI0/XI6/XI6/NET35_XI0/XI6/XI6/MM7_g N_VSS_XI0/XI6/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI6/MM8 N_XI0/XI6/XI6/NET35_XI0/XI6/XI6/MM8_d N_WL<9>_XI0/XI6/XI6/MM8_g
+ N_BLN<9>_XI0/XI6/XI6/MM8_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI6/MM5 N_XI0/XI6/XI6/NET34_XI0/XI6/XI6/MM5_d
+ N_XI0/XI6/XI6/NET33_XI0/XI6/XI6/MM5_g N_VDD_XI0/XI6/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI6/MM4 N_XI0/XI6/XI6/NET33_XI0/XI6/XI6/MM4_d
+ N_XI0/XI6/XI6/NET34_XI0/XI6/XI6/MM4_g N_VDD_XI0/XI6/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI6/MM10 N_XI0/XI6/XI6/NET35_XI0/XI6/XI6/MM10_d
+ N_XI0/XI6/XI6/NET36_XI0/XI6/XI6/MM10_g N_VDD_XI0/XI6/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI6/MM11 N_XI0/XI6/XI6/NET36_XI0/XI6/XI6/MM11_d
+ N_XI0/XI6/XI6/NET35_XI0/XI6/XI6/MM11_g N_VDD_XI0/XI6/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI7/MM2 N_XI0/XI6/XI7/NET34_XI0/XI6/XI7/MM2_d
+ N_XI0/XI6/XI7/NET33_XI0/XI6/XI7/MM2_g N_VSS_XI0/XI6/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI7/MM3 N_XI0/XI6/XI7/NET33_XI0/XI6/XI7/MM3_d N_WL<8>_XI0/XI6/XI7/MM3_g
+ N_BLN<8>_XI0/XI6/XI7/MM3_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI7/MM0 N_XI0/XI6/XI7/NET34_XI0/XI6/XI7/MM0_d N_WL<8>_XI0/XI6/XI7/MM0_g
+ N_BL<8>_XI0/XI6/XI7/MM0_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI7/MM1 N_XI0/XI6/XI7/NET33_XI0/XI6/XI7/MM1_d
+ N_XI0/XI6/XI7/NET34_XI0/XI6/XI7/MM1_g N_VSS_XI0/XI6/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI7/MM9 N_XI0/XI6/XI7/NET36_XI0/XI6/XI7/MM9_d N_WL<9>_XI0/XI6/XI7/MM9_g
+ N_BL<8>_XI0/XI6/XI7/MM9_s N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI7/MM6 N_XI0/XI6/XI7/NET35_XI0/XI6/XI7/MM6_d
+ N_XI0/XI6/XI7/NET36_XI0/XI6/XI7/MM6_g N_VSS_XI0/XI6/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI7/MM7 N_XI0/XI6/XI7/NET36_XI0/XI6/XI7/MM7_d
+ N_XI0/XI6/XI7/NET35_XI0/XI6/XI7/MM7_g N_VSS_XI0/XI6/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI7/MM8 N_XI0/XI6/XI7/NET35_XI0/XI6/XI7/MM8_d N_WL<9>_XI0/XI6/XI7/MM8_g
+ N_BLN<8>_XI0/XI6/XI7/MM8_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI7/MM5 N_XI0/XI6/XI7/NET34_XI0/XI6/XI7/MM5_d
+ N_XI0/XI6/XI7/NET33_XI0/XI6/XI7/MM5_g N_VDD_XI0/XI6/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI7/MM4 N_XI0/XI6/XI7/NET33_XI0/XI6/XI7/MM4_d
+ N_XI0/XI6/XI7/NET34_XI0/XI6/XI7/MM4_g N_VDD_XI0/XI6/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI7/MM10 N_XI0/XI6/XI7/NET35_XI0/XI6/XI7/MM10_d
+ N_XI0/XI6/XI7/NET36_XI0/XI6/XI7/MM10_g N_VDD_XI0/XI6/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI7/MM11 N_XI0/XI6/XI7/NET36_XI0/XI6/XI7/MM11_d
+ N_XI0/XI6/XI7/NET35_XI0/XI6/XI7/MM11_g N_VDD_XI0/XI6/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI8/MM2 N_XI0/XI6/XI8/NET34_XI0/XI6/XI8/MM2_d
+ N_XI0/XI6/XI8/NET33_XI0/XI6/XI8/MM2_g N_VSS_XI0/XI6/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI8/MM3 N_XI0/XI6/XI8/NET33_XI0/XI6/XI8/MM3_d N_WL<8>_XI0/XI6/XI8/MM3_g
+ N_BLN<7>_XI0/XI6/XI8/MM3_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI8/MM0 N_XI0/XI6/XI8/NET34_XI0/XI6/XI8/MM0_d N_WL<8>_XI0/XI6/XI8/MM0_g
+ N_BL<7>_XI0/XI6/XI8/MM0_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI8/MM1 N_XI0/XI6/XI8/NET33_XI0/XI6/XI8/MM1_d
+ N_XI0/XI6/XI8/NET34_XI0/XI6/XI8/MM1_g N_VSS_XI0/XI6/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI8/MM9 N_XI0/XI6/XI8/NET36_XI0/XI6/XI8/MM9_d N_WL<9>_XI0/XI6/XI8/MM9_g
+ N_BL<7>_XI0/XI6/XI8/MM9_s N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI8/MM6 N_XI0/XI6/XI8/NET35_XI0/XI6/XI8/MM6_d
+ N_XI0/XI6/XI8/NET36_XI0/XI6/XI8/MM6_g N_VSS_XI0/XI6/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI8/MM7 N_XI0/XI6/XI8/NET36_XI0/XI6/XI8/MM7_d
+ N_XI0/XI6/XI8/NET35_XI0/XI6/XI8/MM7_g N_VSS_XI0/XI6/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI8/MM8 N_XI0/XI6/XI8/NET35_XI0/XI6/XI8/MM8_d N_WL<9>_XI0/XI6/XI8/MM8_g
+ N_BLN<7>_XI0/XI6/XI8/MM8_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI8/MM5 N_XI0/XI6/XI8/NET34_XI0/XI6/XI8/MM5_d
+ N_XI0/XI6/XI8/NET33_XI0/XI6/XI8/MM5_g N_VDD_XI0/XI6/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI8/MM4 N_XI0/XI6/XI8/NET33_XI0/XI6/XI8/MM4_d
+ N_XI0/XI6/XI8/NET34_XI0/XI6/XI8/MM4_g N_VDD_XI0/XI6/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI8/MM10 N_XI0/XI6/XI8/NET35_XI0/XI6/XI8/MM10_d
+ N_XI0/XI6/XI8/NET36_XI0/XI6/XI8/MM10_g N_VDD_XI0/XI6/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI8/MM11 N_XI0/XI6/XI8/NET36_XI0/XI6/XI8/MM11_d
+ N_XI0/XI6/XI8/NET35_XI0/XI6/XI8/MM11_g N_VDD_XI0/XI6/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI9/MM2 N_XI0/XI6/XI9/NET34_XI0/XI6/XI9/MM2_d
+ N_XI0/XI6/XI9/NET33_XI0/XI6/XI9/MM2_g N_VSS_XI0/XI6/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI9/MM3 N_XI0/XI6/XI9/NET33_XI0/XI6/XI9/MM3_d N_WL<8>_XI0/XI6/XI9/MM3_g
+ N_BLN<6>_XI0/XI6/XI9/MM3_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI9/MM0 N_XI0/XI6/XI9/NET34_XI0/XI6/XI9/MM0_d N_WL<8>_XI0/XI6/XI9/MM0_g
+ N_BL<6>_XI0/XI6/XI9/MM0_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI9/MM1 N_XI0/XI6/XI9/NET33_XI0/XI6/XI9/MM1_d
+ N_XI0/XI6/XI9/NET34_XI0/XI6/XI9/MM1_g N_VSS_XI0/XI6/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI9/MM9 N_XI0/XI6/XI9/NET36_XI0/XI6/XI9/MM9_d N_WL<9>_XI0/XI6/XI9/MM9_g
+ N_BL<6>_XI0/XI6/XI9/MM9_s N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI9/MM6 N_XI0/XI6/XI9/NET35_XI0/XI6/XI9/MM6_d
+ N_XI0/XI6/XI9/NET36_XI0/XI6/XI9/MM6_g N_VSS_XI0/XI6/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI9/MM7 N_XI0/XI6/XI9/NET36_XI0/XI6/XI9/MM7_d
+ N_XI0/XI6/XI9/NET35_XI0/XI6/XI9/MM7_g N_VSS_XI0/XI6/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI9/MM8 N_XI0/XI6/XI9/NET35_XI0/XI6/XI9/MM8_d N_WL<9>_XI0/XI6/XI9/MM8_g
+ N_BLN<6>_XI0/XI6/XI9/MM8_s N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI6/XI9/MM5 N_XI0/XI6/XI9/NET34_XI0/XI6/XI9/MM5_d
+ N_XI0/XI6/XI9/NET33_XI0/XI6/XI9/MM5_g N_VDD_XI0/XI6/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI9/MM4 N_XI0/XI6/XI9/NET33_XI0/XI6/XI9/MM4_d
+ N_XI0/XI6/XI9/NET34_XI0/XI6/XI9/MM4_g N_VDD_XI0/XI6/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI9/MM10 N_XI0/XI6/XI9/NET35_XI0/XI6/XI9/MM10_d
+ N_XI0/XI6/XI9/NET36_XI0/XI6/XI9/MM10_g N_VDD_XI0/XI6/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI9/MM11 N_XI0/XI6/XI9/NET36_XI0/XI6/XI9/MM11_d
+ N_XI0/XI6/XI9/NET35_XI0/XI6/XI9/MM11_g N_VDD_XI0/XI6/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI10/MM2 N_XI0/XI6/XI10/NET34_XI0/XI6/XI10/MM2_d
+ N_XI0/XI6/XI10/NET33_XI0/XI6/XI10/MM2_g N_VSS_XI0/XI6/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM3 N_XI0/XI6/XI10/NET33_XI0/XI6/XI10/MM3_d
+ N_WL<8>_XI0/XI6/XI10/MM3_g N_BLN<5>_XI0/XI6/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM0 N_XI0/XI6/XI10/NET34_XI0/XI6/XI10/MM0_d
+ N_WL<8>_XI0/XI6/XI10/MM0_g N_BL<5>_XI0/XI6/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM1 N_XI0/XI6/XI10/NET33_XI0/XI6/XI10/MM1_d
+ N_XI0/XI6/XI10/NET34_XI0/XI6/XI10/MM1_g N_VSS_XI0/XI6/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM9 N_XI0/XI6/XI10/NET36_XI0/XI6/XI10/MM9_d
+ N_WL<9>_XI0/XI6/XI10/MM9_g N_BL<5>_XI0/XI6/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM6 N_XI0/XI6/XI10/NET35_XI0/XI6/XI10/MM6_d
+ N_XI0/XI6/XI10/NET36_XI0/XI6/XI10/MM6_g N_VSS_XI0/XI6/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM7 N_XI0/XI6/XI10/NET36_XI0/XI6/XI10/MM7_d
+ N_XI0/XI6/XI10/NET35_XI0/XI6/XI10/MM7_g N_VSS_XI0/XI6/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM8 N_XI0/XI6/XI10/NET35_XI0/XI6/XI10/MM8_d
+ N_WL<9>_XI0/XI6/XI10/MM8_g N_BLN<5>_XI0/XI6/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI10/MM5 N_XI0/XI6/XI10/NET34_XI0/XI6/XI10/MM5_d
+ N_XI0/XI6/XI10/NET33_XI0/XI6/XI10/MM5_g N_VDD_XI0/XI6/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI10/MM4 N_XI0/XI6/XI10/NET33_XI0/XI6/XI10/MM4_d
+ N_XI0/XI6/XI10/NET34_XI0/XI6/XI10/MM4_g N_VDD_XI0/XI6/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI10/MM10 N_XI0/XI6/XI10/NET35_XI0/XI6/XI10/MM10_d
+ N_XI0/XI6/XI10/NET36_XI0/XI6/XI10/MM10_g N_VDD_XI0/XI6/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI10/MM11 N_XI0/XI6/XI10/NET36_XI0/XI6/XI10/MM11_d
+ N_XI0/XI6/XI10/NET35_XI0/XI6/XI10/MM11_g N_VDD_XI0/XI6/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI11/MM2 N_XI0/XI6/XI11/NET34_XI0/XI6/XI11/MM2_d
+ N_XI0/XI6/XI11/NET33_XI0/XI6/XI11/MM2_g N_VSS_XI0/XI6/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM3 N_XI0/XI6/XI11/NET33_XI0/XI6/XI11/MM3_d
+ N_WL<8>_XI0/XI6/XI11/MM3_g N_BLN<4>_XI0/XI6/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM0 N_XI0/XI6/XI11/NET34_XI0/XI6/XI11/MM0_d
+ N_WL<8>_XI0/XI6/XI11/MM0_g N_BL<4>_XI0/XI6/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM1 N_XI0/XI6/XI11/NET33_XI0/XI6/XI11/MM1_d
+ N_XI0/XI6/XI11/NET34_XI0/XI6/XI11/MM1_g N_VSS_XI0/XI6/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM9 N_XI0/XI6/XI11/NET36_XI0/XI6/XI11/MM9_d
+ N_WL<9>_XI0/XI6/XI11/MM9_g N_BL<4>_XI0/XI6/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM6 N_XI0/XI6/XI11/NET35_XI0/XI6/XI11/MM6_d
+ N_XI0/XI6/XI11/NET36_XI0/XI6/XI11/MM6_g N_VSS_XI0/XI6/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM7 N_XI0/XI6/XI11/NET36_XI0/XI6/XI11/MM7_d
+ N_XI0/XI6/XI11/NET35_XI0/XI6/XI11/MM7_g N_VSS_XI0/XI6/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM8 N_XI0/XI6/XI11/NET35_XI0/XI6/XI11/MM8_d
+ N_WL<9>_XI0/XI6/XI11/MM8_g N_BLN<4>_XI0/XI6/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI11/MM5 N_XI0/XI6/XI11/NET34_XI0/XI6/XI11/MM5_d
+ N_XI0/XI6/XI11/NET33_XI0/XI6/XI11/MM5_g N_VDD_XI0/XI6/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI11/MM4 N_XI0/XI6/XI11/NET33_XI0/XI6/XI11/MM4_d
+ N_XI0/XI6/XI11/NET34_XI0/XI6/XI11/MM4_g N_VDD_XI0/XI6/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI11/MM10 N_XI0/XI6/XI11/NET35_XI0/XI6/XI11/MM10_d
+ N_XI0/XI6/XI11/NET36_XI0/XI6/XI11/MM10_g N_VDD_XI0/XI6/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI11/MM11 N_XI0/XI6/XI11/NET36_XI0/XI6/XI11/MM11_d
+ N_XI0/XI6/XI11/NET35_XI0/XI6/XI11/MM11_g N_VDD_XI0/XI6/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI12/MM2 N_XI0/XI6/XI12/NET34_XI0/XI6/XI12/MM2_d
+ N_XI0/XI6/XI12/NET33_XI0/XI6/XI12/MM2_g N_VSS_XI0/XI6/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM3 N_XI0/XI6/XI12/NET33_XI0/XI6/XI12/MM3_d
+ N_WL<8>_XI0/XI6/XI12/MM3_g N_BLN<3>_XI0/XI6/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM0 N_XI0/XI6/XI12/NET34_XI0/XI6/XI12/MM0_d
+ N_WL<8>_XI0/XI6/XI12/MM0_g N_BL<3>_XI0/XI6/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM1 N_XI0/XI6/XI12/NET33_XI0/XI6/XI12/MM1_d
+ N_XI0/XI6/XI12/NET34_XI0/XI6/XI12/MM1_g N_VSS_XI0/XI6/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM9 N_XI0/XI6/XI12/NET36_XI0/XI6/XI12/MM9_d
+ N_WL<9>_XI0/XI6/XI12/MM9_g N_BL<3>_XI0/XI6/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM6 N_XI0/XI6/XI12/NET35_XI0/XI6/XI12/MM6_d
+ N_XI0/XI6/XI12/NET36_XI0/XI6/XI12/MM6_g N_VSS_XI0/XI6/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM7 N_XI0/XI6/XI12/NET36_XI0/XI6/XI12/MM7_d
+ N_XI0/XI6/XI12/NET35_XI0/XI6/XI12/MM7_g N_VSS_XI0/XI6/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM8 N_XI0/XI6/XI12/NET35_XI0/XI6/XI12/MM8_d
+ N_WL<9>_XI0/XI6/XI12/MM8_g N_BLN<3>_XI0/XI6/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI12/MM5 N_XI0/XI6/XI12/NET34_XI0/XI6/XI12/MM5_d
+ N_XI0/XI6/XI12/NET33_XI0/XI6/XI12/MM5_g N_VDD_XI0/XI6/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI12/MM4 N_XI0/XI6/XI12/NET33_XI0/XI6/XI12/MM4_d
+ N_XI0/XI6/XI12/NET34_XI0/XI6/XI12/MM4_g N_VDD_XI0/XI6/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI12/MM10 N_XI0/XI6/XI12/NET35_XI0/XI6/XI12/MM10_d
+ N_XI0/XI6/XI12/NET36_XI0/XI6/XI12/MM10_g N_VDD_XI0/XI6/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI12/MM11 N_XI0/XI6/XI12/NET36_XI0/XI6/XI12/MM11_d
+ N_XI0/XI6/XI12/NET35_XI0/XI6/XI12/MM11_g N_VDD_XI0/XI6/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI13/MM2 N_XI0/XI6/XI13/NET34_XI0/XI6/XI13/MM2_d
+ N_XI0/XI6/XI13/NET33_XI0/XI6/XI13/MM2_g N_VSS_XI0/XI6/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM3 N_XI0/XI6/XI13/NET33_XI0/XI6/XI13/MM3_d
+ N_WL<8>_XI0/XI6/XI13/MM3_g N_BLN<2>_XI0/XI6/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM0 N_XI0/XI6/XI13/NET34_XI0/XI6/XI13/MM0_d
+ N_WL<8>_XI0/XI6/XI13/MM0_g N_BL<2>_XI0/XI6/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM1 N_XI0/XI6/XI13/NET33_XI0/XI6/XI13/MM1_d
+ N_XI0/XI6/XI13/NET34_XI0/XI6/XI13/MM1_g N_VSS_XI0/XI6/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM9 N_XI0/XI6/XI13/NET36_XI0/XI6/XI13/MM9_d
+ N_WL<9>_XI0/XI6/XI13/MM9_g N_BL<2>_XI0/XI6/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM6 N_XI0/XI6/XI13/NET35_XI0/XI6/XI13/MM6_d
+ N_XI0/XI6/XI13/NET36_XI0/XI6/XI13/MM6_g N_VSS_XI0/XI6/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM7 N_XI0/XI6/XI13/NET36_XI0/XI6/XI13/MM7_d
+ N_XI0/XI6/XI13/NET35_XI0/XI6/XI13/MM7_g N_VSS_XI0/XI6/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM8 N_XI0/XI6/XI13/NET35_XI0/XI6/XI13/MM8_d
+ N_WL<9>_XI0/XI6/XI13/MM8_g N_BLN<2>_XI0/XI6/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI13/MM5 N_XI0/XI6/XI13/NET34_XI0/XI6/XI13/MM5_d
+ N_XI0/XI6/XI13/NET33_XI0/XI6/XI13/MM5_g N_VDD_XI0/XI6/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI13/MM4 N_XI0/XI6/XI13/NET33_XI0/XI6/XI13/MM4_d
+ N_XI0/XI6/XI13/NET34_XI0/XI6/XI13/MM4_g N_VDD_XI0/XI6/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI13/MM10 N_XI0/XI6/XI13/NET35_XI0/XI6/XI13/MM10_d
+ N_XI0/XI6/XI13/NET36_XI0/XI6/XI13/MM10_g N_VDD_XI0/XI6/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI13/MM11 N_XI0/XI6/XI13/NET36_XI0/XI6/XI13/MM11_d
+ N_XI0/XI6/XI13/NET35_XI0/XI6/XI13/MM11_g N_VDD_XI0/XI6/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI14/MM2 N_XI0/XI6/XI14/NET34_XI0/XI6/XI14/MM2_d
+ N_XI0/XI6/XI14/NET33_XI0/XI6/XI14/MM2_g N_VSS_XI0/XI6/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM3 N_XI0/XI6/XI14/NET33_XI0/XI6/XI14/MM3_d
+ N_WL<8>_XI0/XI6/XI14/MM3_g N_BLN<1>_XI0/XI6/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM0 N_XI0/XI6/XI14/NET34_XI0/XI6/XI14/MM0_d
+ N_WL<8>_XI0/XI6/XI14/MM0_g N_BL<1>_XI0/XI6/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM1 N_XI0/XI6/XI14/NET33_XI0/XI6/XI14/MM1_d
+ N_XI0/XI6/XI14/NET34_XI0/XI6/XI14/MM1_g N_VSS_XI0/XI6/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM9 N_XI0/XI6/XI14/NET36_XI0/XI6/XI14/MM9_d
+ N_WL<9>_XI0/XI6/XI14/MM9_g N_BL<1>_XI0/XI6/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM6 N_XI0/XI6/XI14/NET35_XI0/XI6/XI14/MM6_d
+ N_XI0/XI6/XI14/NET36_XI0/XI6/XI14/MM6_g N_VSS_XI0/XI6/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM7 N_XI0/XI6/XI14/NET36_XI0/XI6/XI14/MM7_d
+ N_XI0/XI6/XI14/NET35_XI0/XI6/XI14/MM7_g N_VSS_XI0/XI6/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM8 N_XI0/XI6/XI14/NET35_XI0/XI6/XI14/MM8_d
+ N_WL<9>_XI0/XI6/XI14/MM8_g N_BLN<1>_XI0/XI6/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI14/MM5 N_XI0/XI6/XI14/NET34_XI0/XI6/XI14/MM5_d
+ N_XI0/XI6/XI14/NET33_XI0/XI6/XI14/MM5_g N_VDD_XI0/XI6/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI14/MM4 N_XI0/XI6/XI14/NET33_XI0/XI6/XI14/MM4_d
+ N_XI0/XI6/XI14/NET34_XI0/XI6/XI14/MM4_g N_VDD_XI0/XI6/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI14/MM10 N_XI0/XI6/XI14/NET35_XI0/XI6/XI14/MM10_d
+ N_XI0/XI6/XI14/NET36_XI0/XI6/XI14/MM10_g N_VDD_XI0/XI6/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI14/MM11 N_XI0/XI6/XI14/NET36_XI0/XI6/XI14/MM11_d
+ N_XI0/XI6/XI14/NET35_XI0/XI6/XI14/MM11_g N_VDD_XI0/XI6/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI15/MM2 N_XI0/XI6/XI15/NET34_XI0/XI6/XI15/MM2_d
+ N_XI0/XI6/XI15/NET33_XI0/XI6/XI15/MM2_g N_VSS_XI0/XI6/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM3 N_XI0/XI6/XI15/NET33_XI0/XI6/XI15/MM3_d
+ N_WL<8>_XI0/XI6/XI15/MM3_g N_BLN<0>_XI0/XI6/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM0 N_XI0/XI6/XI15/NET34_XI0/XI6/XI15/MM0_d
+ N_WL<8>_XI0/XI6/XI15/MM0_g N_BL<0>_XI0/XI6/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM1 N_XI0/XI6/XI15/NET33_XI0/XI6/XI15/MM1_d
+ N_XI0/XI6/XI15/NET34_XI0/XI6/XI15/MM1_g N_VSS_XI0/XI6/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM9 N_XI0/XI6/XI15/NET36_XI0/XI6/XI15/MM9_d
+ N_WL<9>_XI0/XI6/XI15/MM9_g N_BL<0>_XI0/XI6/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM6 N_XI0/XI6/XI15/NET35_XI0/XI6/XI15/MM6_d
+ N_XI0/XI6/XI15/NET36_XI0/XI6/XI15/MM6_g N_VSS_XI0/XI6/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM7 N_XI0/XI6/XI15/NET36_XI0/XI6/XI15/MM7_d
+ N_XI0/XI6/XI15/NET35_XI0/XI6/XI15/MM7_g N_VSS_XI0/XI6/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM8 N_XI0/XI6/XI15/NET35_XI0/XI6/XI15/MM8_d
+ N_WL<9>_XI0/XI6/XI15/MM8_g N_BLN<0>_XI0/XI6/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/XI15/MM5 N_XI0/XI6/XI15/NET34_XI0/XI6/XI15/MM5_d
+ N_XI0/XI6/XI15/NET33_XI0/XI6/XI15/MM5_g N_VDD_XI0/XI6/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI15/MM4 N_XI0/XI6/XI15/NET33_XI0/XI6/XI15/MM4_d
+ N_XI0/XI6/XI15/NET34_XI0/XI6/XI15/MM4_g N_VDD_XI0/XI6/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI15/MM10 N_XI0/XI6/XI15/NET35_XI0/XI6/XI15/MM10_d
+ N_XI0/XI6/XI15/NET36_XI0/XI6/XI15/MM10_g N_VDD_XI0/XI6/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/XI15/MM11 N_XI0/XI6/XI15/NET36_XI0/XI6/XI15/MM11_d
+ N_XI0/XI6/XI15/NET35_XI0/XI6/XI15/MM11_g N_VDD_XI0/XI6/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI0/MM2 N_XI0/XI7/XI0/NET34_XI0/XI7/XI0/MM2_d
+ N_XI0/XI7/XI0/NET33_XI0/XI7/XI0/MM2_g N_VSS_XI0/XI7/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM3 N_XI0/XI7/XI0/NET33_XI0/XI7/XI0/MM3_d
+ N_WL<10>_XI0/XI7/XI0/MM3_g N_BLN<15>_XI0/XI7/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM0 N_XI0/XI7/XI0/NET34_XI0/XI7/XI0/MM0_d
+ N_WL<10>_XI0/XI7/XI0/MM0_g N_BL<15>_XI0/XI7/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM1 N_XI0/XI7/XI0/NET33_XI0/XI7/XI0/MM1_d
+ N_XI0/XI7/XI0/NET34_XI0/XI7/XI0/MM1_g N_VSS_XI0/XI7/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM9 N_XI0/XI7/XI0/NET36_XI0/XI7/XI0/MM9_d
+ N_WL<11>_XI0/XI7/XI0/MM9_g N_BL<15>_XI0/XI7/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM6 N_XI0/XI7/XI0/NET35_XI0/XI7/XI0/MM6_d
+ N_XI0/XI7/XI0/NET36_XI0/XI7/XI0/MM6_g N_VSS_XI0/XI7/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM7 N_XI0/XI7/XI0/NET36_XI0/XI7/XI0/MM7_d
+ N_XI0/XI7/XI0/NET35_XI0/XI7/XI0/MM7_g N_VSS_XI0/XI7/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM8 N_XI0/XI7/XI0/NET35_XI0/XI7/XI0/MM8_d
+ N_WL<11>_XI0/XI7/XI0/MM8_g N_BLN<15>_XI0/XI7/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI0/MM5 N_XI0/XI7/XI0/NET34_XI0/XI7/XI0/MM5_d
+ N_XI0/XI7/XI0/NET33_XI0/XI7/XI0/MM5_g N_VDD_XI0/XI7/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI0/MM4 N_XI0/XI7/XI0/NET33_XI0/XI7/XI0/MM4_d
+ N_XI0/XI7/XI0/NET34_XI0/XI7/XI0/MM4_g N_VDD_XI0/XI7/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI0/MM10 N_XI0/XI7/XI0/NET35_XI0/XI7/XI0/MM10_d
+ N_XI0/XI7/XI0/NET36_XI0/XI7/XI0/MM10_g N_VDD_XI0/XI7/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI0/MM11 N_XI0/XI7/XI0/NET36_XI0/XI7/XI0/MM11_d
+ N_XI0/XI7/XI0/NET35_XI0/XI7/XI0/MM11_g N_VDD_XI0/XI7/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI1/MM2 N_XI0/XI7/XI1/NET34_XI0/XI7/XI1/MM2_d
+ N_XI0/XI7/XI1/NET33_XI0/XI7/XI1/MM2_g N_VSS_XI0/XI7/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM3 N_XI0/XI7/XI1/NET33_XI0/XI7/XI1/MM3_d
+ N_WL<10>_XI0/XI7/XI1/MM3_g N_BLN<14>_XI0/XI7/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM0 N_XI0/XI7/XI1/NET34_XI0/XI7/XI1/MM0_d
+ N_WL<10>_XI0/XI7/XI1/MM0_g N_BL<14>_XI0/XI7/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM1 N_XI0/XI7/XI1/NET33_XI0/XI7/XI1/MM1_d
+ N_XI0/XI7/XI1/NET34_XI0/XI7/XI1/MM1_g N_VSS_XI0/XI7/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM9 N_XI0/XI7/XI1/NET36_XI0/XI7/XI1/MM9_d
+ N_WL<11>_XI0/XI7/XI1/MM9_g N_BL<14>_XI0/XI7/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM6 N_XI0/XI7/XI1/NET35_XI0/XI7/XI1/MM6_d
+ N_XI0/XI7/XI1/NET36_XI0/XI7/XI1/MM6_g N_VSS_XI0/XI7/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM7 N_XI0/XI7/XI1/NET36_XI0/XI7/XI1/MM7_d
+ N_XI0/XI7/XI1/NET35_XI0/XI7/XI1/MM7_g N_VSS_XI0/XI7/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM8 N_XI0/XI7/XI1/NET35_XI0/XI7/XI1/MM8_d
+ N_WL<11>_XI0/XI7/XI1/MM8_g N_BLN<14>_XI0/XI7/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI1/MM5 N_XI0/XI7/XI1/NET34_XI0/XI7/XI1/MM5_d
+ N_XI0/XI7/XI1/NET33_XI0/XI7/XI1/MM5_g N_VDD_XI0/XI7/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI1/MM4 N_XI0/XI7/XI1/NET33_XI0/XI7/XI1/MM4_d
+ N_XI0/XI7/XI1/NET34_XI0/XI7/XI1/MM4_g N_VDD_XI0/XI7/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI1/MM10 N_XI0/XI7/XI1/NET35_XI0/XI7/XI1/MM10_d
+ N_XI0/XI7/XI1/NET36_XI0/XI7/XI1/MM10_g N_VDD_XI0/XI7/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI1/MM11 N_XI0/XI7/XI1/NET36_XI0/XI7/XI1/MM11_d
+ N_XI0/XI7/XI1/NET35_XI0/XI7/XI1/MM11_g N_VDD_XI0/XI7/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI2/MM2 N_XI0/XI7/XI2/NET34_XI0/XI7/XI2/MM2_d
+ N_XI0/XI7/XI2/NET33_XI0/XI7/XI2/MM2_g N_VSS_XI0/XI7/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM3 N_XI0/XI7/XI2/NET33_XI0/XI7/XI2/MM3_d
+ N_WL<10>_XI0/XI7/XI2/MM3_g N_BLN<13>_XI0/XI7/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM0 N_XI0/XI7/XI2/NET34_XI0/XI7/XI2/MM0_d
+ N_WL<10>_XI0/XI7/XI2/MM0_g N_BL<13>_XI0/XI7/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM1 N_XI0/XI7/XI2/NET33_XI0/XI7/XI2/MM1_d
+ N_XI0/XI7/XI2/NET34_XI0/XI7/XI2/MM1_g N_VSS_XI0/XI7/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM9 N_XI0/XI7/XI2/NET36_XI0/XI7/XI2/MM9_d
+ N_WL<11>_XI0/XI7/XI2/MM9_g N_BL<13>_XI0/XI7/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM6 N_XI0/XI7/XI2/NET35_XI0/XI7/XI2/MM6_d
+ N_XI0/XI7/XI2/NET36_XI0/XI7/XI2/MM6_g N_VSS_XI0/XI7/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM7 N_XI0/XI7/XI2/NET36_XI0/XI7/XI2/MM7_d
+ N_XI0/XI7/XI2/NET35_XI0/XI7/XI2/MM7_g N_VSS_XI0/XI7/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM8 N_XI0/XI7/XI2/NET35_XI0/XI7/XI2/MM8_d
+ N_WL<11>_XI0/XI7/XI2/MM8_g N_BLN<13>_XI0/XI7/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI2/MM5 N_XI0/XI7/XI2/NET34_XI0/XI7/XI2/MM5_d
+ N_XI0/XI7/XI2/NET33_XI0/XI7/XI2/MM5_g N_VDD_XI0/XI7/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI2/MM4 N_XI0/XI7/XI2/NET33_XI0/XI7/XI2/MM4_d
+ N_XI0/XI7/XI2/NET34_XI0/XI7/XI2/MM4_g N_VDD_XI0/XI7/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI2/MM10 N_XI0/XI7/XI2/NET35_XI0/XI7/XI2/MM10_d
+ N_XI0/XI7/XI2/NET36_XI0/XI7/XI2/MM10_g N_VDD_XI0/XI7/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI2/MM11 N_XI0/XI7/XI2/NET36_XI0/XI7/XI2/MM11_d
+ N_XI0/XI7/XI2/NET35_XI0/XI7/XI2/MM11_g N_VDD_XI0/XI7/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI3/MM2 N_XI0/XI7/XI3/NET34_XI0/XI7/XI3/MM2_d
+ N_XI0/XI7/XI3/NET33_XI0/XI7/XI3/MM2_g N_VSS_XI0/XI7/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM3 N_XI0/XI7/XI3/NET33_XI0/XI7/XI3/MM3_d
+ N_WL<10>_XI0/XI7/XI3/MM3_g N_BLN<12>_XI0/XI7/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM0 N_XI0/XI7/XI3/NET34_XI0/XI7/XI3/MM0_d
+ N_WL<10>_XI0/XI7/XI3/MM0_g N_BL<12>_XI0/XI7/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM1 N_XI0/XI7/XI3/NET33_XI0/XI7/XI3/MM1_d
+ N_XI0/XI7/XI3/NET34_XI0/XI7/XI3/MM1_g N_VSS_XI0/XI7/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM9 N_XI0/XI7/XI3/NET36_XI0/XI7/XI3/MM9_d
+ N_WL<11>_XI0/XI7/XI3/MM9_g N_BL<12>_XI0/XI7/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM6 N_XI0/XI7/XI3/NET35_XI0/XI7/XI3/MM6_d
+ N_XI0/XI7/XI3/NET36_XI0/XI7/XI3/MM6_g N_VSS_XI0/XI7/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM7 N_XI0/XI7/XI3/NET36_XI0/XI7/XI3/MM7_d
+ N_XI0/XI7/XI3/NET35_XI0/XI7/XI3/MM7_g N_VSS_XI0/XI7/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM8 N_XI0/XI7/XI3/NET35_XI0/XI7/XI3/MM8_d
+ N_WL<11>_XI0/XI7/XI3/MM8_g N_BLN<12>_XI0/XI7/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI3/MM5 N_XI0/XI7/XI3/NET34_XI0/XI7/XI3/MM5_d
+ N_XI0/XI7/XI3/NET33_XI0/XI7/XI3/MM5_g N_VDD_XI0/XI7/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI3/MM4 N_XI0/XI7/XI3/NET33_XI0/XI7/XI3/MM4_d
+ N_XI0/XI7/XI3/NET34_XI0/XI7/XI3/MM4_g N_VDD_XI0/XI7/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI3/MM10 N_XI0/XI7/XI3/NET35_XI0/XI7/XI3/MM10_d
+ N_XI0/XI7/XI3/NET36_XI0/XI7/XI3/MM10_g N_VDD_XI0/XI7/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI3/MM11 N_XI0/XI7/XI3/NET36_XI0/XI7/XI3/MM11_d
+ N_XI0/XI7/XI3/NET35_XI0/XI7/XI3/MM11_g N_VDD_XI0/XI7/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI4/MM2 N_XI0/XI7/XI4/NET34_XI0/XI7/XI4/MM2_d
+ N_XI0/XI7/XI4/NET33_XI0/XI7/XI4/MM2_g N_VSS_XI0/XI7/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM3 N_XI0/XI7/XI4/NET33_XI0/XI7/XI4/MM3_d
+ N_WL<10>_XI0/XI7/XI4/MM3_g N_BLN<11>_XI0/XI7/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM0 N_XI0/XI7/XI4/NET34_XI0/XI7/XI4/MM0_d
+ N_WL<10>_XI0/XI7/XI4/MM0_g N_BL<11>_XI0/XI7/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM1 N_XI0/XI7/XI4/NET33_XI0/XI7/XI4/MM1_d
+ N_XI0/XI7/XI4/NET34_XI0/XI7/XI4/MM1_g N_VSS_XI0/XI7/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM9 N_XI0/XI7/XI4/NET36_XI0/XI7/XI4/MM9_d
+ N_WL<11>_XI0/XI7/XI4/MM9_g N_BL<11>_XI0/XI7/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM6 N_XI0/XI7/XI4/NET35_XI0/XI7/XI4/MM6_d
+ N_XI0/XI7/XI4/NET36_XI0/XI7/XI4/MM6_g N_VSS_XI0/XI7/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM7 N_XI0/XI7/XI4/NET36_XI0/XI7/XI4/MM7_d
+ N_XI0/XI7/XI4/NET35_XI0/XI7/XI4/MM7_g N_VSS_XI0/XI7/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM8 N_XI0/XI7/XI4/NET35_XI0/XI7/XI4/MM8_d
+ N_WL<11>_XI0/XI7/XI4/MM8_g N_BLN<11>_XI0/XI7/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI4/MM5 N_XI0/XI7/XI4/NET34_XI0/XI7/XI4/MM5_d
+ N_XI0/XI7/XI4/NET33_XI0/XI7/XI4/MM5_g N_VDD_XI0/XI7/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI4/MM4 N_XI0/XI7/XI4/NET33_XI0/XI7/XI4/MM4_d
+ N_XI0/XI7/XI4/NET34_XI0/XI7/XI4/MM4_g N_VDD_XI0/XI7/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI4/MM10 N_XI0/XI7/XI4/NET35_XI0/XI7/XI4/MM10_d
+ N_XI0/XI7/XI4/NET36_XI0/XI7/XI4/MM10_g N_VDD_XI0/XI7/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI4/MM11 N_XI0/XI7/XI4/NET36_XI0/XI7/XI4/MM11_d
+ N_XI0/XI7/XI4/NET35_XI0/XI7/XI4/MM11_g N_VDD_XI0/XI7/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI5/MM2 N_XI0/XI7/XI5/NET34_XI0/XI7/XI5/MM2_d
+ N_XI0/XI7/XI5/NET33_XI0/XI7/XI5/MM2_g N_VSS_XI0/XI7/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM3 N_XI0/XI7/XI5/NET33_XI0/XI7/XI5/MM3_d
+ N_WL<10>_XI0/XI7/XI5/MM3_g N_BLN<10>_XI0/XI7/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM0 N_XI0/XI7/XI5/NET34_XI0/XI7/XI5/MM0_d
+ N_WL<10>_XI0/XI7/XI5/MM0_g N_BL<10>_XI0/XI7/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM1 N_XI0/XI7/XI5/NET33_XI0/XI7/XI5/MM1_d
+ N_XI0/XI7/XI5/NET34_XI0/XI7/XI5/MM1_g N_VSS_XI0/XI7/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM9 N_XI0/XI7/XI5/NET36_XI0/XI7/XI5/MM9_d
+ N_WL<11>_XI0/XI7/XI5/MM9_g N_BL<10>_XI0/XI7/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM6 N_XI0/XI7/XI5/NET35_XI0/XI7/XI5/MM6_d
+ N_XI0/XI7/XI5/NET36_XI0/XI7/XI5/MM6_g N_VSS_XI0/XI7/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM7 N_XI0/XI7/XI5/NET36_XI0/XI7/XI5/MM7_d
+ N_XI0/XI7/XI5/NET35_XI0/XI7/XI5/MM7_g N_VSS_XI0/XI7/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM8 N_XI0/XI7/XI5/NET35_XI0/XI7/XI5/MM8_d
+ N_WL<11>_XI0/XI7/XI5/MM8_g N_BLN<10>_XI0/XI7/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI5/MM5 N_XI0/XI7/XI5/NET34_XI0/XI7/XI5/MM5_d
+ N_XI0/XI7/XI5/NET33_XI0/XI7/XI5/MM5_g N_VDD_XI0/XI7/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI5/MM4 N_XI0/XI7/XI5/NET33_XI0/XI7/XI5/MM4_d
+ N_XI0/XI7/XI5/NET34_XI0/XI7/XI5/MM4_g N_VDD_XI0/XI7/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI5/MM10 N_XI0/XI7/XI5/NET35_XI0/XI7/XI5/MM10_d
+ N_XI0/XI7/XI5/NET36_XI0/XI7/XI5/MM10_g N_VDD_XI0/XI7/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI5/MM11 N_XI0/XI7/XI5/NET36_XI0/XI7/XI5/MM11_d
+ N_XI0/XI7/XI5/NET35_XI0/XI7/XI5/MM11_g N_VDD_XI0/XI7/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI6/MM2 N_XI0/XI7/XI6/NET34_XI0/XI7/XI6/MM2_d
+ N_XI0/XI7/XI6/NET33_XI0/XI7/XI6/MM2_g N_VSS_XI0/XI7/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM3 N_XI0/XI7/XI6/NET33_XI0/XI7/XI6/MM3_d
+ N_WL<10>_XI0/XI7/XI6/MM3_g N_BLN<9>_XI0/XI7/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM0 N_XI0/XI7/XI6/NET34_XI0/XI7/XI6/MM0_d
+ N_WL<10>_XI0/XI7/XI6/MM0_g N_BL<9>_XI0/XI7/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM1 N_XI0/XI7/XI6/NET33_XI0/XI7/XI6/MM1_d
+ N_XI0/XI7/XI6/NET34_XI0/XI7/XI6/MM1_g N_VSS_XI0/XI7/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM9 N_XI0/XI7/XI6/NET36_XI0/XI7/XI6/MM9_d
+ N_WL<11>_XI0/XI7/XI6/MM9_g N_BL<9>_XI0/XI7/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM6 N_XI0/XI7/XI6/NET35_XI0/XI7/XI6/MM6_d
+ N_XI0/XI7/XI6/NET36_XI0/XI7/XI6/MM6_g N_VSS_XI0/XI7/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM7 N_XI0/XI7/XI6/NET36_XI0/XI7/XI6/MM7_d
+ N_XI0/XI7/XI6/NET35_XI0/XI7/XI6/MM7_g N_VSS_XI0/XI7/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM8 N_XI0/XI7/XI6/NET35_XI0/XI7/XI6/MM8_d
+ N_WL<11>_XI0/XI7/XI6/MM8_g N_BLN<9>_XI0/XI7/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI6/MM5 N_XI0/XI7/XI6/NET34_XI0/XI7/XI6/MM5_d
+ N_XI0/XI7/XI6/NET33_XI0/XI7/XI6/MM5_g N_VDD_XI0/XI7/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI6/MM4 N_XI0/XI7/XI6/NET33_XI0/XI7/XI6/MM4_d
+ N_XI0/XI7/XI6/NET34_XI0/XI7/XI6/MM4_g N_VDD_XI0/XI7/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI6/MM10 N_XI0/XI7/XI6/NET35_XI0/XI7/XI6/MM10_d
+ N_XI0/XI7/XI6/NET36_XI0/XI7/XI6/MM10_g N_VDD_XI0/XI7/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI6/MM11 N_XI0/XI7/XI6/NET36_XI0/XI7/XI6/MM11_d
+ N_XI0/XI7/XI6/NET35_XI0/XI7/XI6/MM11_g N_VDD_XI0/XI7/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI7/MM2 N_XI0/XI7/XI7/NET34_XI0/XI7/XI7/MM2_d
+ N_XI0/XI7/XI7/NET33_XI0/XI7/XI7/MM2_g N_VSS_XI0/XI7/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM3 N_XI0/XI7/XI7/NET33_XI0/XI7/XI7/MM3_d
+ N_WL<10>_XI0/XI7/XI7/MM3_g N_BLN<8>_XI0/XI7/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM0 N_XI0/XI7/XI7/NET34_XI0/XI7/XI7/MM0_d
+ N_WL<10>_XI0/XI7/XI7/MM0_g N_BL<8>_XI0/XI7/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM1 N_XI0/XI7/XI7/NET33_XI0/XI7/XI7/MM1_d
+ N_XI0/XI7/XI7/NET34_XI0/XI7/XI7/MM1_g N_VSS_XI0/XI7/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM9 N_XI0/XI7/XI7/NET36_XI0/XI7/XI7/MM9_d
+ N_WL<11>_XI0/XI7/XI7/MM9_g N_BL<8>_XI0/XI7/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM6 N_XI0/XI7/XI7/NET35_XI0/XI7/XI7/MM6_d
+ N_XI0/XI7/XI7/NET36_XI0/XI7/XI7/MM6_g N_VSS_XI0/XI7/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM7 N_XI0/XI7/XI7/NET36_XI0/XI7/XI7/MM7_d
+ N_XI0/XI7/XI7/NET35_XI0/XI7/XI7/MM7_g N_VSS_XI0/XI7/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM8 N_XI0/XI7/XI7/NET35_XI0/XI7/XI7/MM8_d
+ N_WL<11>_XI0/XI7/XI7/MM8_g N_BLN<8>_XI0/XI7/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI7/MM5 N_XI0/XI7/XI7/NET34_XI0/XI7/XI7/MM5_d
+ N_XI0/XI7/XI7/NET33_XI0/XI7/XI7/MM5_g N_VDD_XI0/XI7/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI7/MM4 N_XI0/XI7/XI7/NET33_XI0/XI7/XI7/MM4_d
+ N_XI0/XI7/XI7/NET34_XI0/XI7/XI7/MM4_g N_VDD_XI0/XI7/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI7/MM10 N_XI0/XI7/XI7/NET35_XI0/XI7/XI7/MM10_d
+ N_XI0/XI7/XI7/NET36_XI0/XI7/XI7/MM10_g N_VDD_XI0/XI7/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI7/MM11 N_XI0/XI7/XI7/NET36_XI0/XI7/XI7/MM11_d
+ N_XI0/XI7/XI7/NET35_XI0/XI7/XI7/MM11_g N_VDD_XI0/XI7/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI8/MM2 N_XI0/XI7/XI8/NET34_XI0/XI7/XI8/MM2_d
+ N_XI0/XI7/XI8/NET33_XI0/XI7/XI8/MM2_g N_VSS_XI0/XI7/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM3 N_XI0/XI7/XI8/NET33_XI0/XI7/XI8/MM3_d
+ N_WL<10>_XI0/XI7/XI8/MM3_g N_BLN<7>_XI0/XI7/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM0 N_XI0/XI7/XI8/NET34_XI0/XI7/XI8/MM0_d
+ N_WL<10>_XI0/XI7/XI8/MM0_g N_BL<7>_XI0/XI7/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM1 N_XI0/XI7/XI8/NET33_XI0/XI7/XI8/MM1_d
+ N_XI0/XI7/XI8/NET34_XI0/XI7/XI8/MM1_g N_VSS_XI0/XI7/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM9 N_XI0/XI7/XI8/NET36_XI0/XI7/XI8/MM9_d
+ N_WL<11>_XI0/XI7/XI8/MM9_g N_BL<7>_XI0/XI7/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM6 N_XI0/XI7/XI8/NET35_XI0/XI7/XI8/MM6_d
+ N_XI0/XI7/XI8/NET36_XI0/XI7/XI8/MM6_g N_VSS_XI0/XI7/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM7 N_XI0/XI7/XI8/NET36_XI0/XI7/XI8/MM7_d
+ N_XI0/XI7/XI8/NET35_XI0/XI7/XI8/MM7_g N_VSS_XI0/XI7/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM8 N_XI0/XI7/XI8/NET35_XI0/XI7/XI8/MM8_d
+ N_WL<11>_XI0/XI7/XI8/MM8_g N_BLN<7>_XI0/XI7/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI8/MM5 N_XI0/XI7/XI8/NET34_XI0/XI7/XI8/MM5_d
+ N_XI0/XI7/XI8/NET33_XI0/XI7/XI8/MM5_g N_VDD_XI0/XI7/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI8/MM4 N_XI0/XI7/XI8/NET33_XI0/XI7/XI8/MM4_d
+ N_XI0/XI7/XI8/NET34_XI0/XI7/XI8/MM4_g N_VDD_XI0/XI7/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI8/MM10 N_XI0/XI7/XI8/NET35_XI0/XI7/XI8/MM10_d
+ N_XI0/XI7/XI8/NET36_XI0/XI7/XI8/MM10_g N_VDD_XI0/XI7/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI8/MM11 N_XI0/XI7/XI8/NET36_XI0/XI7/XI8/MM11_d
+ N_XI0/XI7/XI8/NET35_XI0/XI7/XI8/MM11_g N_VDD_XI0/XI7/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI9/MM2 N_XI0/XI7/XI9/NET34_XI0/XI7/XI9/MM2_d
+ N_XI0/XI7/XI9/NET33_XI0/XI7/XI9/MM2_g N_VSS_XI0/XI7/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM3 N_XI0/XI7/XI9/NET33_XI0/XI7/XI9/MM3_d
+ N_WL<10>_XI0/XI7/XI9/MM3_g N_BLN<6>_XI0/XI7/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM0 N_XI0/XI7/XI9/NET34_XI0/XI7/XI9/MM0_d
+ N_WL<10>_XI0/XI7/XI9/MM0_g N_BL<6>_XI0/XI7/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM1 N_XI0/XI7/XI9/NET33_XI0/XI7/XI9/MM1_d
+ N_XI0/XI7/XI9/NET34_XI0/XI7/XI9/MM1_g N_VSS_XI0/XI7/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM9 N_XI0/XI7/XI9/NET36_XI0/XI7/XI9/MM9_d
+ N_WL<11>_XI0/XI7/XI9/MM9_g N_BL<6>_XI0/XI7/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM6 N_XI0/XI7/XI9/NET35_XI0/XI7/XI9/MM6_d
+ N_XI0/XI7/XI9/NET36_XI0/XI7/XI9/MM6_g N_VSS_XI0/XI7/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM7 N_XI0/XI7/XI9/NET36_XI0/XI7/XI9/MM7_d
+ N_XI0/XI7/XI9/NET35_XI0/XI7/XI9/MM7_g N_VSS_XI0/XI7/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM8 N_XI0/XI7/XI9/NET35_XI0/XI7/XI9/MM8_d
+ N_WL<11>_XI0/XI7/XI9/MM8_g N_BLN<6>_XI0/XI7/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI9/MM5 N_XI0/XI7/XI9/NET34_XI0/XI7/XI9/MM5_d
+ N_XI0/XI7/XI9/NET33_XI0/XI7/XI9/MM5_g N_VDD_XI0/XI7/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI9/MM4 N_XI0/XI7/XI9/NET33_XI0/XI7/XI9/MM4_d
+ N_XI0/XI7/XI9/NET34_XI0/XI7/XI9/MM4_g N_VDD_XI0/XI7/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI9/MM10 N_XI0/XI7/XI9/NET35_XI0/XI7/XI9/MM10_d
+ N_XI0/XI7/XI9/NET36_XI0/XI7/XI9/MM10_g N_VDD_XI0/XI7/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI9/MM11 N_XI0/XI7/XI9/NET36_XI0/XI7/XI9/MM11_d
+ N_XI0/XI7/XI9/NET35_XI0/XI7/XI9/MM11_g N_VDD_XI0/XI7/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI10/MM2 N_XI0/XI7/XI10/NET34_XI0/XI7/XI10/MM2_d
+ N_XI0/XI7/XI10/NET33_XI0/XI7/XI10/MM2_g N_VSS_XI0/XI7/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM3 N_XI0/XI7/XI10/NET33_XI0/XI7/XI10/MM3_d
+ N_WL<10>_XI0/XI7/XI10/MM3_g N_BLN<5>_XI0/XI7/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM0 N_XI0/XI7/XI10/NET34_XI0/XI7/XI10/MM0_d
+ N_WL<10>_XI0/XI7/XI10/MM0_g N_BL<5>_XI0/XI7/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM1 N_XI0/XI7/XI10/NET33_XI0/XI7/XI10/MM1_d
+ N_XI0/XI7/XI10/NET34_XI0/XI7/XI10/MM1_g N_VSS_XI0/XI7/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM9 N_XI0/XI7/XI10/NET36_XI0/XI7/XI10/MM9_d
+ N_WL<11>_XI0/XI7/XI10/MM9_g N_BL<5>_XI0/XI7/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM6 N_XI0/XI7/XI10/NET35_XI0/XI7/XI10/MM6_d
+ N_XI0/XI7/XI10/NET36_XI0/XI7/XI10/MM6_g N_VSS_XI0/XI7/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM7 N_XI0/XI7/XI10/NET36_XI0/XI7/XI10/MM7_d
+ N_XI0/XI7/XI10/NET35_XI0/XI7/XI10/MM7_g N_VSS_XI0/XI7/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM8 N_XI0/XI7/XI10/NET35_XI0/XI7/XI10/MM8_d
+ N_WL<11>_XI0/XI7/XI10/MM8_g N_BLN<5>_XI0/XI7/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI10/MM5 N_XI0/XI7/XI10/NET34_XI0/XI7/XI10/MM5_d
+ N_XI0/XI7/XI10/NET33_XI0/XI7/XI10/MM5_g N_VDD_XI0/XI7/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI10/MM4 N_XI0/XI7/XI10/NET33_XI0/XI7/XI10/MM4_d
+ N_XI0/XI7/XI10/NET34_XI0/XI7/XI10/MM4_g N_VDD_XI0/XI7/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI10/MM10 N_XI0/XI7/XI10/NET35_XI0/XI7/XI10/MM10_d
+ N_XI0/XI7/XI10/NET36_XI0/XI7/XI10/MM10_g N_VDD_XI0/XI7/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI10/MM11 N_XI0/XI7/XI10/NET36_XI0/XI7/XI10/MM11_d
+ N_XI0/XI7/XI10/NET35_XI0/XI7/XI10/MM11_g N_VDD_XI0/XI7/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI11/MM2 N_XI0/XI7/XI11/NET34_XI0/XI7/XI11/MM2_d
+ N_XI0/XI7/XI11/NET33_XI0/XI7/XI11/MM2_g N_VSS_XI0/XI7/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM3 N_XI0/XI7/XI11/NET33_XI0/XI7/XI11/MM3_d
+ N_WL<10>_XI0/XI7/XI11/MM3_g N_BLN<4>_XI0/XI7/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM0 N_XI0/XI7/XI11/NET34_XI0/XI7/XI11/MM0_d
+ N_WL<10>_XI0/XI7/XI11/MM0_g N_BL<4>_XI0/XI7/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM1 N_XI0/XI7/XI11/NET33_XI0/XI7/XI11/MM1_d
+ N_XI0/XI7/XI11/NET34_XI0/XI7/XI11/MM1_g N_VSS_XI0/XI7/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM9 N_XI0/XI7/XI11/NET36_XI0/XI7/XI11/MM9_d
+ N_WL<11>_XI0/XI7/XI11/MM9_g N_BL<4>_XI0/XI7/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM6 N_XI0/XI7/XI11/NET35_XI0/XI7/XI11/MM6_d
+ N_XI0/XI7/XI11/NET36_XI0/XI7/XI11/MM6_g N_VSS_XI0/XI7/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM7 N_XI0/XI7/XI11/NET36_XI0/XI7/XI11/MM7_d
+ N_XI0/XI7/XI11/NET35_XI0/XI7/XI11/MM7_g N_VSS_XI0/XI7/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM8 N_XI0/XI7/XI11/NET35_XI0/XI7/XI11/MM8_d
+ N_WL<11>_XI0/XI7/XI11/MM8_g N_BLN<4>_XI0/XI7/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI11/MM5 N_XI0/XI7/XI11/NET34_XI0/XI7/XI11/MM5_d
+ N_XI0/XI7/XI11/NET33_XI0/XI7/XI11/MM5_g N_VDD_XI0/XI7/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI11/MM4 N_XI0/XI7/XI11/NET33_XI0/XI7/XI11/MM4_d
+ N_XI0/XI7/XI11/NET34_XI0/XI7/XI11/MM4_g N_VDD_XI0/XI7/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI11/MM10 N_XI0/XI7/XI11/NET35_XI0/XI7/XI11/MM10_d
+ N_XI0/XI7/XI11/NET36_XI0/XI7/XI11/MM10_g N_VDD_XI0/XI7/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI11/MM11 N_XI0/XI7/XI11/NET36_XI0/XI7/XI11/MM11_d
+ N_XI0/XI7/XI11/NET35_XI0/XI7/XI11/MM11_g N_VDD_XI0/XI7/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI12/MM2 N_XI0/XI7/XI12/NET34_XI0/XI7/XI12/MM2_d
+ N_XI0/XI7/XI12/NET33_XI0/XI7/XI12/MM2_g N_VSS_XI0/XI7/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM3 N_XI0/XI7/XI12/NET33_XI0/XI7/XI12/MM3_d
+ N_WL<10>_XI0/XI7/XI12/MM3_g N_BLN<3>_XI0/XI7/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM0 N_XI0/XI7/XI12/NET34_XI0/XI7/XI12/MM0_d
+ N_WL<10>_XI0/XI7/XI12/MM0_g N_BL<3>_XI0/XI7/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM1 N_XI0/XI7/XI12/NET33_XI0/XI7/XI12/MM1_d
+ N_XI0/XI7/XI12/NET34_XI0/XI7/XI12/MM1_g N_VSS_XI0/XI7/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM9 N_XI0/XI7/XI12/NET36_XI0/XI7/XI12/MM9_d
+ N_WL<11>_XI0/XI7/XI12/MM9_g N_BL<3>_XI0/XI7/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM6 N_XI0/XI7/XI12/NET35_XI0/XI7/XI12/MM6_d
+ N_XI0/XI7/XI12/NET36_XI0/XI7/XI12/MM6_g N_VSS_XI0/XI7/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM7 N_XI0/XI7/XI12/NET36_XI0/XI7/XI12/MM7_d
+ N_XI0/XI7/XI12/NET35_XI0/XI7/XI12/MM7_g N_VSS_XI0/XI7/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM8 N_XI0/XI7/XI12/NET35_XI0/XI7/XI12/MM8_d
+ N_WL<11>_XI0/XI7/XI12/MM8_g N_BLN<3>_XI0/XI7/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI12/MM5 N_XI0/XI7/XI12/NET34_XI0/XI7/XI12/MM5_d
+ N_XI0/XI7/XI12/NET33_XI0/XI7/XI12/MM5_g N_VDD_XI0/XI7/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI12/MM4 N_XI0/XI7/XI12/NET33_XI0/XI7/XI12/MM4_d
+ N_XI0/XI7/XI12/NET34_XI0/XI7/XI12/MM4_g N_VDD_XI0/XI7/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI12/MM10 N_XI0/XI7/XI12/NET35_XI0/XI7/XI12/MM10_d
+ N_XI0/XI7/XI12/NET36_XI0/XI7/XI12/MM10_g N_VDD_XI0/XI7/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI12/MM11 N_XI0/XI7/XI12/NET36_XI0/XI7/XI12/MM11_d
+ N_XI0/XI7/XI12/NET35_XI0/XI7/XI12/MM11_g N_VDD_XI0/XI7/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI13/MM2 N_XI0/XI7/XI13/NET34_XI0/XI7/XI13/MM2_d
+ N_XI0/XI7/XI13/NET33_XI0/XI7/XI13/MM2_g N_VSS_XI0/XI7/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM3 N_XI0/XI7/XI13/NET33_XI0/XI7/XI13/MM3_d
+ N_WL<10>_XI0/XI7/XI13/MM3_g N_BLN<2>_XI0/XI7/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM0 N_XI0/XI7/XI13/NET34_XI0/XI7/XI13/MM0_d
+ N_WL<10>_XI0/XI7/XI13/MM0_g N_BL<2>_XI0/XI7/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM1 N_XI0/XI7/XI13/NET33_XI0/XI7/XI13/MM1_d
+ N_XI0/XI7/XI13/NET34_XI0/XI7/XI13/MM1_g N_VSS_XI0/XI7/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM9 N_XI0/XI7/XI13/NET36_XI0/XI7/XI13/MM9_d
+ N_WL<11>_XI0/XI7/XI13/MM9_g N_BL<2>_XI0/XI7/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM6 N_XI0/XI7/XI13/NET35_XI0/XI7/XI13/MM6_d
+ N_XI0/XI7/XI13/NET36_XI0/XI7/XI13/MM6_g N_VSS_XI0/XI7/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM7 N_XI0/XI7/XI13/NET36_XI0/XI7/XI13/MM7_d
+ N_XI0/XI7/XI13/NET35_XI0/XI7/XI13/MM7_g N_VSS_XI0/XI7/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM8 N_XI0/XI7/XI13/NET35_XI0/XI7/XI13/MM8_d
+ N_WL<11>_XI0/XI7/XI13/MM8_g N_BLN<2>_XI0/XI7/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI13/MM5 N_XI0/XI7/XI13/NET34_XI0/XI7/XI13/MM5_d
+ N_XI0/XI7/XI13/NET33_XI0/XI7/XI13/MM5_g N_VDD_XI0/XI7/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI13/MM4 N_XI0/XI7/XI13/NET33_XI0/XI7/XI13/MM4_d
+ N_XI0/XI7/XI13/NET34_XI0/XI7/XI13/MM4_g N_VDD_XI0/XI7/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI13/MM10 N_XI0/XI7/XI13/NET35_XI0/XI7/XI13/MM10_d
+ N_XI0/XI7/XI13/NET36_XI0/XI7/XI13/MM10_g N_VDD_XI0/XI7/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI13/MM11 N_XI0/XI7/XI13/NET36_XI0/XI7/XI13/MM11_d
+ N_XI0/XI7/XI13/NET35_XI0/XI7/XI13/MM11_g N_VDD_XI0/XI7/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI14/MM2 N_XI0/XI7/XI14/NET34_XI0/XI7/XI14/MM2_d
+ N_XI0/XI7/XI14/NET33_XI0/XI7/XI14/MM2_g N_VSS_XI0/XI7/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM3 N_XI0/XI7/XI14/NET33_XI0/XI7/XI14/MM3_d
+ N_WL<10>_XI0/XI7/XI14/MM3_g N_BLN<1>_XI0/XI7/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM0 N_XI0/XI7/XI14/NET34_XI0/XI7/XI14/MM0_d
+ N_WL<10>_XI0/XI7/XI14/MM0_g N_BL<1>_XI0/XI7/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM1 N_XI0/XI7/XI14/NET33_XI0/XI7/XI14/MM1_d
+ N_XI0/XI7/XI14/NET34_XI0/XI7/XI14/MM1_g N_VSS_XI0/XI7/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM9 N_XI0/XI7/XI14/NET36_XI0/XI7/XI14/MM9_d
+ N_WL<11>_XI0/XI7/XI14/MM9_g N_BL<1>_XI0/XI7/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM6 N_XI0/XI7/XI14/NET35_XI0/XI7/XI14/MM6_d
+ N_XI0/XI7/XI14/NET36_XI0/XI7/XI14/MM6_g N_VSS_XI0/XI7/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM7 N_XI0/XI7/XI14/NET36_XI0/XI7/XI14/MM7_d
+ N_XI0/XI7/XI14/NET35_XI0/XI7/XI14/MM7_g N_VSS_XI0/XI7/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM8 N_XI0/XI7/XI14/NET35_XI0/XI7/XI14/MM8_d
+ N_WL<11>_XI0/XI7/XI14/MM8_g N_BLN<1>_XI0/XI7/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI14/MM5 N_XI0/XI7/XI14/NET34_XI0/XI7/XI14/MM5_d
+ N_XI0/XI7/XI14/NET33_XI0/XI7/XI14/MM5_g N_VDD_XI0/XI7/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI14/MM4 N_XI0/XI7/XI14/NET33_XI0/XI7/XI14/MM4_d
+ N_XI0/XI7/XI14/NET34_XI0/XI7/XI14/MM4_g N_VDD_XI0/XI7/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI14/MM10 N_XI0/XI7/XI14/NET35_XI0/XI7/XI14/MM10_d
+ N_XI0/XI7/XI14/NET36_XI0/XI7/XI14/MM10_g N_VDD_XI0/XI7/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI14/MM11 N_XI0/XI7/XI14/NET36_XI0/XI7/XI14/MM11_d
+ N_XI0/XI7/XI14/NET35_XI0/XI7/XI14/MM11_g N_VDD_XI0/XI7/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI15/MM2 N_XI0/XI7/XI15/NET34_XI0/XI7/XI15/MM2_d
+ N_XI0/XI7/XI15/NET33_XI0/XI7/XI15/MM2_g N_VSS_XI0/XI7/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM3 N_XI0/XI7/XI15/NET33_XI0/XI7/XI15/MM3_d
+ N_WL<10>_XI0/XI7/XI15/MM3_g N_BLN<0>_XI0/XI7/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM0 N_XI0/XI7/XI15/NET34_XI0/XI7/XI15/MM0_d
+ N_WL<10>_XI0/XI7/XI15/MM0_g N_BL<0>_XI0/XI7/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM1 N_XI0/XI7/XI15/NET33_XI0/XI7/XI15/MM1_d
+ N_XI0/XI7/XI15/NET34_XI0/XI7/XI15/MM1_g N_VSS_XI0/XI7/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM9 N_XI0/XI7/XI15/NET36_XI0/XI7/XI15/MM9_d
+ N_WL<11>_XI0/XI7/XI15/MM9_g N_BL<0>_XI0/XI7/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM6 N_XI0/XI7/XI15/NET35_XI0/XI7/XI15/MM6_d
+ N_XI0/XI7/XI15/NET36_XI0/XI7/XI15/MM6_g N_VSS_XI0/XI7/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM7 N_XI0/XI7/XI15/NET36_XI0/XI7/XI15/MM7_d
+ N_XI0/XI7/XI15/NET35_XI0/XI7/XI15/MM7_g N_VSS_XI0/XI7/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM8 N_XI0/XI7/XI15/NET35_XI0/XI7/XI15/MM8_d
+ N_WL<11>_XI0/XI7/XI15/MM8_g N_BLN<0>_XI0/XI7/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/XI15/MM5 N_XI0/XI7/XI15/NET34_XI0/XI7/XI15/MM5_d
+ N_XI0/XI7/XI15/NET33_XI0/XI7/XI15/MM5_g N_VDD_XI0/XI7/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI15/MM4 N_XI0/XI7/XI15/NET33_XI0/XI7/XI15/MM4_d
+ N_XI0/XI7/XI15/NET34_XI0/XI7/XI15/MM4_g N_VDD_XI0/XI7/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI15/MM10 N_XI0/XI7/XI15/NET35_XI0/XI7/XI15/MM10_d
+ N_XI0/XI7/XI15/NET36_XI0/XI7/XI15/MM10_g N_VDD_XI0/XI7/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/XI15/MM11 N_XI0/XI7/XI15/NET36_XI0/XI7/XI15/MM11_d
+ N_XI0/XI7/XI15/NET35_XI0/XI7/XI15/MM11_g N_VDD_XI0/XI7/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI0/MM2 N_XI0/XI8/XI0/NET34_XI0/XI8/XI0/MM2_d
+ N_XI0/XI8/XI0/NET33_XI0/XI8/XI0/MM2_g N_VSS_XI0/XI8/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM3 N_XI0/XI8/XI0/NET33_XI0/XI8/XI0/MM3_d
+ N_WL<12>_XI0/XI8/XI0/MM3_g N_BLN<15>_XI0/XI8/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM0 N_XI0/XI8/XI0/NET34_XI0/XI8/XI0/MM0_d
+ N_WL<12>_XI0/XI8/XI0/MM0_g N_BL<15>_XI0/XI8/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM1 N_XI0/XI8/XI0/NET33_XI0/XI8/XI0/MM1_d
+ N_XI0/XI8/XI0/NET34_XI0/XI8/XI0/MM1_g N_VSS_XI0/XI8/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM9 N_XI0/XI8/XI0/NET36_XI0/XI8/XI0/MM9_d
+ N_WL<13>_XI0/XI8/XI0/MM9_g N_BL<15>_XI0/XI8/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM6 N_XI0/XI8/XI0/NET35_XI0/XI8/XI0/MM6_d
+ N_XI0/XI8/XI0/NET36_XI0/XI8/XI0/MM6_g N_VSS_XI0/XI8/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM7 N_XI0/XI8/XI0/NET36_XI0/XI8/XI0/MM7_d
+ N_XI0/XI8/XI0/NET35_XI0/XI8/XI0/MM7_g N_VSS_XI0/XI8/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM8 N_XI0/XI8/XI0/NET35_XI0/XI8/XI0/MM8_d
+ N_WL<13>_XI0/XI8/XI0/MM8_g N_BLN<15>_XI0/XI8/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI0/MM5 N_XI0/XI8/XI0/NET34_XI0/XI8/XI0/MM5_d
+ N_XI0/XI8/XI0/NET33_XI0/XI8/XI0/MM5_g N_VDD_XI0/XI8/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI0/MM4 N_XI0/XI8/XI0/NET33_XI0/XI8/XI0/MM4_d
+ N_XI0/XI8/XI0/NET34_XI0/XI8/XI0/MM4_g N_VDD_XI0/XI8/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI0/MM10 N_XI0/XI8/XI0/NET35_XI0/XI8/XI0/MM10_d
+ N_XI0/XI8/XI0/NET36_XI0/XI8/XI0/MM10_g N_VDD_XI0/XI8/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI0/MM11 N_XI0/XI8/XI0/NET36_XI0/XI8/XI0/MM11_d
+ N_XI0/XI8/XI0/NET35_XI0/XI8/XI0/MM11_g N_VDD_XI0/XI8/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI1/MM2 N_XI0/XI8/XI1/NET34_XI0/XI8/XI1/MM2_d
+ N_XI0/XI8/XI1/NET33_XI0/XI8/XI1/MM2_g N_VSS_XI0/XI8/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM3 N_XI0/XI8/XI1/NET33_XI0/XI8/XI1/MM3_d
+ N_WL<12>_XI0/XI8/XI1/MM3_g N_BLN<14>_XI0/XI8/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM0 N_XI0/XI8/XI1/NET34_XI0/XI8/XI1/MM0_d
+ N_WL<12>_XI0/XI8/XI1/MM0_g N_BL<14>_XI0/XI8/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM1 N_XI0/XI8/XI1/NET33_XI0/XI8/XI1/MM1_d
+ N_XI0/XI8/XI1/NET34_XI0/XI8/XI1/MM1_g N_VSS_XI0/XI8/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM9 N_XI0/XI8/XI1/NET36_XI0/XI8/XI1/MM9_d
+ N_WL<13>_XI0/XI8/XI1/MM9_g N_BL<14>_XI0/XI8/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM6 N_XI0/XI8/XI1/NET35_XI0/XI8/XI1/MM6_d
+ N_XI0/XI8/XI1/NET36_XI0/XI8/XI1/MM6_g N_VSS_XI0/XI8/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM7 N_XI0/XI8/XI1/NET36_XI0/XI8/XI1/MM7_d
+ N_XI0/XI8/XI1/NET35_XI0/XI8/XI1/MM7_g N_VSS_XI0/XI8/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM8 N_XI0/XI8/XI1/NET35_XI0/XI8/XI1/MM8_d
+ N_WL<13>_XI0/XI8/XI1/MM8_g N_BLN<14>_XI0/XI8/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI1/MM5 N_XI0/XI8/XI1/NET34_XI0/XI8/XI1/MM5_d
+ N_XI0/XI8/XI1/NET33_XI0/XI8/XI1/MM5_g N_VDD_XI0/XI8/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI1/MM4 N_XI0/XI8/XI1/NET33_XI0/XI8/XI1/MM4_d
+ N_XI0/XI8/XI1/NET34_XI0/XI8/XI1/MM4_g N_VDD_XI0/XI8/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI1/MM10 N_XI0/XI8/XI1/NET35_XI0/XI8/XI1/MM10_d
+ N_XI0/XI8/XI1/NET36_XI0/XI8/XI1/MM10_g N_VDD_XI0/XI8/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI1/MM11 N_XI0/XI8/XI1/NET36_XI0/XI8/XI1/MM11_d
+ N_XI0/XI8/XI1/NET35_XI0/XI8/XI1/MM11_g N_VDD_XI0/XI8/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI2/MM2 N_XI0/XI8/XI2/NET34_XI0/XI8/XI2/MM2_d
+ N_XI0/XI8/XI2/NET33_XI0/XI8/XI2/MM2_g N_VSS_XI0/XI8/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM3 N_XI0/XI8/XI2/NET33_XI0/XI8/XI2/MM3_d
+ N_WL<12>_XI0/XI8/XI2/MM3_g N_BLN<13>_XI0/XI8/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM0 N_XI0/XI8/XI2/NET34_XI0/XI8/XI2/MM0_d
+ N_WL<12>_XI0/XI8/XI2/MM0_g N_BL<13>_XI0/XI8/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM1 N_XI0/XI8/XI2/NET33_XI0/XI8/XI2/MM1_d
+ N_XI0/XI8/XI2/NET34_XI0/XI8/XI2/MM1_g N_VSS_XI0/XI8/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM9 N_XI0/XI8/XI2/NET36_XI0/XI8/XI2/MM9_d
+ N_WL<13>_XI0/XI8/XI2/MM9_g N_BL<13>_XI0/XI8/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM6 N_XI0/XI8/XI2/NET35_XI0/XI8/XI2/MM6_d
+ N_XI0/XI8/XI2/NET36_XI0/XI8/XI2/MM6_g N_VSS_XI0/XI8/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM7 N_XI0/XI8/XI2/NET36_XI0/XI8/XI2/MM7_d
+ N_XI0/XI8/XI2/NET35_XI0/XI8/XI2/MM7_g N_VSS_XI0/XI8/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM8 N_XI0/XI8/XI2/NET35_XI0/XI8/XI2/MM8_d
+ N_WL<13>_XI0/XI8/XI2/MM8_g N_BLN<13>_XI0/XI8/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI2/MM5 N_XI0/XI8/XI2/NET34_XI0/XI8/XI2/MM5_d
+ N_XI0/XI8/XI2/NET33_XI0/XI8/XI2/MM5_g N_VDD_XI0/XI8/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI2/MM4 N_XI0/XI8/XI2/NET33_XI0/XI8/XI2/MM4_d
+ N_XI0/XI8/XI2/NET34_XI0/XI8/XI2/MM4_g N_VDD_XI0/XI8/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI2/MM10 N_XI0/XI8/XI2/NET35_XI0/XI8/XI2/MM10_d
+ N_XI0/XI8/XI2/NET36_XI0/XI8/XI2/MM10_g N_VDD_XI0/XI8/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI2/MM11 N_XI0/XI8/XI2/NET36_XI0/XI8/XI2/MM11_d
+ N_XI0/XI8/XI2/NET35_XI0/XI8/XI2/MM11_g N_VDD_XI0/XI8/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI3/MM2 N_XI0/XI8/XI3/NET34_XI0/XI8/XI3/MM2_d
+ N_XI0/XI8/XI3/NET33_XI0/XI8/XI3/MM2_g N_VSS_XI0/XI8/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM3 N_XI0/XI8/XI3/NET33_XI0/XI8/XI3/MM3_d
+ N_WL<12>_XI0/XI8/XI3/MM3_g N_BLN<12>_XI0/XI8/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM0 N_XI0/XI8/XI3/NET34_XI0/XI8/XI3/MM0_d
+ N_WL<12>_XI0/XI8/XI3/MM0_g N_BL<12>_XI0/XI8/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM1 N_XI0/XI8/XI3/NET33_XI0/XI8/XI3/MM1_d
+ N_XI0/XI8/XI3/NET34_XI0/XI8/XI3/MM1_g N_VSS_XI0/XI8/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM9 N_XI0/XI8/XI3/NET36_XI0/XI8/XI3/MM9_d
+ N_WL<13>_XI0/XI8/XI3/MM9_g N_BL<12>_XI0/XI8/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM6 N_XI0/XI8/XI3/NET35_XI0/XI8/XI3/MM6_d
+ N_XI0/XI8/XI3/NET36_XI0/XI8/XI3/MM6_g N_VSS_XI0/XI8/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM7 N_XI0/XI8/XI3/NET36_XI0/XI8/XI3/MM7_d
+ N_XI0/XI8/XI3/NET35_XI0/XI8/XI3/MM7_g N_VSS_XI0/XI8/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM8 N_XI0/XI8/XI3/NET35_XI0/XI8/XI3/MM8_d
+ N_WL<13>_XI0/XI8/XI3/MM8_g N_BLN<12>_XI0/XI8/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI3/MM5 N_XI0/XI8/XI3/NET34_XI0/XI8/XI3/MM5_d
+ N_XI0/XI8/XI3/NET33_XI0/XI8/XI3/MM5_g N_VDD_XI0/XI8/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI3/MM4 N_XI0/XI8/XI3/NET33_XI0/XI8/XI3/MM4_d
+ N_XI0/XI8/XI3/NET34_XI0/XI8/XI3/MM4_g N_VDD_XI0/XI8/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI3/MM10 N_XI0/XI8/XI3/NET35_XI0/XI8/XI3/MM10_d
+ N_XI0/XI8/XI3/NET36_XI0/XI8/XI3/MM10_g N_VDD_XI0/XI8/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI3/MM11 N_XI0/XI8/XI3/NET36_XI0/XI8/XI3/MM11_d
+ N_XI0/XI8/XI3/NET35_XI0/XI8/XI3/MM11_g N_VDD_XI0/XI8/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI4/MM2 N_XI0/XI8/XI4/NET34_XI0/XI8/XI4/MM2_d
+ N_XI0/XI8/XI4/NET33_XI0/XI8/XI4/MM2_g N_VSS_XI0/XI8/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM3 N_XI0/XI8/XI4/NET33_XI0/XI8/XI4/MM3_d
+ N_WL<12>_XI0/XI8/XI4/MM3_g N_BLN<11>_XI0/XI8/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM0 N_XI0/XI8/XI4/NET34_XI0/XI8/XI4/MM0_d
+ N_WL<12>_XI0/XI8/XI4/MM0_g N_BL<11>_XI0/XI8/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM1 N_XI0/XI8/XI4/NET33_XI0/XI8/XI4/MM1_d
+ N_XI0/XI8/XI4/NET34_XI0/XI8/XI4/MM1_g N_VSS_XI0/XI8/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM9 N_XI0/XI8/XI4/NET36_XI0/XI8/XI4/MM9_d
+ N_WL<13>_XI0/XI8/XI4/MM9_g N_BL<11>_XI0/XI8/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM6 N_XI0/XI8/XI4/NET35_XI0/XI8/XI4/MM6_d
+ N_XI0/XI8/XI4/NET36_XI0/XI8/XI4/MM6_g N_VSS_XI0/XI8/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM7 N_XI0/XI8/XI4/NET36_XI0/XI8/XI4/MM7_d
+ N_XI0/XI8/XI4/NET35_XI0/XI8/XI4/MM7_g N_VSS_XI0/XI8/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM8 N_XI0/XI8/XI4/NET35_XI0/XI8/XI4/MM8_d
+ N_WL<13>_XI0/XI8/XI4/MM8_g N_BLN<11>_XI0/XI8/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI4/MM5 N_XI0/XI8/XI4/NET34_XI0/XI8/XI4/MM5_d
+ N_XI0/XI8/XI4/NET33_XI0/XI8/XI4/MM5_g N_VDD_XI0/XI8/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI4/MM4 N_XI0/XI8/XI4/NET33_XI0/XI8/XI4/MM4_d
+ N_XI0/XI8/XI4/NET34_XI0/XI8/XI4/MM4_g N_VDD_XI0/XI8/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI4/MM10 N_XI0/XI8/XI4/NET35_XI0/XI8/XI4/MM10_d
+ N_XI0/XI8/XI4/NET36_XI0/XI8/XI4/MM10_g N_VDD_XI0/XI8/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI4/MM11 N_XI0/XI8/XI4/NET36_XI0/XI8/XI4/MM11_d
+ N_XI0/XI8/XI4/NET35_XI0/XI8/XI4/MM11_g N_VDD_XI0/XI8/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI5/MM2 N_XI0/XI8/XI5/NET34_XI0/XI8/XI5/MM2_d
+ N_XI0/XI8/XI5/NET33_XI0/XI8/XI5/MM2_g N_VSS_XI0/XI8/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM3 N_XI0/XI8/XI5/NET33_XI0/XI8/XI5/MM3_d
+ N_WL<12>_XI0/XI8/XI5/MM3_g N_BLN<10>_XI0/XI8/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM0 N_XI0/XI8/XI5/NET34_XI0/XI8/XI5/MM0_d
+ N_WL<12>_XI0/XI8/XI5/MM0_g N_BL<10>_XI0/XI8/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM1 N_XI0/XI8/XI5/NET33_XI0/XI8/XI5/MM1_d
+ N_XI0/XI8/XI5/NET34_XI0/XI8/XI5/MM1_g N_VSS_XI0/XI8/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM9 N_XI0/XI8/XI5/NET36_XI0/XI8/XI5/MM9_d
+ N_WL<13>_XI0/XI8/XI5/MM9_g N_BL<10>_XI0/XI8/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM6 N_XI0/XI8/XI5/NET35_XI0/XI8/XI5/MM6_d
+ N_XI0/XI8/XI5/NET36_XI0/XI8/XI5/MM6_g N_VSS_XI0/XI8/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM7 N_XI0/XI8/XI5/NET36_XI0/XI8/XI5/MM7_d
+ N_XI0/XI8/XI5/NET35_XI0/XI8/XI5/MM7_g N_VSS_XI0/XI8/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM8 N_XI0/XI8/XI5/NET35_XI0/XI8/XI5/MM8_d
+ N_WL<13>_XI0/XI8/XI5/MM8_g N_BLN<10>_XI0/XI8/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI5/MM5 N_XI0/XI8/XI5/NET34_XI0/XI8/XI5/MM5_d
+ N_XI0/XI8/XI5/NET33_XI0/XI8/XI5/MM5_g N_VDD_XI0/XI8/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI5/MM4 N_XI0/XI8/XI5/NET33_XI0/XI8/XI5/MM4_d
+ N_XI0/XI8/XI5/NET34_XI0/XI8/XI5/MM4_g N_VDD_XI0/XI8/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI5/MM10 N_XI0/XI8/XI5/NET35_XI0/XI8/XI5/MM10_d
+ N_XI0/XI8/XI5/NET36_XI0/XI8/XI5/MM10_g N_VDD_XI0/XI8/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI5/MM11 N_XI0/XI8/XI5/NET36_XI0/XI8/XI5/MM11_d
+ N_XI0/XI8/XI5/NET35_XI0/XI8/XI5/MM11_g N_VDD_XI0/XI8/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI6/MM2 N_XI0/XI8/XI6/NET34_XI0/XI8/XI6/MM2_d
+ N_XI0/XI8/XI6/NET33_XI0/XI8/XI6/MM2_g N_VSS_XI0/XI8/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM3 N_XI0/XI8/XI6/NET33_XI0/XI8/XI6/MM3_d
+ N_WL<12>_XI0/XI8/XI6/MM3_g N_BLN<9>_XI0/XI8/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM0 N_XI0/XI8/XI6/NET34_XI0/XI8/XI6/MM0_d
+ N_WL<12>_XI0/XI8/XI6/MM0_g N_BL<9>_XI0/XI8/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM1 N_XI0/XI8/XI6/NET33_XI0/XI8/XI6/MM1_d
+ N_XI0/XI8/XI6/NET34_XI0/XI8/XI6/MM1_g N_VSS_XI0/XI8/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM9 N_XI0/XI8/XI6/NET36_XI0/XI8/XI6/MM9_d
+ N_WL<13>_XI0/XI8/XI6/MM9_g N_BL<9>_XI0/XI8/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM6 N_XI0/XI8/XI6/NET35_XI0/XI8/XI6/MM6_d
+ N_XI0/XI8/XI6/NET36_XI0/XI8/XI6/MM6_g N_VSS_XI0/XI8/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM7 N_XI0/XI8/XI6/NET36_XI0/XI8/XI6/MM7_d
+ N_XI0/XI8/XI6/NET35_XI0/XI8/XI6/MM7_g N_VSS_XI0/XI8/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM8 N_XI0/XI8/XI6/NET35_XI0/XI8/XI6/MM8_d
+ N_WL<13>_XI0/XI8/XI6/MM8_g N_BLN<9>_XI0/XI8/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI6/MM5 N_XI0/XI8/XI6/NET34_XI0/XI8/XI6/MM5_d
+ N_XI0/XI8/XI6/NET33_XI0/XI8/XI6/MM5_g N_VDD_XI0/XI8/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI6/MM4 N_XI0/XI8/XI6/NET33_XI0/XI8/XI6/MM4_d
+ N_XI0/XI8/XI6/NET34_XI0/XI8/XI6/MM4_g N_VDD_XI0/XI8/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI6/MM10 N_XI0/XI8/XI6/NET35_XI0/XI8/XI6/MM10_d
+ N_XI0/XI8/XI6/NET36_XI0/XI8/XI6/MM10_g N_VDD_XI0/XI8/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI6/MM11 N_XI0/XI8/XI6/NET36_XI0/XI8/XI6/MM11_d
+ N_XI0/XI8/XI6/NET35_XI0/XI8/XI6/MM11_g N_VDD_XI0/XI8/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI7/MM2 N_XI0/XI8/XI7/NET34_XI0/XI8/XI7/MM2_d
+ N_XI0/XI8/XI7/NET33_XI0/XI8/XI7/MM2_g N_VSS_XI0/XI8/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM3 N_XI0/XI8/XI7/NET33_XI0/XI8/XI7/MM3_d
+ N_WL<12>_XI0/XI8/XI7/MM3_g N_BLN<8>_XI0/XI8/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM0 N_XI0/XI8/XI7/NET34_XI0/XI8/XI7/MM0_d
+ N_WL<12>_XI0/XI8/XI7/MM0_g N_BL<8>_XI0/XI8/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM1 N_XI0/XI8/XI7/NET33_XI0/XI8/XI7/MM1_d
+ N_XI0/XI8/XI7/NET34_XI0/XI8/XI7/MM1_g N_VSS_XI0/XI8/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM9 N_XI0/XI8/XI7/NET36_XI0/XI8/XI7/MM9_d
+ N_WL<13>_XI0/XI8/XI7/MM9_g N_BL<8>_XI0/XI8/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM6 N_XI0/XI8/XI7/NET35_XI0/XI8/XI7/MM6_d
+ N_XI0/XI8/XI7/NET36_XI0/XI8/XI7/MM6_g N_VSS_XI0/XI8/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM7 N_XI0/XI8/XI7/NET36_XI0/XI8/XI7/MM7_d
+ N_XI0/XI8/XI7/NET35_XI0/XI8/XI7/MM7_g N_VSS_XI0/XI8/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM8 N_XI0/XI8/XI7/NET35_XI0/XI8/XI7/MM8_d
+ N_WL<13>_XI0/XI8/XI7/MM8_g N_BLN<8>_XI0/XI8/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI7/MM5 N_XI0/XI8/XI7/NET34_XI0/XI8/XI7/MM5_d
+ N_XI0/XI8/XI7/NET33_XI0/XI8/XI7/MM5_g N_VDD_XI0/XI8/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI7/MM4 N_XI0/XI8/XI7/NET33_XI0/XI8/XI7/MM4_d
+ N_XI0/XI8/XI7/NET34_XI0/XI8/XI7/MM4_g N_VDD_XI0/XI8/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI7/MM10 N_XI0/XI8/XI7/NET35_XI0/XI8/XI7/MM10_d
+ N_XI0/XI8/XI7/NET36_XI0/XI8/XI7/MM10_g N_VDD_XI0/XI8/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI7/MM11 N_XI0/XI8/XI7/NET36_XI0/XI8/XI7/MM11_d
+ N_XI0/XI8/XI7/NET35_XI0/XI8/XI7/MM11_g N_VDD_XI0/XI8/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI8/MM2 N_XI0/XI8/XI8/NET34_XI0/XI8/XI8/MM2_d
+ N_XI0/XI8/XI8/NET33_XI0/XI8/XI8/MM2_g N_VSS_XI0/XI8/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM3 N_XI0/XI8/XI8/NET33_XI0/XI8/XI8/MM3_d
+ N_WL<12>_XI0/XI8/XI8/MM3_g N_BLN<7>_XI0/XI8/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM0 N_XI0/XI8/XI8/NET34_XI0/XI8/XI8/MM0_d
+ N_WL<12>_XI0/XI8/XI8/MM0_g N_BL<7>_XI0/XI8/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM1 N_XI0/XI8/XI8/NET33_XI0/XI8/XI8/MM1_d
+ N_XI0/XI8/XI8/NET34_XI0/XI8/XI8/MM1_g N_VSS_XI0/XI8/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM9 N_XI0/XI8/XI8/NET36_XI0/XI8/XI8/MM9_d
+ N_WL<13>_XI0/XI8/XI8/MM9_g N_BL<7>_XI0/XI8/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM6 N_XI0/XI8/XI8/NET35_XI0/XI8/XI8/MM6_d
+ N_XI0/XI8/XI8/NET36_XI0/XI8/XI8/MM6_g N_VSS_XI0/XI8/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM7 N_XI0/XI8/XI8/NET36_XI0/XI8/XI8/MM7_d
+ N_XI0/XI8/XI8/NET35_XI0/XI8/XI8/MM7_g N_VSS_XI0/XI8/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM8 N_XI0/XI8/XI8/NET35_XI0/XI8/XI8/MM8_d
+ N_WL<13>_XI0/XI8/XI8/MM8_g N_BLN<7>_XI0/XI8/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI8/MM5 N_XI0/XI8/XI8/NET34_XI0/XI8/XI8/MM5_d
+ N_XI0/XI8/XI8/NET33_XI0/XI8/XI8/MM5_g N_VDD_XI0/XI8/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI8/MM4 N_XI0/XI8/XI8/NET33_XI0/XI8/XI8/MM4_d
+ N_XI0/XI8/XI8/NET34_XI0/XI8/XI8/MM4_g N_VDD_XI0/XI8/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI8/MM10 N_XI0/XI8/XI8/NET35_XI0/XI8/XI8/MM10_d
+ N_XI0/XI8/XI8/NET36_XI0/XI8/XI8/MM10_g N_VDD_XI0/XI8/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI8/MM11 N_XI0/XI8/XI8/NET36_XI0/XI8/XI8/MM11_d
+ N_XI0/XI8/XI8/NET35_XI0/XI8/XI8/MM11_g N_VDD_XI0/XI8/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI9/MM2 N_XI0/XI8/XI9/NET34_XI0/XI8/XI9/MM2_d
+ N_XI0/XI8/XI9/NET33_XI0/XI8/XI9/MM2_g N_VSS_XI0/XI8/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM3 N_XI0/XI8/XI9/NET33_XI0/XI8/XI9/MM3_d
+ N_WL<12>_XI0/XI8/XI9/MM3_g N_BLN<6>_XI0/XI8/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM0 N_XI0/XI8/XI9/NET34_XI0/XI8/XI9/MM0_d
+ N_WL<12>_XI0/XI8/XI9/MM0_g N_BL<6>_XI0/XI8/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM1 N_XI0/XI8/XI9/NET33_XI0/XI8/XI9/MM1_d
+ N_XI0/XI8/XI9/NET34_XI0/XI8/XI9/MM1_g N_VSS_XI0/XI8/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM9 N_XI0/XI8/XI9/NET36_XI0/XI8/XI9/MM9_d
+ N_WL<13>_XI0/XI8/XI9/MM9_g N_BL<6>_XI0/XI8/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM6 N_XI0/XI8/XI9/NET35_XI0/XI8/XI9/MM6_d
+ N_XI0/XI8/XI9/NET36_XI0/XI8/XI9/MM6_g N_VSS_XI0/XI8/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM7 N_XI0/XI8/XI9/NET36_XI0/XI8/XI9/MM7_d
+ N_XI0/XI8/XI9/NET35_XI0/XI8/XI9/MM7_g N_VSS_XI0/XI8/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM8 N_XI0/XI8/XI9/NET35_XI0/XI8/XI9/MM8_d
+ N_WL<13>_XI0/XI8/XI9/MM8_g N_BLN<6>_XI0/XI8/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI9/MM5 N_XI0/XI8/XI9/NET34_XI0/XI8/XI9/MM5_d
+ N_XI0/XI8/XI9/NET33_XI0/XI8/XI9/MM5_g N_VDD_XI0/XI8/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI9/MM4 N_XI0/XI8/XI9/NET33_XI0/XI8/XI9/MM4_d
+ N_XI0/XI8/XI9/NET34_XI0/XI8/XI9/MM4_g N_VDD_XI0/XI8/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI9/MM10 N_XI0/XI8/XI9/NET35_XI0/XI8/XI9/MM10_d
+ N_XI0/XI8/XI9/NET36_XI0/XI8/XI9/MM10_g N_VDD_XI0/XI8/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI9/MM11 N_XI0/XI8/XI9/NET36_XI0/XI8/XI9/MM11_d
+ N_XI0/XI8/XI9/NET35_XI0/XI8/XI9/MM11_g N_VDD_XI0/XI8/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI10/MM2 N_XI0/XI8/XI10/NET34_XI0/XI8/XI10/MM2_d
+ N_XI0/XI8/XI10/NET33_XI0/XI8/XI10/MM2_g N_VSS_XI0/XI8/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM3 N_XI0/XI8/XI10/NET33_XI0/XI8/XI10/MM3_d
+ N_WL<12>_XI0/XI8/XI10/MM3_g N_BLN<5>_XI0/XI8/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM0 N_XI0/XI8/XI10/NET34_XI0/XI8/XI10/MM0_d
+ N_WL<12>_XI0/XI8/XI10/MM0_g N_BL<5>_XI0/XI8/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM1 N_XI0/XI8/XI10/NET33_XI0/XI8/XI10/MM1_d
+ N_XI0/XI8/XI10/NET34_XI0/XI8/XI10/MM1_g N_VSS_XI0/XI8/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM9 N_XI0/XI8/XI10/NET36_XI0/XI8/XI10/MM9_d
+ N_WL<13>_XI0/XI8/XI10/MM9_g N_BL<5>_XI0/XI8/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM6 N_XI0/XI8/XI10/NET35_XI0/XI8/XI10/MM6_d
+ N_XI0/XI8/XI10/NET36_XI0/XI8/XI10/MM6_g N_VSS_XI0/XI8/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM7 N_XI0/XI8/XI10/NET36_XI0/XI8/XI10/MM7_d
+ N_XI0/XI8/XI10/NET35_XI0/XI8/XI10/MM7_g N_VSS_XI0/XI8/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM8 N_XI0/XI8/XI10/NET35_XI0/XI8/XI10/MM8_d
+ N_WL<13>_XI0/XI8/XI10/MM8_g N_BLN<5>_XI0/XI8/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI10/MM5 N_XI0/XI8/XI10/NET34_XI0/XI8/XI10/MM5_d
+ N_XI0/XI8/XI10/NET33_XI0/XI8/XI10/MM5_g N_VDD_XI0/XI8/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI10/MM4 N_XI0/XI8/XI10/NET33_XI0/XI8/XI10/MM4_d
+ N_XI0/XI8/XI10/NET34_XI0/XI8/XI10/MM4_g N_VDD_XI0/XI8/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI10/MM10 N_XI0/XI8/XI10/NET35_XI0/XI8/XI10/MM10_d
+ N_XI0/XI8/XI10/NET36_XI0/XI8/XI10/MM10_g N_VDD_XI0/XI8/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI10/MM11 N_XI0/XI8/XI10/NET36_XI0/XI8/XI10/MM11_d
+ N_XI0/XI8/XI10/NET35_XI0/XI8/XI10/MM11_g N_VDD_XI0/XI8/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI11/MM2 N_XI0/XI8/XI11/NET34_XI0/XI8/XI11/MM2_d
+ N_XI0/XI8/XI11/NET33_XI0/XI8/XI11/MM2_g N_VSS_XI0/XI8/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM3 N_XI0/XI8/XI11/NET33_XI0/XI8/XI11/MM3_d
+ N_WL<12>_XI0/XI8/XI11/MM3_g N_BLN<4>_XI0/XI8/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM0 N_XI0/XI8/XI11/NET34_XI0/XI8/XI11/MM0_d
+ N_WL<12>_XI0/XI8/XI11/MM0_g N_BL<4>_XI0/XI8/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM1 N_XI0/XI8/XI11/NET33_XI0/XI8/XI11/MM1_d
+ N_XI0/XI8/XI11/NET34_XI0/XI8/XI11/MM1_g N_VSS_XI0/XI8/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM9 N_XI0/XI8/XI11/NET36_XI0/XI8/XI11/MM9_d
+ N_WL<13>_XI0/XI8/XI11/MM9_g N_BL<4>_XI0/XI8/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM6 N_XI0/XI8/XI11/NET35_XI0/XI8/XI11/MM6_d
+ N_XI0/XI8/XI11/NET36_XI0/XI8/XI11/MM6_g N_VSS_XI0/XI8/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM7 N_XI0/XI8/XI11/NET36_XI0/XI8/XI11/MM7_d
+ N_XI0/XI8/XI11/NET35_XI0/XI8/XI11/MM7_g N_VSS_XI0/XI8/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM8 N_XI0/XI8/XI11/NET35_XI0/XI8/XI11/MM8_d
+ N_WL<13>_XI0/XI8/XI11/MM8_g N_BLN<4>_XI0/XI8/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI11/MM5 N_XI0/XI8/XI11/NET34_XI0/XI8/XI11/MM5_d
+ N_XI0/XI8/XI11/NET33_XI0/XI8/XI11/MM5_g N_VDD_XI0/XI8/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI11/MM4 N_XI0/XI8/XI11/NET33_XI0/XI8/XI11/MM4_d
+ N_XI0/XI8/XI11/NET34_XI0/XI8/XI11/MM4_g N_VDD_XI0/XI8/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI11/MM10 N_XI0/XI8/XI11/NET35_XI0/XI8/XI11/MM10_d
+ N_XI0/XI8/XI11/NET36_XI0/XI8/XI11/MM10_g N_VDD_XI0/XI8/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI11/MM11 N_XI0/XI8/XI11/NET36_XI0/XI8/XI11/MM11_d
+ N_XI0/XI8/XI11/NET35_XI0/XI8/XI11/MM11_g N_VDD_XI0/XI8/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI12/MM2 N_XI0/XI8/XI12/NET34_XI0/XI8/XI12/MM2_d
+ N_XI0/XI8/XI12/NET33_XI0/XI8/XI12/MM2_g N_VSS_XI0/XI8/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM3 N_XI0/XI8/XI12/NET33_XI0/XI8/XI12/MM3_d
+ N_WL<12>_XI0/XI8/XI12/MM3_g N_BLN<3>_XI0/XI8/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM0 N_XI0/XI8/XI12/NET34_XI0/XI8/XI12/MM0_d
+ N_WL<12>_XI0/XI8/XI12/MM0_g N_BL<3>_XI0/XI8/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM1 N_XI0/XI8/XI12/NET33_XI0/XI8/XI12/MM1_d
+ N_XI0/XI8/XI12/NET34_XI0/XI8/XI12/MM1_g N_VSS_XI0/XI8/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM9 N_XI0/XI8/XI12/NET36_XI0/XI8/XI12/MM9_d
+ N_WL<13>_XI0/XI8/XI12/MM9_g N_BL<3>_XI0/XI8/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM6 N_XI0/XI8/XI12/NET35_XI0/XI8/XI12/MM6_d
+ N_XI0/XI8/XI12/NET36_XI0/XI8/XI12/MM6_g N_VSS_XI0/XI8/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM7 N_XI0/XI8/XI12/NET36_XI0/XI8/XI12/MM7_d
+ N_XI0/XI8/XI12/NET35_XI0/XI8/XI12/MM7_g N_VSS_XI0/XI8/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM8 N_XI0/XI8/XI12/NET35_XI0/XI8/XI12/MM8_d
+ N_WL<13>_XI0/XI8/XI12/MM8_g N_BLN<3>_XI0/XI8/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI12/MM5 N_XI0/XI8/XI12/NET34_XI0/XI8/XI12/MM5_d
+ N_XI0/XI8/XI12/NET33_XI0/XI8/XI12/MM5_g N_VDD_XI0/XI8/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI12/MM4 N_XI0/XI8/XI12/NET33_XI0/XI8/XI12/MM4_d
+ N_XI0/XI8/XI12/NET34_XI0/XI8/XI12/MM4_g N_VDD_XI0/XI8/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI12/MM10 N_XI0/XI8/XI12/NET35_XI0/XI8/XI12/MM10_d
+ N_XI0/XI8/XI12/NET36_XI0/XI8/XI12/MM10_g N_VDD_XI0/XI8/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI12/MM11 N_XI0/XI8/XI12/NET36_XI0/XI8/XI12/MM11_d
+ N_XI0/XI8/XI12/NET35_XI0/XI8/XI12/MM11_g N_VDD_XI0/XI8/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI13/MM2 N_XI0/XI8/XI13/NET34_XI0/XI8/XI13/MM2_d
+ N_XI0/XI8/XI13/NET33_XI0/XI8/XI13/MM2_g N_VSS_XI0/XI8/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM3 N_XI0/XI8/XI13/NET33_XI0/XI8/XI13/MM3_d
+ N_WL<12>_XI0/XI8/XI13/MM3_g N_BLN<2>_XI0/XI8/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM0 N_XI0/XI8/XI13/NET34_XI0/XI8/XI13/MM0_d
+ N_WL<12>_XI0/XI8/XI13/MM0_g N_BL<2>_XI0/XI8/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM1 N_XI0/XI8/XI13/NET33_XI0/XI8/XI13/MM1_d
+ N_XI0/XI8/XI13/NET34_XI0/XI8/XI13/MM1_g N_VSS_XI0/XI8/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM9 N_XI0/XI8/XI13/NET36_XI0/XI8/XI13/MM9_d
+ N_WL<13>_XI0/XI8/XI13/MM9_g N_BL<2>_XI0/XI8/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM6 N_XI0/XI8/XI13/NET35_XI0/XI8/XI13/MM6_d
+ N_XI0/XI8/XI13/NET36_XI0/XI8/XI13/MM6_g N_VSS_XI0/XI8/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM7 N_XI0/XI8/XI13/NET36_XI0/XI8/XI13/MM7_d
+ N_XI0/XI8/XI13/NET35_XI0/XI8/XI13/MM7_g N_VSS_XI0/XI8/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM8 N_XI0/XI8/XI13/NET35_XI0/XI8/XI13/MM8_d
+ N_WL<13>_XI0/XI8/XI13/MM8_g N_BLN<2>_XI0/XI8/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI13/MM5 N_XI0/XI8/XI13/NET34_XI0/XI8/XI13/MM5_d
+ N_XI0/XI8/XI13/NET33_XI0/XI8/XI13/MM5_g N_VDD_XI0/XI8/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI13/MM4 N_XI0/XI8/XI13/NET33_XI0/XI8/XI13/MM4_d
+ N_XI0/XI8/XI13/NET34_XI0/XI8/XI13/MM4_g N_VDD_XI0/XI8/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI13/MM10 N_XI0/XI8/XI13/NET35_XI0/XI8/XI13/MM10_d
+ N_XI0/XI8/XI13/NET36_XI0/XI8/XI13/MM10_g N_VDD_XI0/XI8/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI13/MM11 N_XI0/XI8/XI13/NET36_XI0/XI8/XI13/MM11_d
+ N_XI0/XI8/XI13/NET35_XI0/XI8/XI13/MM11_g N_VDD_XI0/XI8/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI14/MM2 N_XI0/XI8/XI14/NET34_XI0/XI8/XI14/MM2_d
+ N_XI0/XI8/XI14/NET33_XI0/XI8/XI14/MM2_g N_VSS_XI0/XI8/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM3 N_XI0/XI8/XI14/NET33_XI0/XI8/XI14/MM3_d
+ N_WL<12>_XI0/XI8/XI14/MM3_g N_BLN<1>_XI0/XI8/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM0 N_XI0/XI8/XI14/NET34_XI0/XI8/XI14/MM0_d
+ N_WL<12>_XI0/XI8/XI14/MM0_g N_BL<1>_XI0/XI8/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM1 N_XI0/XI8/XI14/NET33_XI0/XI8/XI14/MM1_d
+ N_XI0/XI8/XI14/NET34_XI0/XI8/XI14/MM1_g N_VSS_XI0/XI8/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM9 N_XI0/XI8/XI14/NET36_XI0/XI8/XI14/MM9_d
+ N_WL<13>_XI0/XI8/XI14/MM9_g N_BL<1>_XI0/XI8/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM6 N_XI0/XI8/XI14/NET35_XI0/XI8/XI14/MM6_d
+ N_XI0/XI8/XI14/NET36_XI0/XI8/XI14/MM6_g N_VSS_XI0/XI8/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM7 N_XI0/XI8/XI14/NET36_XI0/XI8/XI14/MM7_d
+ N_XI0/XI8/XI14/NET35_XI0/XI8/XI14/MM7_g N_VSS_XI0/XI8/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM8 N_XI0/XI8/XI14/NET35_XI0/XI8/XI14/MM8_d
+ N_WL<13>_XI0/XI8/XI14/MM8_g N_BLN<1>_XI0/XI8/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI14/MM5 N_XI0/XI8/XI14/NET34_XI0/XI8/XI14/MM5_d
+ N_XI0/XI8/XI14/NET33_XI0/XI8/XI14/MM5_g N_VDD_XI0/XI8/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI14/MM4 N_XI0/XI8/XI14/NET33_XI0/XI8/XI14/MM4_d
+ N_XI0/XI8/XI14/NET34_XI0/XI8/XI14/MM4_g N_VDD_XI0/XI8/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI14/MM10 N_XI0/XI8/XI14/NET35_XI0/XI8/XI14/MM10_d
+ N_XI0/XI8/XI14/NET36_XI0/XI8/XI14/MM10_g N_VDD_XI0/XI8/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI14/MM11 N_XI0/XI8/XI14/NET36_XI0/XI8/XI14/MM11_d
+ N_XI0/XI8/XI14/NET35_XI0/XI8/XI14/MM11_g N_VDD_XI0/XI8/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI15/MM2 N_XI0/XI8/XI15/NET34_XI0/XI8/XI15/MM2_d
+ N_XI0/XI8/XI15/NET33_XI0/XI8/XI15/MM2_g N_VSS_XI0/XI8/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM3 N_XI0/XI8/XI15/NET33_XI0/XI8/XI15/MM3_d
+ N_WL<12>_XI0/XI8/XI15/MM3_g N_BLN<0>_XI0/XI8/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM0 N_XI0/XI8/XI15/NET34_XI0/XI8/XI15/MM0_d
+ N_WL<12>_XI0/XI8/XI15/MM0_g N_BL<0>_XI0/XI8/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM1 N_XI0/XI8/XI15/NET33_XI0/XI8/XI15/MM1_d
+ N_XI0/XI8/XI15/NET34_XI0/XI8/XI15/MM1_g N_VSS_XI0/XI8/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM9 N_XI0/XI8/XI15/NET36_XI0/XI8/XI15/MM9_d
+ N_WL<13>_XI0/XI8/XI15/MM9_g N_BL<0>_XI0/XI8/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM6 N_XI0/XI8/XI15/NET35_XI0/XI8/XI15/MM6_d
+ N_XI0/XI8/XI15/NET36_XI0/XI8/XI15/MM6_g N_VSS_XI0/XI8/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM7 N_XI0/XI8/XI15/NET36_XI0/XI8/XI15/MM7_d
+ N_XI0/XI8/XI15/NET35_XI0/XI8/XI15/MM7_g N_VSS_XI0/XI8/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM8 N_XI0/XI8/XI15/NET35_XI0/XI8/XI15/MM8_d
+ N_WL<13>_XI0/XI8/XI15/MM8_g N_BLN<0>_XI0/XI8/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/XI15/MM5 N_XI0/XI8/XI15/NET34_XI0/XI8/XI15/MM5_d
+ N_XI0/XI8/XI15/NET33_XI0/XI8/XI15/MM5_g N_VDD_XI0/XI8/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI15/MM4 N_XI0/XI8/XI15/NET33_XI0/XI8/XI15/MM4_d
+ N_XI0/XI8/XI15/NET34_XI0/XI8/XI15/MM4_g N_VDD_XI0/XI8/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI15/MM10 N_XI0/XI8/XI15/NET35_XI0/XI8/XI15/MM10_d
+ N_XI0/XI8/XI15/NET36_XI0/XI8/XI15/MM10_g N_VDD_XI0/XI8/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/XI15/MM11 N_XI0/XI8/XI15/NET36_XI0/XI8/XI15/MM11_d
+ N_XI0/XI8/XI15/NET35_XI0/XI8/XI15/MM11_g N_VDD_XI0/XI8/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI0/MM2 N_XI0/XI9/XI0/NET34_XI0/XI9/XI0/MM2_d
+ N_XI0/XI9/XI0/NET33_XI0/XI9/XI0/MM2_g N_VSS_XI0/XI9/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM3 N_XI0/XI9/XI0/NET33_XI0/XI9/XI0/MM3_d
+ N_WL<14>_XI0/XI9/XI0/MM3_g N_BLN<15>_XI0/XI9/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM0 N_XI0/XI9/XI0/NET34_XI0/XI9/XI0/MM0_d
+ N_WL<14>_XI0/XI9/XI0/MM0_g N_BL<15>_XI0/XI9/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM1 N_XI0/XI9/XI0/NET33_XI0/XI9/XI0/MM1_d
+ N_XI0/XI9/XI0/NET34_XI0/XI9/XI0/MM1_g N_VSS_XI0/XI9/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM9 N_XI0/XI9/XI0/NET36_XI0/XI9/XI0/MM9_d
+ N_WL<15>_XI0/XI9/XI0/MM9_g N_BL<15>_XI0/XI9/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM6 N_XI0/XI9/XI0/NET35_XI0/XI9/XI0/MM6_d
+ N_XI0/XI9/XI0/NET36_XI0/XI9/XI0/MM6_g N_VSS_XI0/XI9/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM7 N_XI0/XI9/XI0/NET36_XI0/XI9/XI0/MM7_d
+ N_XI0/XI9/XI0/NET35_XI0/XI9/XI0/MM7_g N_VSS_XI0/XI9/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM8 N_XI0/XI9/XI0/NET35_XI0/XI9/XI0/MM8_d
+ N_WL<15>_XI0/XI9/XI0/MM8_g N_BLN<15>_XI0/XI9/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI0/MM5 N_XI0/XI9/XI0/NET34_XI0/XI9/XI0/MM5_d
+ N_XI0/XI9/XI0/NET33_XI0/XI9/XI0/MM5_g N_VDD_XI0/XI9/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI0/MM4 N_XI0/XI9/XI0/NET33_XI0/XI9/XI0/MM4_d
+ N_XI0/XI9/XI0/NET34_XI0/XI9/XI0/MM4_g N_VDD_XI0/XI9/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI0/MM10 N_XI0/XI9/XI0/NET35_XI0/XI9/XI0/MM10_d
+ N_XI0/XI9/XI0/NET36_XI0/XI9/XI0/MM10_g N_VDD_XI0/XI9/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI0/MM11 N_XI0/XI9/XI0/NET36_XI0/XI9/XI0/MM11_d
+ N_XI0/XI9/XI0/NET35_XI0/XI9/XI0/MM11_g N_VDD_XI0/XI9/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI1/MM2 N_XI0/XI9/XI1/NET34_XI0/XI9/XI1/MM2_d
+ N_XI0/XI9/XI1/NET33_XI0/XI9/XI1/MM2_g N_VSS_XI0/XI9/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM3 N_XI0/XI9/XI1/NET33_XI0/XI9/XI1/MM3_d
+ N_WL<14>_XI0/XI9/XI1/MM3_g N_BLN<14>_XI0/XI9/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM0 N_XI0/XI9/XI1/NET34_XI0/XI9/XI1/MM0_d
+ N_WL<14>_XI0/XI9/XI1/MM0_g N_BL<14>_XI0/XI9/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM1 N_XI0/XI9/XI1/NET33_XI0/XI9/XI1/MM1_d
+ N_XI0/XI9/XI1/NET34_XI0/XI9/XI1/MM1_g N_VSS_XI0/XI9/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM9 N_XI0/XI9/XI1/NET36_XI0/XI9/XI1/MM9_d
+ N_WL<15>_XI0/XI9/XI1/MM9_g N_BL<14>_XI0/XI9/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM6 N_XI0/XI9/XI1/NET35_XI0/XI9/XI1/MM6_d
+ N_XI0/XI9/XI1/NET36_XI0/XI9/XI1/MM6_g N_VSS_XI0/XI9/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM7 N_XI0/XI9/XI1/NET36_XI0/XI9/XI1/MM7_d
+ N_XI0/XI9/XI1/NET35_XI0/XI9/XI1/MM7_g N_VSS_XI0/XI9/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM8 N_XI0/XI9/XI1/NET35_XI0/XI9/XI1/MM8_d
+ N_WL<15>_XI0/XI9/XI1/MM8_g N_BLN<14>_XI0/XI9/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI1/MM5 N_XI0/XI9/XI1/NET34_XI0/XI9/XI1/MM5_d
+ N_XI0/XI9/XI1/NET33_XI0/XI9/XI1/MM5_g N_VDD_XI0/XI9/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI1/MM4 N_XI0/XI9/XI1/NET33_XI0/XI9/XI1/MM4_d
+ N_XI0/XI9/XI1/NET34_XI0/XI9/XI1/MM4_g N_VDD_XI0/XI9/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI1/MM10 N_XI0/XI9/XI1/NET35_XI0/XI9/XI1/MM10_d
+ N_XI0/XI9/XI1/NET36_XI0/XI9/XI1/MM10_g N_VDD_XI0/XI9/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI1/MM11 N_XI0/XI9/XI1/NET36_XI0/XI9/XI1/MM11_d
+ N_XI0/XI9/XI1/NET35_XI0/XI9/XI1/MM11_g N_VDD_XI0/XI9/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI2/MM2 N_XI0/XI9/XI2/NET34_XI0/XI9/XI2/MM2_d
+ N_XI0/XI9/XI2/NET33_XI0/XI9/XI2/MM2_g N_VSS_XI0/XI9/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM3 N_XI0/XI9/XI2/NET33_XI0/XI9/XI2/MM3_d
+ N_WL<14>_XI0/XI9/XI2/MM3_g N_BLN<13>_XI0/XI9/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM0 N_XI0/XI9/XI2/NET34_XI0/XI9/XI2/MM0_d
+ N_WL<14>_XI0/XI9/XI2/MM0_g N_BL<13>_XI0/XI9/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM1 N_XI0/XI9/XI2/NET33_XI0/XI9/XI2/MM1_d
+ N_XI0/XI9/XI2/NET34_XI0/XI9/XI2/MM1_g N_VSS_XI0/XI9/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM9 N_XI0/XI9/XI2/NET36_XI0/XI9/XI2/MM9_d
+ N_WL<15>_XI0/XI9/XI2/MM9_g N_BL<13>_XI0/XI9/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM6 N_XI0/XI9/XI2/NET35_XI0/XI9/XI2/MM6_d
+ N_XI0/XI9/XI2/NET36_XI0/XI9/XI2/MM6_g N_VSS_XI0/XI9/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM7 N_XI0/XI9/XI2/NET36_XI0/XI9/XI2/MM7_d
+ N_XI0/XI9/XI2/NET35_XI0/XI9/XI2/MM7_g N_VSS_XI0/XI9/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM8 N_XI0/XI9/XI2/NET35_XI0/XI9/XI2/MM8_d
+ N_WL<15>_XI0/XI9/XI2/MM8_g N_BLN<13>_XI0/XI9/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI2/MM5 N_XI0/XI9/XI2/NET34_XI0/XI9/XI2/MM5_d
+ N_XI0/XI9/XI2/NET33_XI0/XI9/XI2/MM5_g N_VDD_XI0/XI9/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI2/MM4 N_XI0/XI9/XI2/NET33_XI0/XI9/XI2/MM4_d
+ N_XI0/XI9/XI2/NET34_XI0/XI9/XI2/MM4_g N_VDD_XI0/XI9/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI2/MM10 N_XI0/XI9/XI2/NET35_XI0/XI9/XI2/MM10_d
+ N_XI0/XI9/XI2/NET36_XI0/XI9/XI2/MM10_g N_VDD_XI0/XI9/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI2/MM11 N_XI0/XI9/XI2/NET36_XI0/XI9/XI2/MM11_d
+ N_XI0/XI9/XI2/NET35_XI0/XI9/XI2/MM11_g N_VDD_XI0/XI9/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI3/MM2 N_XI0/XI9/XI3/NET34_XI0/XI9/XI3/MM2_d
+ N_XI0/XI9/XI3/NET33_XI0/XI9/XI3/MM2_g N_VSS_XI0/XI9/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM3 N_XI0/XI9/XI3/NET33_XI0/XI9/XI3/MM3_d
+ N_WL<14>_XI0/XI9/XI3/MM3_g N_BLN<12>_XI0/XI9/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM0 N_XI0/XI9/XI3/NET34_XI0/XI9/XI3/MM0_d
+ N_WL<14>_XI0/XI9/XI3/MM0_g N_BL<12>_XI0/XI9/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM1 N_XI0/XI9/XI3/NET33_XI0/XI9/XI3/MM1_d
+ N_XI0/XI9/XI3/NET34_XI0/XI9/XI3/MM1_g N_VSS_XI0/XI9/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM9 N_XI0/XI9/XI3/NET36_XI0/XI9/XI3/MM9_d
+ N_WL<15>_XI0/XI9/XI3/MM9_g N_BL<12>_XI0/XI9/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM6 N_XI0/XI9/XI3/NET35_XI0/XI9/XI3/MM6_d
+ N_XI0/XI9/XI3/NET36_XI0/XI9/XI3/MM6_g N_VSS_XI0/XI9/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM7 N_XI0/XI9/XI3/NET36_XI0/XI9/XI3/MM7_d
+ N_XI0/XI9/XI3/NET35_XI0/XI9/XI3/MM7_g N_VSS_XI0/XI9/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM8 N_XI0/XI9/XI3/NET35_XI0/XI9/XI3/MM8_d
+ N_WL<15>_XI0/XI9/XI3/MM8_g N_BLN<12>_XI0/XI9/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI3/MM5 N_XI0/XI9/XI3/NET34_XI0/XI9/XI3/MM5_d
+ N_XI0/XI9/XI3/NET33_XI0/XI9/XI3/MM5_g N_VDD_XI0/XI9/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI3/MM4 N_XI0/XI9/XI3/NET33_XI0/XI9/XI3/MM4_d
+ N_XI0/XI9/XI3/NET34_XI0/XI9/XI3/MM4_g N_VDD_XI0/XI9/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI3/MM10 N_XI0/XI9/XI3/NET35_XI0/XI9/XI3/MM10_d
+ N_XI0/XI9/XI3/NET36_XI0/XI9/XI3/MM10_g N_VDD_XI0/XI9/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI3/MM11 N_XI0/XI9/XI3/NET36_XI0/XI9/XI3/MM11_d
+ N_XI0/XI9/XI3/NET35_XI0/XI9/XI3/MM11_g N_VDD_XI0/XI9/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI4/MM2 N_XI0/XI9/XI4/NET34_XI0/XI9/XI4/MM2_d
+ N_XI0/XI9/XI4/NET33_XI0/XI9/XI4/MM2_g N_VSS_XI0/XI9/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM3 N_XI0/XI9/XI4/NET33_XI0/XI9/XI4/MM3_d
+ N_WL<14>_XI0/XI9/XI4/MM3_g N_BLN<11>_XI0/XI9/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM0 N_XI0/XI9/XI4/NET34_XI0/XI9/XI4/MM0_d
+ N_WL<14>_XI0/XI9/XI4/MM0_g N_BL<11>_XI0/XI9/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM1 N_XI0/XI9/XI4/NET33_XI0/XI9/XI4/MM1_d
+ N_XI0/XI9/XI4/NET34_XI0/XI9/XI4/MM1_g N_VSS_XI0/XI9/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM9 N_XI0/XI9/XI4/NET36_XI0/XI9/XI4/MM9_d
+ N_WL<15>_XI0/XI9/XI4/MM9_g N_BL<11>_XI0/XI9/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM6 N_XI0/XI9/XI4/NET35_XI0/XI9/XI4/MM6_d
+ N_XI0/XI9/XI4/NET36_XI0/XI9/XI4/MM6_g N_VSS_XI0/XI9/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM7 N_XI0/XI9/XI4/NET36_XI0/XI9/XI4/MM7_d
+ N_XI0/XI9/XI4/NET35_XI0/XI9/XI4/MM7_g N_VSS_XI0/XI9/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM8 N_XI0/XI9/XI4/NET35_XI0/XI9/XI4/MM8_d
+ N_WL<15>_XI0/XI9/XI4/MM8_g N_BLN<11>_XI0/XI9/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI4/MM5 N_XI0/XI9/XI4/NET34_XI0/XI9/XI4/MM5_d
+ N_XI0/XI9/XI4/NET33_XI0/XI9/XI4/MM5_g N_VDD_XI0/XI9/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI4/MM4 N_XI0/XI9/XI4/NET33_XI0/XI9/XI4/MM4_d
+ N_XI0/XI9/XI4/NET34_XI0/XI9/XI4/MM4_g N_VDD_XI0/XI9/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI4/MM10 N_XI0/XI9/XI4/NET35_XI0/XI9/XI4/MM10_d
+ N_XI0/XI9/XI4/NET36_XI0/XI9/XI4/MM10_g N_VDD_XI0/XI9/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI4/MM11 N_XI0/XI9/XI4/NET36_XI0/XI9/XI4/MM11_d
+ N_XI0/XI9/XI4/NET35_XI0/XI9/XI4/MM11_g N_VDD_XI0/XI9/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI5/MM2 N_XI0/XI9/XI5/NET34_XI0/XI9/XI5/MM2_d
+ N_XI0/XI9/XI5/NET33_XI0/XI9/XI5/MM2_g N_VSS_XI0/XI9/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM3 N_XI0/XI9/XI5/NET33_XI0/XI9/XI5/MM3_d
+ N_WL<14>_XI0/XI9/XI5/MM3_g N_BLN<10>_XI0/XI9/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM0 N_XI0/XI9/XI5/NET34_XI0/XI9/XI5/MM0_d
+ N_WL<14>_XI0/XI9/XI5/MM0_g N_BL<10>_XI0/XI9/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM1 N_XI0/XI9/XI5/NET33_XI0/XI9/XI5/MM1_d
+ N_XI0/XI9/XI5/NET34_XI0/XI9/XI5/MM1_g N_VSS_XI0/XI9/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM9 N_XI0/XI9/XI5/NET36_XI0/XI9/XI5/MM9_d
+ N_WL<15>_XI0/XI9/XI5/MM9_g N_BL<10>_XI0/XI9/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM6 N_XI0/XI9/XI5/NET35_XI0/XI9/XI5/MM6_d
+ N_XI0/XI9/XI5/NET36_XI0/XI9/XI5/MM6_g N_VSS_XI0/XI9/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM7 N_XI0/XI9/XI5/NET36_XI0/XI9/XI5/MM7_d
+ N_XI0/XI9/XI5/NET35_XI0/XI9/XI5/MM7_g N_VSS_XI0/XI9/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM8 N_XI0/XI9/XI5/NET35_XI0/XI9/XI5/MM8_d
+ N_WL<15>_XI0/XI9/XI5/MM8_g N_BLN<10>_XI0/XI9/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI5/MM5 N_XI0/XI9/XI5/NET34_XI0/XI9/XI5/MM5_d
+ N_XI0/XI9/XI5/NET33_XI0/XI9/XI5/MM5_g N_VDD_XI0/XI9/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI5/MM4 N_XI0/XI9/XI5/NET33_XI0/XI9/XI5/MM4_d
+ N_XI0/XI9/XI5/NET34_XI0/XI9/XI5/MM4_g N_VDD_XI0/XI9/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI5/MM10 N_XI0/XI9/XI5/NET35_XI0/XI9/XI5/MM10_d
+ N_XI0/XI9/XI5/NET36_XI0/XI9/XI5/MM10_g N_VDD_XI0/XI9/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI5/MM11 N_XI0/XI9/XI5/NET36_XI0/XI9/XI5/MM11_d
+ N_XI0/XI9/XI5/NET35_XI0/XI9/XI5/MM11_g N_VDD_XI0/XI9/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI6/MM2 N_XI0/XI9/XI6/NET34_XI0/XI9/XI6/MM2_d
+ N_XI0/XI9/XI6/NET33_XI0/XI9/XI6/MM2_g N_VSS_XI0/XI9/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM3 N_XI0/XI9/XI6/NET33_XI0/XI9/XI6/MM3_d
+ N_WL<14>_XI0/XI9/XI6/MM3_g N_BLN<9>_XI0/XI9/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM0 N_XI0/XI9/XI6/NET34_XI0/XI9/XI6/MM0_d
+ N_WL<14>_XI0/XI9/XI6/MM0_g N_BL<9>_XI0/XI9/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM1 N_XI0/XI9/XI6/NET33_XI0/XI9/XI6/MM1_d
+ N_XI0/XI9/XI6/NET34_XI0/XI9/XI6/MM1_g N_VSS_XI0/XI9/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM9 N_XI0/XI9/XI6/NET36_XI0/XI9/XI6/MM9_d
+ N_WL<15>_XI0/XI9/XI6/MM9_g N_BL<9>_XI0/XI9/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM6 N_XI0/XI9/XI6/NET35_XI0/XI9/XI6/MM6_d
+ N_XI0/XI9/XI6/NET36_XI0/XI9/XI6/MM6_g N_VSS_XI0/XI9/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM7 N_XI0/XI9/XI6/NET36_XI0/XI9/XI6/MM7_d
+ N_XI0/XI9/XI6/NET35_XI0/XI9/XI6/MM7_g N_VSS_XI0/XI9/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM8 N_XI0/XI9/XI6/NET35_XI0/XI9/XI6/MM8_d
+ N_WL<15>_XI0/XI9/XI6/MM8_g N_BLN<9>_XI0/XI9/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI6/MM5 N_XI0/XI9/XI6/NET34_XI0/XI9/XI6/MM5_d
+ N_XI0/XI9/XI6/NET33_XI0/XI9/XI6/MM5_g N_VDD_XI0/XI9/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI6/MM4 N_XI0/XI9/XI6/NET33_XI0/XI9/XI6/MM4_d
+ N_XI0/XI9/XI6/NET34_XI0/XI9/XI6/MM4_g N_VDD_XI0/XI9/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI6/MM10 N_XI0/XI9/XI6/NET35_XI0/XI9/XI6/MM10_d
+ N_XI0/XI9/XI6/NET36_XI0/XI9/XI6/MM10_g N_VDD_XI0/XI9/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI6/MM11 N_XI0/XI9/XI6/NET36_XI0/XI9/XI6/MM11_d
+ N_XI0/XI9/XI6/NET35_XI0/XI9/XI6/MM11_g N_VDD_XI0/XI9/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI7/MM2 N_XI0/XI9/XI7/NET34_XI0/XI9/XI7/MM2_d
+ N_XI0/XI9/XI7/NET33_XI0/XI9/XI7/MM2_g N_VSS_XI0/XI9/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM3 N_XI0/XI9/XI7/NET33_XI0/XI9/XI7/MM3_d
+ N_WL<14>_XI0/XI9/XI7/MM3_g N_BLN<8>_XI0/XI9/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM0 N_XI0/XI9/XI7/NET34_XI0/XI9/XI7/MM0_d
+ N_WL<14>_XI0/XI9/XI7/MM0_g N_BL<8>_XI0/XI9/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM1 N_XI0/XI9/XI7/NET33_XI0/XI9/XI7/MM1_d
+ N_XI0/XI9/XI7/NET34_XI0/XI9/XI7/MM1_g N_VSS_XI0/XI9/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM9 N_XI0/XI9/XI7/NET36_XI0/XI9/XI7/MM9_d
+ N_WL<15>_XI0/XI9/XI7/MM9_g N_BL<8>_XI0/XI9/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM6 N_XI0/XI9/XI7/NET35_XI0/XI9/XI7/MM6_d
+ N_XI0/XI9/XI7/NET36_XI0/XI9/XI7/MM6_g N_VSS_XI0/XI9/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM7 N_XI0/XI9/XI7/NET36_XI0/XI9/XI7/MM7_d
+ N_XI0/XI9/XI7/NET35_XI0/XI9/XI7/MM7_g N_VSS_XI0/XI9/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM8 N_XI0/XI9/XI7/NET35_XI0/XI9/XI7/MM8_d
+ N_WL<15>_XI0/XI9/XI7/MM8_g N_BLN<8>_XI0/XI9/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI7/MM5 N_XI0/XI9/XI7/NET34_XI0/XI9/XI7/MM5_d
+ N_XI0/XI9/XI7/NET33_XI0/XI9/XI7/MM5_g N_VDD_XI0/XI9/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI7/MM4 N_XI0/XI9/XI7/NET33_XI0/XI9/XI7/MM4_d
+ N_XI0/XI9/XI7/NET34_XI0/XI9/XI7/MM4_g N_VDD_XI0/XI9/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI7/MM10 N_XI0/XI9/XI7/NET35_XI0/XI9/XI7/MM10_d
+ N_XI0/XI9/XI7/NET36_XI0/XI9/XI7/MM10_g N_VDD_XI0/XI9/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI7/MM11 N_XI0/XI9/XI7/NET36_XI0/XI9/XI7/MM11_d
+ N_XI0/XI9/XI7/NET35_XI0/XI9/XI7/MM11_g N_VDD_XI0/XI9/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI8/MM2 N_XI0/XI9/XI8/NET34_XI0/XI9/XI8/MM2_d
+ N_XI0/XI9/XI8/NET33_XI0/XI9/XI8/MM2_g N_VSS_XI0/XI9/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM3 N_XI0/XI9/XI8/NET33_XI0/XI9/XI8/MM3_d
+ N_WL<14>_XI0/XI9/XI8/MM3_g N_BLN<7>_XI0/XI9/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM0 N_XI0/XI9/XI8/NET34_XI0/XI9/XI8/MM0_d
+ N_WL<14>_XI0/XI9/XI8/MM0_g N_BL<7>_XI0/XI9/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM1 N_XI0/XI9/XI8/NET33_XI0/XI9/XI8/MM1_d
+ N_XI0/XI9/XI8/NET34_XI0/XI9/XI8/MM1_g N_VSS_XI0/XI9/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM9 N_XI0/XI9/XI8/NET36_XI0/XI9/XI8/MM9_d
+ N_WL<15>_XI0/XI9/XI8/MM9_g N_BL<7>_XI0/XI9/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM6 N_XI0/XI9/XI8/NET35_XI0/XI9/XI8/MM6_d
+ N_XI0/XI9/XI8/NET36_XI0/XI9/XI8/MM6_g N_VSS_XI0/XI9/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM7 N_XI0/XI9/XI8/NET36_XI0/XI9/XI8/MM7_d
+ N_XI0/XI9/XI8/NET35_XI0/XI9/XI8/MM7_g N_VSS_XI0/XI9/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM8 N_XI0/XI9/XI8/NET35_XI0/XI9/XI8/MM8_d
+ N_WL<15>_XI0/XI9/XI8/MM8_g N_BLN<7>_XI0/XI9/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI8/MM5 N_XI0/XI9/XI8/NET34_XI0/XI9/XI8/MM5_d
+ N_XI0/XI9/XI8/NET33_XI0/XI9/XI8/MM5_g N_VDD_XI0/XI9/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI8/MM4 N_XI0/XI9/XI8/NET33_XI0/XI9/XI8/MM4_d
+ N_XI0/XI9/XI8/NET34_XI0/XI9/XI8/MM4_g N_VDD_XI0/XI9/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI8/MM10 N_XI0/XI9/XI8/NET35_XI0/XI9/XI8/MM10_d
+ N_XI0/XI9/XI8/NET36_XI0/XI9/XI8/MM10_g N_VDD_XI0/XI9/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI8/MM11 N_XI0/XI9/XI8/NET36_XI0/XI9/XI8/MM11_d
+ N_XI0/XI9/XI8/NET35_XI0/XI9/XI8/MM11_g N_VDD_XI0/XI9/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI9/MM2 N_XI0/XI9/XI9/NET34_XI0/XI9/XI9/MM2_d
+ N_XI0/XI9/XI9/NET33_XI0/XI9/XI9/MM2_g N_VSS_XI0/XI9/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM3 N_XI0/XI9/XI9/NET33_XI0/XI9/XI9/MM3_d
+ N_WL<14>_XI0/XI9/XI9/MM3_g N_BLN<6>_XI0/XI9/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM0 N_XI0/XI9/XI9/NET34_XI0/XI9/XI9/MM0_d
+ N_WL<14>_XI0/XI9/XI9/MM0_g N_BL<6>_XI0/XI9/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM1 N_XI0/XI9/XI9/NET33_XI0/XI9/XI9/MM1_d
+ N_XI0/XI9/XI9/NET34_XI0/XI9/XI9/MM1_g N_VSS_XI0/XI9/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM9 N_XI0/XI9/XI9/NET36_XI0/XI9/XI9/MM9_d
+ N_WL<15>_XI0/XI9/XI9/MM9_g N_BL<6>_XI0/XI9/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM6 N_XI0/XI9/XI9/NET35_XI0/XI9/XI9/MM6_d
+ N_XI0/XI9/XI9/NET36_XI0/XI9/XI9/MM6_g N_VSS_XI0/XI9/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM7 N_XI0/XI9/XI9/NET36_XI0/XI9/XI9/MM7_d
+ N_XI0/XI9/XI9/NET35_XI0/XI9/XI9/MM7_g N_VSS_XI0/XI9/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM8 N_XI0/XI9/XI9/NET35_XI0/XI9/XI9/MM8_d
+ N_WL<15>_XI0/XI9/XI9/MM8_g N_BLN<6>_XI0/XI9/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI9/MM5 N_XI0/XI9/XI9/NET34_XI0/XI9/XI9/MM5_d
+ N_XI0/XI9/XI9/NET33_XI0/XI9/XI9/MM5_g N_VDD_XI0/XI9/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI9/MM4 N_XI0/XI9/XI9/NET33_XI0/XI9/XI9/MM4_d
+ N_XI0/XI9/XI9/NET34_XI0/XI9/XI9/MM4_g N_VDD_XI0/XI9/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI9/MM10 N_XI0/XI9/XI9/NET35_XI0/XI9/XI9/MM10_d
+ N_XI0/XI9/XI9/NET36_XI0/XI9/XI9/MM10_g N_VDD_XI0/XI9/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI9/MM11 N_XI0/XI9/XI9/NET36_XI0/XI9/XI9/MM11_d
+ N_XI0/XI9/XI9/NET35_XI0/XI9/XI9/MM11_g N_VDD_XI0/XI9/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI10/MM2 N_XI0/XI9/XI10/NET34_XI0/XI9/XI10/MM2_d
+ N_XI0/XI9/XI10/NET33_XI0/XI9/XI10/MM2_g N_VSS_XI0/XI9/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM3 N_XI0/XI9/XI10/NET33_XI0/XI9/XI10/MM3_d
+ N_WL<14>_XI0/XI9/XI10/MM3_g N_BLN<5>_XI0/XI9/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM0 N_XI0/XI9/XI10/NET34_XI0/XI9/XI10/MM0_d
+ N_WL<14>_XI0/XI9/XI10/MM0_g N_BL<5>_XI0/XI9/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM1 N_XI0/XI9/XI10/NET33_XI0/XI9/XI10/MM1_d
+ N_XI0/XI9/XI10/NET34_XI0/XI9/XI10/MM1_g N_VSS_XI0/XI9/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM9 N_XI0/XI9/XI10/NET36_XI0/XI9/XI10/MM9_d
+ N_WL<15>_XI0/XI9/XI10/MM9_g N_BL<5>_XI0/XI9/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM6 N_XI0/XI9/XI10/NET35_XI0/XI9/XI10/MM6_d
+ N_XI0/XI9/XI10/NET36_XI0/XI9/XI10/MM6_g N_VSS_XI0/XI9/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM7 N_XI0/XI9/XI10/NET36_XI0/XI9/XI10/MM7_d
+ N_XI0/XI9/XI10/NET35_XI0/XI9/XI10/MM7_g N_VSS_XI0/XI9/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM8 N_XI0/XI9/XI10/NET35_XI0/XI9/XI10/MM8_d
+ N_WL<15>_XI0/XI9/XI10/MM8_g N_BLN<5>_XI0/XI9/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI10/MM5 N_XI0/XI9/XI10/NET34_XI0/XI9/XI10/MM5_d
+ N_XI0/XI9/XI10/NET33_XI0/XI9/XI10/MM5_g N_VDD_XI0/XI9/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI10/MM4 N_XI0/XI9/XI10/NET33_XI0/XI9/XI10/MM4_d
+ N_XI0/XI9/XI10/NET34_XI0/XI9/XI10/MM4_g N_VDD_XI0/XI9/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI10/MM10 N_XI0/XI9/XI10/NET35_XI0/XI9/XI10/MM10_d
+ N_XI0/XI9/XI10/NET36_XI0/XI9/XI10/MM10_g N_VDD_XI0/XI9/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI10/MM11 N_XI0/XI9/XI10/NET36_XI0/XI9/XI10/MM11_d
+ N_XI0/XI9/XI10/NET35_XI0/XI9/XI10/MM11_g N_VDD_XI0/XI9/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI11/MM2 N_XI0/XI9/XI11/NET34_XI0/XI9/XI11/MM2_d
+ N_XI0/XI9/XI11/NET33_XI0/XI9/XI11/MM2_g N_VSS_XI0/XI9/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM3 N_XI0/XI9/XI11/NET33_XI0/XI9/XI11/MM3_d
+ N_WL<14>_XI0/XI9/XI11/MM3_g N_BLN<4>_XI0/XI9/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM0 N_XI0/XI9/XI11/NET34_XI0/XI9/XI11/MM0_d
+ N_WL<14>_XI0/XI9/XI11/MM0_g N_BL<4>_XI0/XI9/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM1 N_XI0/XI9/XI11/NET33_XI0/XI9/XI11/MM1_d
+ N_XI0/XI9/XI11/NET34_XI0/XI9/XI11/MM1_g N_VSS_XI0/XI9/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM9 N_XI0/XI9/XI11/NET36_XI0/XI9/XI11/MM9_d
+ N_WL<15>_XI0/XI9/XI11/MM9_g N_BL<4>_XI0/XI9/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM6 N_XI0/XI9/XI11/NET35_XI0/XI9/XI11/MM6_d
+ N_XI0/XI9/XI11/NET36_XI0/XI9/XI11/MM6_g N_VSS_XI0/XI9/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM7 N_XI0/XI9/XI11/NET36_XI0/XI9/XI11/MM7_d
+ N_XI0/XI9/XI11/NET35_XI0/XI9/XI11/MM7_g N_VSS_XI0/XI9/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM8 N_XI0/XI9/XI11/NET35_XI0/XI9/XI11/MM8_d
+ N_WL<15>_XI0/XI9/XI11/MM8_g N_BLN<4>_XI0/XI9/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI11/MM5 N_XI0/XI9/XI11/NET34_XI0/XI9/XI11/MM5_d
+ N_XI0/XI9/XI11/NET33_XI0/XI9/XI11/MM5_g N_VDD_XI0/XI9/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI11/MM4 N_XI0/XI9/XI11/NET33_XI0/XI9/XI11/MM4_d
+ N_XI0/XI9/XI11/NET34_XI0/XI9/XI11/MM4_g N_VDD_XI0/XI9/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI11/MM10 N_XI0/XI9/XI11/NET35_XI0/XI9/XI11/MM10_d
+ N_XI0/XI9/XI11/NET36_XI0/XI9/XI11/MM10_g N_VDD_XI0/XI9/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI11/MM11 N_XI0/XI9/XI11/NET36_XI0/XI9/XI11/MM11_d
+ N_XI0/XI9/XI11/NET35_XI0/XI9/XI11/MM11_g N_VDD_XI0/XI9/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI12/MM2 N_XI0/XI9/XI12/NET34_XI0/XI9/XI12/MM2_d
+ N_XI0/XI9/XI12/NET33_XI0/XI9/XI12/MM2_g N_VSS_XI0/XI9/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM3 N_XI0/XI9/XI12/NET33_XI0/XI9/XI12/MM3_d
+ N_WL<14>_XI0/XI9/XI12/MM3_g N_BLN<3>_XI0/XI9/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM0 N_XI0/XI9/XI12/NET34_XI0/XI9/XI12/MM0_d
+ N_WL<14>_XI0/XI9/XI12/MM0_g N_BL<3>_XI0/XI9/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM1 N_XI0/XI9/XI12/NET33_XI0/XI9/XI12/MM1_d
+ N_XI0/XI9/XI12/NET34_XI0/XI9/XI12/MM1_g N_VSS_XI0/XI9/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM9 N_XI0/XI9/XI12/NET36_XI0/XI9/XI12/MM9_d
+ N_WL<15>_XI0/XI9/XI12/MM9_g N_BL<3>_XI0/XI9/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM6 N_XI0/XI9/XI12/NET35_XI0/XI9/XI12/MM6_d
+ N_XI0/XI9/XI12/NET36_XI0/XI9/XI12/MM6_g N_VSS_XI0/XI9/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM7 N_XI0/XI9/XI12/NET36_XI0/XI9/XI12/MM7_d
+ N_XI0/XI9/XI12/NET35_XI0/XI9/XI12/MM7_g N_VSS_XI0/XI9/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM8 N_XI0/XI9/XI12/NET35_XI0/XI9/XI12/MM8_d
+ N_WL<15>_XI0/XI9/XI12/MM8_g N_BLN<3>_XI0/XI9/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI12/MM5 N_XI0/XI9/XI12/NET34_XI0/XI9/XI12/MM5_d
+ N_XI0/XI9/XI12/NET33_XI0/XI9/XI12/MM5_g N_VDD_XI0/XI9/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI12/MM4 N_XI0/XI9/XI12/NET33_XI0/XI9/XI12/MM4_d
+ N_XI0/XI9/XI12/NET34_XI0/XI9/XI12/MM4_g N_VDD_XI0/XI9/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI12/MM10 N_XI0/XI9/XI12/NET35_XI0/XI9/XI12/MM10_d
+ N_XI0/XI9/XI12/NET36_XI0/XI9/XI12/MM10_g N_VDD_XI0/XI9/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI12/MM11 N_XI0/XI9/XI12/NET36_XI0/XI9/XI12/MM11_d
+ N_XI0/XI9/XI12/NET35_XI0/XI9/XI12/MM11_g N_VDD_XI0/XI9/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI13/MM2 N_XI0/XI9/XI13/NET34_XI0/XI9/XI13/MM2_d
+ N_XI0/XI9/XI13/NET33_XI0/XI9/XI13/MM2_g N_VSS_XI0/XI9/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM3 N_XI0/XI9/XI13/NET33_XI0/XI9/XI13/MM3_d
+ N_WL<14>_XI0/XI9/XI13/MM3_g N_BLN<2>_XI0/XI9/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM0 N_XI0/XI9/XI13/NET34_XI0/XI9/XI13/MM0_d
+ N_WL<14>_XI0/XI9/XI13/MM0_g N_BL<2>_XI0/XI9/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM1 N_XI0/XI9/XI13/NET33_XI0/XI9/XI13/MM1_d
+ N_XI0/XI9/XI13/NET34_XI0/XI9/XI13/MM1_g N_VSS_XI0/XI9/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM9 N_XI0/XI9/XI13/NET36_XI0/XI9/XI13/MM9_d
+ N_WL<15>_XI0/XI9/XI13/MM9_g N_BL<2>_XI0/XI9/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM6 N_XI0/XI9/XI13/NET35_XI0/XI9/XI13/MM6_d
+ N_XI0/XI9/XI13/NET36_XI0/XI9/XI13/MM6_g N_VSS_XI0/XI9/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM7 N_XI0/XI9/XI13/NET36_XI0/XI9/XI13/MM7_d
+ N_XI0/XI9/XI13/NET35_XI0/XI9/XI13/MM7_g N_VSS_XI0/XI9/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM8 N_XI0/XI9/XI13/NET35_XI0/XI9/XI13/MM8_d
+ N_WL<15>_XI0/XI9/XI13/MM8_g N_BLN<2>_XI0/XI9/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI13/MM5 N_XI0/XI9/XI13/NET34_XI0/XI9/XI13/MM5_d
+ N_XI0/XI9/XI13/NET33_XI0/XI9/XI13/MM5_g N_VDD_XI0/XI9/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI13/MM4 N_XI0/XI9/XI13/NET33_XI0/XI9/XI13/MM4_d
+ N_XI0/XI9/XI13/NET34_XI0/XI9/XI13/MM4_g N_VDD_XI0/XI9/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI13/MM10 N_XI0/XI9/XI13/NET35_XI0/XI9/XI13/MM10_d
+ N_XI0/XI9/XI13/NET36_XI0/XI9/XI13/MM10_g N_VDD_XI0/XI9/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI13/MM11 N_XI0/XI9/XI13/NET36_XI0/XI9/XI13/MM11_d
+ N_XI0/XI9/XI13/NET35_XI0/XI9/XI13/MM11_g N_VDD_XI0/XI9/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI14/MM2 N_XI0/XI9/XI14/NET34_XI0/XI9/XI14/MM2_d
+ N_XI0/XI9/XI14/NET33_XI0/XI9/XI14/MM2_g N_VSS_XI0/XI9/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM3 N_XI0/XI9/XI14/NET33_XI0/XI9/XI14/MM3_d
+ N_WL<14>_XI0/XI9/XI14/MM3_g N_BLN<1>_XI0/XI9/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM0 N_XI0/XI9/XI14/NET34_XI0/XI9/XI14/MM0_d
+ N_WL<14>_XI0/XI9/XI14/MM0_g N_BL<1>_XI0/XI9/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM1 N_XI0/XI9/XI14/NET33_XI0/XI9/XI14/MM1_d
+ N_XI0/XI9/XI14/NET34_XI0/XI9/XI14/MM1_g N_VSS_XI0/XI9/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM9 N_XI0/XI9/XI14/NET36_XI0/XI9/XI14/MM9_d
+ N_WL<15>_XI0/XI9/XI14/MM9_g N_BL<1>_XI0/XI9/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM6 N_XI0/XI9/XI14/NET35_XI0/XI9/XI14/MM6_d
+ N_XI0/XI9/XI14/NET36_XI0/XI9/XI14/MM6_g N_VSS_XI0/XI9/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM7 N_XI0/XI9/XI14/NET36_XI0/XI9/XI14/MM7_d
+ N_XI0/XI9/XI14/NET35_XI0/XI9/XI14/MM7_g N_VSS_XI0/XI9/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM8 N_XI0/XI9/XI14/NET35_XI0/XI9/XI14/MM8_d
+ N_WL<15>_XI0/XI9/XI14/MM8_g N_BLN<1>_XI0/XI9/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI14/MM5 N_XI0/XI9/XI14/NET34_XI0/XI9/XI14/MM5_d
+ N_XI0/XI9/XI14/NET33_XI0/XI9/XI14/MM5_g N_VDD_XI0/XI9/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI14/MM4 N_XI0/XI9/XI14/NET33_XI0/XI9/XI14/MM4_d
+ N_XI0/XI9/XI14/NET34_XI0/XI9/XI14/MM4_g N_VDD_XI0/XI9/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI14/MM10 N_XI0/XI9/XI14/NET35_XI0/XI9/XI14/MM10_d
+ N_XI0/XI9/XI14/NET36_XI0/XI9/XI14/MM10_g N_VDD_XI0/XI9/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI14/MM11 N_XI0/XI9/XI14/NET36_XI0/XI9/XI14/MM11_d
+ N_XI0/XI9/XI14/NET35_XI0/XI9/XI14/MM11_g N_VDD_XI0/XI9/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI15/MM2 N_XI0/XI9/XI15/NET34_XI0/XI9/XI15/MM2_d
+ N_XI0/XI9/XI15/NET33_XI0/XI9/XI15/MM2_g N_VSS_XI0/XI9/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM3 N_XI0/XI9/XI15/NET33_XI0/XI9/XI15/MM3_d
+ N_WL<14>_XI0/XI9/XI15/MM3_g N_BLN<0>_XI0/XI9/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM0 N_XI0/XI9/XI15/NET34_XI0/XI9/XI15/MM0_d
+ N_WL<14>_XI0/XI9/XI15/MM0_g N_BL<0>_XI0/XI9/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM1 N_XI0/XI9/XI15/NET33_XI0/XI9/XI15/MM1_d
+ N_XI0/XI9/XI15/NET34_XI0/XI9/XI15/MM1_g N_VSS_XI0/XI9/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM9 N_XI0/XI9/XI15/NET36_XI0/XI9/XI15/MM9_d
+ N_WL<15>_XI0/XI9/XI15/MM9_g N_BL<0>_XI0/XI9/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM6 N_XI0/XI9/XI15/NET35_XI0/XI9/XI15/MM6_d
+ N_XI0/XI9/XI15/NET36_XI0/XI9/XI15/MM6_g N_VSS_XI0/XI9/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM7 N_XI0/XI9/XI15/NET36_XI0/XI9/XI15/MM7_d
+ N_XI0/XI9/XI15/NET35_XI0/XI9/XI15/MM7_g N_VSS_XI0/XI9/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM8 N_XI0/XI9/XI15/NET35_XI0/XI9/XI15/MM8_d
+ N_WL<15>_XI0/XI9/XI15/MM8_g N_BLN<0>_XI0/XI9/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/XI15/MM5 N_XI0/XI9/XI15/NET34_XI0/XI9/XI15/MM5_d
+ N_XI0/XI9/XI15/NET33_XI0/XI9/XI15/MM5_g N_VDD_XI0/XI9/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI15/MM4 N_XI0/XI9/XI15/NET33_XI0/XI9/XI15/MM4_d
+ N_XI0/XI9/XI15/NET34_XI0/XI9/XI15/MM4_g N_VDD_XI0/XI9/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI15/MM10 N_XI0/XI9/XI15/NET35_XI0/XI9/XI15/MM10_d
+ N_XI0/XI9/XI15/NET36_XI0/XI9/XI15/MM10_g N_VDD_XI0/XI9/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/XI15/MM11 N_XI0/XI9/XI15/NET36_XI0/XI9/XI15/MM11_d
+ N_XI0/XI9/XI15/NET35_XI0/XI9/XI15/MM11_g N_VDD_XI0/XI9/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI0/MM2 N_XI0/XI10/XI0/NET34_XI0/XI10/XI0/MM2_d
+ N_XI0/XI10/XI0/NET33_XI0/XI10/XI0/MM2_g N_VSS_XI0/XI10/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM3 N_XI0/XI10/XI0/NET33_XI0/XI10/XI0/MM3_d
+ N_WL<16>_XI0/XI10/XI0/MM3_g N_BLN<15>_XI0/XI10/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM0 N_XI0/XI10/XI0/NET34_XI0/XI10/XI0/MM0_d
+ N_WL<16>_XI0/XI10/XI0/MM0_g N_BL<15>_XI0/XI10/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM1 N_XI0/XI10/XI0/NET33_XI0/XI10/XI0/MM1_d
+ N_XI0/XI10/XI0/NET34_XI0/XI10/XI0/MM1_g N_VSS_XI0/XI10/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM9 N_XI0/XI10/XI0/NET36_XI0/XI10/XI0/MM9_d
+ N_WL<17>_XI0/XI10/XI0/MM9_g N_BL<15>_XI0/XI10/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM6 N_XI0/XI10/XI0/NET35_XI0/XI10/XI0/MM6_d
+ N_XI0/XI10/XI0/NET36_XI0/XI10/XI0/MM6_g N_VSS_XI0/XI10/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM7 N_XI0/XI10/XI0/NET36_XI0/XI10/XI0/MM7_d
+ N_XI0/XI10/XI0/NET35_XI0/XI10/XI0/MM7_g N_VSS_XI0/XI10/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM8 N_XI0/XI10/XI0/NET35_XI0/XI10/XI0/MM8_d
+ N_WL<17>_XI0/XI10/XI0/MM8_g N_BLN<15>_XI0/XI10/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI0/MM5 N_XI0/XI10/XI0/NET34_XI0/XI10/XI0/MM5_d
+ N_XI0/XI10/XI0/NET33_XI0/XI10/XI0/MM5_g N_VDD_XI0/XI10/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI0/MM4 N_XI0/XI10/XI0/NET33_XI0/XI10/XI0/MM4_d
+ N_XI0/XI10/XI0/NET34_XI0/XI10/XI0/MM4_g N_VDD_XI0/XI10/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI0/MM10 N_XI0/XI10/XI0/NET35_XI0/XI10/XI0/MM10_d
+ N_XI0/XI10/XI0/NET36_XI0/XI10/XI0/MM10_g N_VDD_XI0/XI10/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI0/MM11 N_XI0/XI10/XI0/NET36_XI0/XI10/XI0/MM11_d
+ N_XI0/XI10/XI0/NET35_XI0/XI10/XI0/MM11_g N_VDD_XI0/XI10/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI1/MM2 N_XI0/XI10/XI1/NET34_XI0/XI10/XI1/MM2_d
+ N_XI0/XI10/XI1/NET33_XI0/XI10/XI1/MM2_g N_VSS_XI0/XI10/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM3 N_XI0/XI10/XI1/NET33_XI0/XI10/XI1/MM3_d
+ N_WL<16>_XI0/XI10/XI1/MM3_g N_BLN<14>_XI0/XI10/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM0 N_XI0/XI10/XI1/NET34_XI0/XI10/XI1/MM0_d
+ N_WL<16>_XI0/XI10/XI1/MM0_g N_BL<14>_XI0/XI10/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM1 N_XI0/XI10/XI1/NET33_XI0/XI10/XI1/MM1_d
+ N_XI0/XI10/XI1/NET34_XI0/XI10/XI1/MM1_g N_VSS_XI0/XI10/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM9 N_XI0/XI10/XI1/NET36_XI0/XI10/XI1/MM9_d
+ N_WL<17>_XI0/XI10/XI1/MM9_g N_BL<14>_XI0/XI10/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM6 N_XI0/XI10/XI1/NET35_XI0/XI10/XI1/MM6_d
+ N_XI0/XI10/XI1/NET36_XI0/XI10/XI1/MM6_g N_VSS_XI0/XI10/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM7 N_XI0/XI10/XI1/NET36_XI0/XI10/XI1/MM7_d
+ N_XI0/XI10/XI1/NET35_XI0/XI10/XI1/MM7_g N_VSS_XI0/XI10/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM8 N_XI0/XI10/XI1/NET35_XI0/XI10/XI1/MM8_d
+ N_WL<17>_XI0/XI10/XI1/MM8_g N_BLN<14>_XI0/XI10/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI1/MM5 N_XI0/XI10/XI1/NET34_XI0/XI10/XI1/MM5_d
+ N_XI0/XI10/XI1/NET33_XI0/XI10/XI1/MM5_g N_VDD_XI0/XI10/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI1/MM4 N_XI0/XI10/XI1/NET33_XI0/XI10/XI1/MM4_d
+ N_XI0/XI10/XI1/NET34_XI0/XI10/XI1/MM4_g N_VDD_XI0/XI10/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI1/MM10 N_XI0/XI10/XI1/NET35_XI0/XI10/XI1/MM10_d
+ N_XI0/XI10/XI1/NET36_XI0/XI10/XI1/MM10_g N_VDD_XI0/XI10/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI1/MM11 N_XI0/XI10/XI1/NET36_XI0/XI10/XI1/MM11_d
+ N_XI0/XI10/XI1/NET35_XI0/XI10/XI1/MM11_g N_VDD_XI0/XI10/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI2/MM2 N_XI0/XI10/XI2/NET34_XI0/XI10/XI2/MM2_d
+ N_XI0/XI10/XI2/NET33_XI0/XI10/XI2/MM2_g N_VSS_XI0/XI10/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM3 N_XI0/XI10/XI2/NET33_XI0/XI10/XI2/MM3_d
+ N_WL<16>_XI0/XI10/XI2/MM3_g N_BLN<13>_XI0/XI10/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM0 N_XI0/XI10/XI2/NET34_XI0/XI10/XI2/MM0_d
+ N_WL<16>_XI0/XI10/XI2/MM0_g N_BL<13>_XI0/XI10/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM1 N_XI0/XI10/XI2/NET33_XI0/XI10/XI2/MM1_d
+ N_XI0/XI10/XI2/NET34_XI0/XI10/XI2/MM1_g N_VSS_XI0/XI10/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM9 N_XI0/XI10/XI2/NET36_XI0/XI10/XI2/MM9_d
+ N_WL<17>_XI0/XI10/XI2/MM9_g N_BL<13>_XI0/XI10/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM6 N_XI0/XI10/XI2/NET35_XI0/XI10/XI2/MM6_d
+ N_XI0/XI10/XI2/NET36_XI0/XI10/XI2/MM6_g N_VSS_XI0/XI10/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM7 N_XI0/XI10/XI2/NET36_XI0/XI10/XI2/MM7_d
+ N_XI0/XI10/XI2/NET35_XI0/XI10/XI2/MM7_g N_VSS_XI0/XI10/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM8 N_XI0/XI10/XI2/NET35_XI0/XI10/XI2/MM8_d
+ N_WL<17>_XI0/XI10/XI2/MM8_g N_BLN<13>_XI0/XI10/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI2/MM5 N_XI0/XI10/XI2/NET34_XI0/XI10/XI2/MM5_d
+ N_XI0/XI10/XI2/NET33_XI0/XI10/XI2/MM5_g N_VDD_XI0/XI10/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI2/MM4 N_XI0/XI10/XI2/NET33_XI0/XI10/XI2/MM4_d
+ N_XI0/XI10/XI2/NET34_XI0/XI10/XI2/MM4_g N_VDD_XI0/XI10/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI2/MM10 N_XI0/XI10/XI2/NET35_XI0/XI10/XI2/MM10_d
+ N_XI0/XI10/XI2/NET36_XI0/XI10/XI2/MM10_g N_VDD_XI0/XI10/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI2/MM11 N_XI0/XI10/XI2/NET36_XI0/XI10/XI2/MM11_d
+ N_XI0/XI10/XI2/NET35_XI0/XI10/XI2/MM11_g N_VDD_XI0/XI10/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI3/MM2 N_XI0/XI10/XI3/NET34_XI0/XI10/XI3/MM2_d
+ N_XI0/XI10/XI3/NET33_XI0/XI10/XI3/MM2_g N_VSS_XI0/XI10/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM3 N_XI0/XI10/XI3/NET33_XI0/XI10/XI3/MM3_d
+ N_WL<16>_XI0/XI10/XI3/MM3_g N_BLN<12>_XI0/XI10/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM0 N_XI0/XI10/XI3/NET34_XI0/XI10/XI3/MM0_d
+ N_WL<16>_XI0/XI10/XI3/MM0_g N_BL<12>_XI0/XI10/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM1 N_XI0/XI10/XI3/NET33_XI0/XI10/XI3/MM1_d
+ N_XI0/XI10/XI3/NET34_XI0/XI10/XI3/MM1_g N_VSS_XI0/XI10/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM9 N_XI0/XI10/XI3/NET36_XI0/XI10/XI3/MM9_d
+ N_WL<17>_XI0/XI10/XI3/MM9_g N_BL<12>_XI0/XI10/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM6 N_XI0/XI10/XI3/NET35_XI0/XI10/XI3/MM6_d
+ N_XI0/XI10/XI3/NET36_XI0/XI10/XI3/MM6_g N_VSS_XI0/XI10/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM7 N_XI0/XI10/XI3/NET36_XI0/XI10/XI3/MM7_d
+ N_XI0/XI10/XI3/NET35_XI0/XI10/XI3/MM7_g N_VSS_XI0/XI10/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM8 N_XI0/XI10/XI3/NET35_XI0/XI10/XI3/MM8_d
+ N_WL<17>_XI0/XI10/XI3/MM8_g N_BLN<12>_XI0/XI10/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI3/MM5 N_XI0/XI10/XI3/NET34_XI0/XI10/XI3/MM5_d
+ N_XI0/XI10/XI3/NET33_XI0/XI10/XI3/MM5_g N_VDD_XI0/XI10/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI3/MM4 N_XI0/XI10/XI3/NET33_XI0/XI10/XI3/MM4_d
+ N_XI0/XI10/XI3/NET34_XI0/XI10/XI3/MM4_g N_VDD_XI0/XI10/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI3/MM10 N_XI0/XI10/XI3/NET35_XI0/XI10/XI3/MM10_d
+ N_XI0/XI10/XI3/NET36_XI0/XI10/XI3/MM10_g N_VDD_XI0/XI10/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI3/MM11 N_XI0/XI10/XI3/NET36_XI0/XI10/XI3/MM11_d
+ N_XI0/XI10/XI3/NET35_XI0/XI10/XI3/MM11_g N_VDD_XI0/XI10/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI4/MM2 N_XI0/XI10/XI4/NET34_XI0/XI10/XI4/MM2_d
+ N_XI0/XI10/XI4/NET33_XI0/XI10/XI4/MM2_g N_VSS_XI0/XI10/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM3 N_XI0/XI10/XI4/NET33_XI0/XI10/XI4/MM3_d
+ N_WL<16>_XI0/XI10/XI4/MM3_g N_BLN<11>_XI0/XI10/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM0 N_XI0/XI10/XI4/NET34_XI0/XI10/XI4/MM0_d
+ N_WL<16>_XI0/XI10/XI4/MM0_g N_BL<11>_XI0/XI10/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM1 N_XI0/XI10/XI4/NET33_XI0/XI10/XI4/MM1_d
+ N_XI0/XI10/XI4/NET34_XI0/XI10/XI4/MM1_g N_VSS_XI0/XI10/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM9 N_XI0/XI10/XI4/NET36_XI0/XI10/XI4/MM9_d
+ N_WL<17>_XI0/XI10/XI4/MM9_g N_BL<11>_XI0/XI10/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM6 N_XI0/XI10/XI4/NET35_XI0/XI10/XI4/MM6_d
+ N_XI0/XI10/XI4/NET36_XI0/XI10/XI4/MM6_g N_VSS_XI0/XI10/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM7 N_XI0/XI10/XI4/NET36_XI0/XI10/XI4/MM7_d
+ N_XI0/XI10/XI4/NET35_XI0/XI10/XI4/MM7_g N_VSS_XI0/XI10/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM8 N_XI0/XI10/XI4/NET35_XI0/XI10/XI4/MM8_d
+ N_WL<17>_XI0/XI10/XI4/MM8_g N_BLN<11>_XI0/XI10/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI4/MM5 N_XI0/XI10/XI4/NET34_XI0/XI10/XI4/MM5_d
+ N_XI0/XI10/XI4/NET33_XI0/XI10/XI4/MM5_g N_VDD_XI0/XI10/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI4/MM4 N_XI0/XI10/XI4/NET33_XI0/XI10/XI4/MM4_d
+ N_XI0/XI10/XI4/NET34_XI0/XI10/XI4/MM4_g N_VDD_XI0/XI10/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI4/MM10 N_XI0/XI10/XI4/NET35_XI0/XI10/XI4/MM10_d
+ N_XI0/XI10/XI4/NET36_XI0/XI10/XI4/MM10_g N_VDD_XI0/XI10/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI4/MM11 N_XI0/XI10/XI4/NET36_XI0/XI10/XI4/MM11_d
+ N_XI0/XI10/XI4/NET35_XI0/XI10/XI4/MM11_g N_VDD_XI0/XI10/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI5/MM2 N_XI0/XI10/XI5/NET34_XI0/XI10/XI5/MM2_d
+ N_XI0/XI10/XI5/NET33_XI0/XI10/XI5/MM2_g N_VSS_XI0/XI10/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM3 N_XI0/XI10/XI5/NET33_XI0/XI10/XI5/MM3_d
+ N_WL<16>_XI0/XI10/XI5/MM3_g N_BLN<10>_XI0/XI10/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM0 N_XI0/XI10/XI5/NET34_XI0/XI10/XI5/MM0_d
+ N_WL<16>_XI0/XI10/XI5/MM0_g N_BL<10>_XI0/XI10/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM1 N_XI0/XI10/XI5/NET33_XI0/XI10/XI5/MM1_d
+ N_XI0/XI10/XI5/NET34_XI0/XI10/XI5/MM1_g N_VSS_XI0/XI10/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM9 N_XI0/XI10/XI5/NET36_XI0/XI10/XI5/MM9_d
+ N_WL<17>_XI0/XI10/XI5/MM9_g N_BL<10>_XI0/XI10/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM6 N_XI0/XI10/XI5/NET35_XI0/XI10/XI5/MM6_d
+ N_XI0/XI10/XI5/NET36_XI0/XI10/XI5/MM6_g N_VSS_XI0/XI10/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM7 N_XI0/XI10/XI5/NET36_XI0/XI10/XI5/MM7_d
+ N_XI0/XI10/XI5/NET35_XI0/XI10/XI5/MM7_g N_VSS_XI0/XI10/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM8 N_XI0/XI10/XI5/NET35_XI0/XI10/XI5/MM8_d
+ N_WL<17>_XI0/XI10/XI5/MM8_g N_BLN<10>_XI0/XI10/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI5/MM5 N_XI0/XI10/XI5/NET34_XI0/XI10/XI5/MM5_d
+ N_XI0/XI10/XI5/NET33_XI0/XI10/XI5/MM5_g N_VDD_XI0/XI10/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI5/MM4 N_XI0/XI10/XI5/NET33_XI0/XI10/XI5/MM4_d
+ N_XI0/XI10/XI5/NET34_XI0/XI10/XI5/MM4_g N_VDD_XI0/XI10/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI5/MM10 N_XI0/XI10/XI5/NET35_XI0/XI10/XI5/MM10_d
+ N_XI0/XI10/XI5/NET36_XI0/XI10/XI5/MM10_g N_VDD_XI0/XI10/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI5/MM11 N_XI0/XI10/XI5/NET36_XI0/XI10/XI5/MM11_d
+ N_XI0/XI10/XI5/NET35_XI0/XI10/XI5/MM11_g N_VDD_XI0/XI10/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI6/MM2 N_XI0/XI10/XI6/NET34_XI0/XI10/XI6/MM2_d
+ N_XI0/XI10/XI6/NET33_XI0/XI10/XI6/MM2_g N_VSS_XI0/XI10/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM3 N_XI0/XI10/XI6/NET33_XI0/XI10/XI6/MM3_d
+ N_WL<16>_XI0/XI10/XI6/MM3_g N_BLN<9>_XI0/XI10/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM0 N_XI0/XI10/XI6/NET34_XI0/XI10/XI6/MM0_d
+ N_WL<16>_XI0/XI10/XI6/MM0_g N_BL<9>_XI0/XI10/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM1 N_XI0/XI10/XI6/NET33_XI0/XI10/XI6/MM1_d
+ N_XI0/XI10/XI6/NET34_XI0/XI10/XI6/MM1_g N_VSS_XI0/XI10/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM9 N_XI0/XI10/XI6/NET36_XI0/XI10/XI6/MM9_d
+ N_WL<17>_XI0/XI10/XI6/MM9_g N_BL<9>_XI0/XI10/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM6 N_XI0/XI10/XI6/NET35_XI0/XI10/XI6/MM6_d
+ N_XI0/XI10/XI6/NET36_XI0/XI10/XI6/MM6_g N_VSS_XI0/XI10/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM7 N_XI0/XI10/XI6/NET36_XI0/XI10/XI6/MM7_d
+ N_XI0/XI10/XI6/NET35_XI0/XI10/XI6/MM7_g N_VSS_XI0/XI10/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM8 N_XI0/XI10/XI6/NET35_XI0/XI10/XI6/MM8_d
+ N_WL<17>_XI0/XI10/XI6/MM8_g N_BLN<9>_XI0/XI10/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI6/MM5 N_XI0/XI10/XI6/NET34_XI0/XI10/XI6/MM5_d
+ N_XI0/XI10/XI6/NET33_XI0/XI10/XI6/MM5_g N_VDD_XI0/XI10/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI6/MM4 N_XI0/XI10/XI6/NET33_XI0/XI10/XI6/MM4_d
+ N_XI0/XI10/XI6/NET34_XI0/XI10/XI6/MM4_g N_VDD_XI0/XI10/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI6/MM10 N_XI0/XI10/XI6/NET35_XI0/XI10/XI6/MM10_d
+ N_XI0/XI10/XI6/NET36_XI0/XI10/XI6/MM10_g N_VDD_XI0/XI10/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI6/MM11 N_XI0/XI10/XI6/NET36_XI0/XI10/XI6/MM11_d
+ N_XI0/XI10/XI6/NET35_XI0/XI10/XI6/MM11_g N_VDD_XI0/XI10/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI7/MM2 N_XI0/XI10/XI7/NET34_XI0/XI10/XI7/MM2_d
+ N_XI0/XI10/XI7/NET33_XI0/XI10/XI7/MM2_g N_VSS_XI0/XI10/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM3 N_XI0/XI10/XI7/NET33_XI0/XI10/XI7/MM3_d
+ N_WL<16>_XI0/XI10/XI7/MM3_g N_BLN<8>_XI0/XI10/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM0 N_XI0/XI10/XI7/NET34_XI0/XI10/XI7/MM0_d
+ N_WL<16>_XI0/XI10/XI7/MM0_g N_BL<8>_XI0/XI10/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM1 N_XI0/XI10/XI7/NET33_XI0/XI10/XI7/MM1_d
+ N_XI0/XI10/XI7/NET34_XI0/XI10/XI7/MM1_g N_VSS_XI0/XI10/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM9 N_XI0/XI10/XI7/NET36_XI0/XI10/XI7/MM9_d
+ N_WL<17>_XI0/XI10/XI7/MM9_g N_BL<8>_XI0/XI10/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM6 N_XI0/XI10/XI7/NET35_XI0/XI10/XI7/MM6_d
+ N_XI0/XI10/XI7/NET36_XI0/XI10/XI7/MM6_g N_VSS_XI0/XI10/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM7 N_XI0/XI10/XI7/NET36_XI0/XI10/XI7/MM7_d
+ N_XI0/XI10/XI7/NET35_XI0/XI10/XI7/MM7_g N_VSS_XI0/XI10/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM8 N_XI0/XI10/XI7/NET35_XI0/XI10/XI7/MM8_d
+ N_WL<17>_XI0/XI10/XI7/MM8_g N_BLN<8>_XI0/XI10/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI7/MM5 N_XI0/XI10/XI7/NET34_XI0/XI10/XI7/MM5_d
+ N_XI0/XI10/XI7/NET33_XI0/XI10/XI7/MM5_g N_VDD_XI0/XI10/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI7/MM4 N_XI0/XI10/XI7/NET33_XI0/XI10/XI7/MM4_d
+ N_XI0/XI10/XI7/NET34_XI0/XI10/XI7/MM4_g N_VDD_XI0/XI10/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI7/MM10 N_XI0/XI10/XI7/NET35_XI0/XI10/XI7/MM10_d
+ N_XI0/XI10/XI7/NET36_XI0/XI10/XI7/MM10_g N_VDD_XI0/XI10/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI7/MM11 N_XI0/XI10/XI7/NET36_XI0/XI10/XI7/MM11_d
+ N_XI0/XI10/XI7/NET35_XI0/XI10/XI7/MM11_g N_VDD_XI0/XI10/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI8/MM2 N_XI0/XI10/XI8/NET34_XI0/XI10/XI8/MM2_d
+ N_XI0/XI10/XI8/NET33_XI0/XI10/XI8/MM2_g N_VSS_XI0/XI10/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM3 N_XI0/XI10/XI8/NET33_XI0/XI10/XI8/MM3_d
+ N_WL<16>_XI0/XI10/XI8/MM3_g N_BLN<7>_XI0/XI10/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM0 N_XI0/XI10/XI8/NET34_XI0/XI10/XI8/MM0_d
+ N_WL<16>_XI0/XI10/XI8/MM0_g N_BL<7>_XI0/XI10/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM1 N_XI0/XI10/XI8/NET33_XI0/XI10/XI8/MM1_d
+ N_XI0/XI10/XI8/NET34_XI0/XI10/XI8/MM1_g N_VSS_XI0/XI10/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM9 N_XI0/XI10/XI8/NET36_XI0/XI10/XI8/MM9_d
+ N_WL<17>_XI0/XI10/XI8/MM9_g N_BL<7>_XI0/XI10/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM6 N_XI0/XI10/XI8/NET35_XI0/XI10/XI8/MM6_d
+ N_XI0/XI10/XI8/NET36_XI0/XI10/XI8/MM6_g N_VSS_XI0/XI10/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM7 N_XI0/XI10/XI8/NET36_XI0/XI10/XI8/MM7_d
+ N_XI0/XI10/XI8/NET35_XI0/XI10/XI8/MM7_g N_VSS_XI0/XI10/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM8 N_XI0/XI10/XI8/NET35_XI0/XI10/XI8/MM8_d
+ N_WL<17>_XI0/XI10/XI8/MM8_g N_BLN<7>_XI0/XI10/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI8/MM5 N_XI0/XI10/XI8/NET34_XI0/XI10/XI8/MM5_d
+ N_XI0/XI10/XI8/NET33_XI0/XI10/XI8/MM5_g N_VDD_XI0/XI10/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI8/MM4 N_XI0/XI10/XI8/NET33_XI0/XI10/XI8/MM4_d
+ N_XI0/XI10/XI8/NET34_XI0/XI10/XI8/MM4_g N_VDD_XI0/XI10/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI8/MM10 N_XI0/XI10/XI8/NET35_XI0/XI10/XI8/MM10_d
+ N_XI0/XI10/XI8/NET36_XI0/XI10/XI8/MM10_g N_VDD_XI0/XI10/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI8/MM11 N_XI0/XI10/XI8/NET36_XI0/XI10/XI8/MM11_d
+ N_XI0/XI10/XI8/NET35_XI0/XI10/XI8/MM11_g N_VDD_XI0/XI10/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI9/MM2 N_XI0/XI10/XI9/NET34_XI0/XI10/XI9/MM2_d
+ N_XI0/XI10/XI9/NET33_XI0/XI10/XI9/MM2_g N_VSS_XI0/XI10/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM3 N_XI0/XI10/XI9/NET33_XI0/XI10/XI9/MM3_d
+ N_WL<16>_XI0/XI10/XI9/MM3_g N_BLN<6>_XI0/XI10/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM0 N_XI0/XI10/XI9/NET34_XI0/XI10/XI9/MM0_d
+ N_WL<16>_XI0/XI10/XI9/MM0_g N_BL<6>_XI0/XI10/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM1 N_XI0/XI10/XI9/NET33_XI0/XI10/XI9/MM1_d
+ N_XI0/XI10/XI9/NET34_XI0/XI10/XI9/MM1_g N_VSS_XI0/XI10/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM9 N_XI0/XI10/XI9/NET36_XI0/XI10/XI9/MM9_d
+ N_WL<17>_XI0/XI10/XI9/MM9_g N_BL<6>_XI0/XI10/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM6 N_XI0/XI10/XI9/NET35_XI0/XI10/XI9/MM6_d
+ N_XI0/XI10/XI9/NET36_XI0/XI10/XI9/MM6_g N_VSS_XI0/XI10/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM7 N_XI0/XI10/XI9/NET36_XI0/XI10/XI9/MM7_d
+ N_XI0/XI10/XI9/NET35_XI0/XI10/XI9/MM7_g N_VSS_XI0/XI10/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM8 N_XI0/XI10/XI9/NET35_XI0/XI10/XI9/MM8_d
+ N_WL<17>_XI0/XI10/XI9/MM8_g N_BLN<6>_XI0/XI10/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI9/MM5 N_XI0/XI10/XI9/NET34_XI0/XI10/XI9/MM5_d
+ N_XI0/XI10/XI9/NET33_XI0/XI10/XI9/MM5_g N_VDD_XI0/XI10/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI9/MM4 N_XI0/XI10/XI9/NET33_XI0/XI10/XI9/MM4_d
+ N_XI0/XI10/XI9/NET34_XI0/XI10/XI9/MM4_g N_VDD_XI0/XI10/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI9/MM10 N_XI0/XI10/XI9/NET35_XI0/XI10/XI9/MM10_d
+ N_XI0/XI10/XI9/NET36_XI0/XI10/XI9/MM10_g N_VDD_XI0/XI10/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI9/MM11 N_XI0/XI10/XI9/NET36_XI0/XI10/XI9/MM11_d
+ N_XI0/XI10/XI9/NET35_XI0/XI10/XI9/MM11_g N_VDD_XI0/XI10/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI10/MM2 N_XI0/XI10/XI10/NET34_XI0/XI10/XI10/MM2_d
+ N_XI0/XI10/XI10/NET33_XI0/XI10/XI10/MM2_g N_VSS_XI0/XI10/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM3 N_XI0/XI10/XI10/NET33_XI0/XI10/XI10/MM3_d
+ N_WL<16>_XI0/XI10/XI10/MM3_g N_BLN<5>_XI0/XI10/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM0 N_XI0/XI10/XI10/NET34_XI0/XI10/XI10/MM0_d
+ N_WL<16>_XI0/XI10/XI10/MM0_g N_BL<5>_XI0/XI10/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM1 N_XI0/XI10/XI10/NET33_XI0/XI10/XI10/MM1_d
+ N_XI0/XI10/XI10/NET34_XI0/XI10/XI10/MM1_g N_VSS_XI0/XI10/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM9 N_XI0/XI10/XI10/NET36_XI0/XI10/XI10/MM9_d
+ N_WL<17>_XI0/XI10/XI10/MM9_g N_BL<5>_XI0/XI10/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM6 N_XI0/XI10/XI10/NET35_XI0/XI10/XI10/MM6_d
+ N_XI0/XI10/XI10/NET36_XI0/XI10/XI10/MM6_g N_VSS_XI0/XI10/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM7 N_XI0/XI10/XI10/NET36_XI0/XI10/XI10/MM7_d
+ N_XI0/XI10/XI10/NET35_XI0/XI10/XI10/MM7_g N_VSS_XI0/XI10/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM8 N_XI0/XI10/XI10/NET35_XI0/XI10/XI10/MM8_d
+ N_WL<17>_XI0/XI10/XI10/MM8_g N_BLN<5>_XI0/XI10/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI10/MM5 N_XI0/XI10/XI10/NET34_XI0/XI10/XI10/MM5_d
+ N_XI0/XI10/XI10/NET33_XI0/XI10/XI10/MM5_g N_VDD_XI0/XI10/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI10/MM4 N_XI0/XI10/XI10/NET33_XI0/XI10/XI10/MM4_d
+ N_XI0/XI10/XI10/NET34_XI0/XI10/XI10/MM4_g N_VDD_XI0/XI10/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI10/MM10 N_XI0/XI10/XI10/NET35_XI0/XI10/XI10/MM10_d
+ N_XI0/XI10/XI10/NET36_XI0/XI10/XI10/MM10_g N_VDD_XI0/XI10/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI10/MM11 N_XI0/XI10/XI10/NET36_XI0/XI10/XI10/MM11_d
+ N_XI0/XI10/XI10/NET35_XI0/XI10/XI10/MM11_g N_VDD_XI0/XI10/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI11/MM2 N_XI0/XI10/XI11/NET34_XI0/XI10/XI11/MM2_d
+ N_XI0/XI10/XI11/NET33_XI0/XI10/XI11/MM2_g N_VSS_XI0/XI10/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM3 N_XI0/XI10/XI11/NET33_XI0/XI10/XI11/MM3_d
+ N_WL<16>_XI0/XI10/XI11/MM3_g N_BLN<4>_XI0/XI10/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM0 N_XI0/XI10/XI11/NET34_XI0/XI10/XI11/MM0_d
+ N_WL<16>_XI0/XI10/XI11/MM0_g N_BL<4>_XI0/XI10/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM1 N_XI0/XI10/XI11/NET33_XI0/XI10/XI11/MM1_d
+ N_XI0/XI10/XI11/NET34_XI0/XI10/XI11/MM1_g N_VSS_XI0/XI10/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM9 N_XI0/XI10/XI11/NET36_XI0/XI10/XI11/MM9_d
+ N_WL<17>_XI0/XI10/XI11/MM9_g N_BL<4>_XI0/XI10/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM6 N_XI0/XI10/XI11/NET35_XI0/XI10/XI11/MM6_d
+ N_XI0/XI10/XI11/NET36_XI0/XI10/XI11/MM6_g N_VSS_XI0/XI10/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM7 N_XI0/XI10/XI11/NET36_XI0/XI10/XI11/MM7_d
+ N_XI0/XI10/XI11/NET35_XI0/XI10/XI11/MM7_g N_VSS_XI0/XI10/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM8 N_XI0/XI10/XI11/NET35_XI0/XI10/XI11/MM8_d
+ N_WL<17>_XI0/XI10/XI11/MM8_g N_BLN<4>_XI0/XI10/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI11/MM5 N_XI0/XI10/XI11/NET34_XI0/XI10/XI11/MM5_d
+ N_XI0/XI10/XI11/NET33_XI0/XI10/XI11/MM5_g N_VDD_XI0/XI10/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI11/MM4 N_XI0/XI10/XI11/NET33_XI0/XI10/XI11/MM4_d
+ N_XI0/XI10/XI11/NET34_XI0/XI10/XI11/MM4_g N_VDD_XI0/XI10/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI11/MM10 N_XI0/XI10/XI11/NET35_XI0/XI10/XI11/MM10_d
+ N_XI0/XI10/XI11/NET36_XI0/XI10/XI11/MM10_g N_VDD_XI0/XI10/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI11/MM11 N_XI0/XI10/XI11/NET36_XI0/XI10/XI11/MM11_d
+ N_XI0/XI10/XI11/NET35_XI0/XI10/XI11/MM11_g N_VDD_XI0/XI10/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI12/MM2 N_XI0/XI10/XI12/NET34_XI0/XI10/XI12/MM2_d
+ N_XI0/XI10/XI12/NET33_XI0/XI10/XI12/MM2_g N_VSS_XI0/XI10/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM3 N_XI0/XI10/XI12/NET33_XI0/XI10/XI12/MM3_d
+ N_WL<16>_XI0/XI10/XI12/MM3_g N_BLN<3>_XI0/XI10/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM0 N_XI0/XI10/XI12/NET34_XI0/XI10/XI12/MM0_d
+ N_WL<16>_XI0/XI10/XI12/MM0_g N_BL<3>_XI0/XI10/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM1 N_XI0/XI10/XI12/NET33_XI0/XI10/XI12/MM1_d
+ N_XI0/XI10/XI12/NET34_XI0/XI10/XI12/MM1_g N_VSS_XI0/XI10/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM9 N_XI0/XI10/XI12/NET36_XI0/XI10/XI12/MM9_d
+ N_WL<17>_XI0/XI10/XI12/MM9_g N_BL<3>_XI0/XI10/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM6 N_XI0/XI10/XI12/NET35_XI0/XI10/XI12/MM6_d
+ N_XI0/XI10/XI12/NET36_XI0/XI10/XI12/MM6_g N_VSS_XI0/XI10/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM7 N_XI0/XI10/XI12/NET36_XI0/XI10/XI12/MM7_d
+ N_XI0/XI10/XI12/NET35_XI0/XI10/XI12/MM7_g N_VSS_XI0/XI10/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM8 N_XI0/XI10/XI12/NET35_XI0/XI10/XI12/MM8_d
+ N_WL<17>_XI0/XI10/XI12/MM8_g N_BLN<3>_XI0/XI10/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI12/MM5 N_XI0/XI10/XI12/NET34_XI0/XI10/XI12/MM5_d
+ N_XI0/XI10/XI12/NET33_XI0/XI10/XI12/MM5_g N_VDD_XI0/XI10/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI12/MM4 N_XI0/XI10/XI12/NET33_XI0/XI10/XI12/MM4_d
+ N_XI0/XI10/XI12/NET34_XI0/XI10/XI12/MM4_g N_VDD_XI0/XI10/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI12/MM10 N_XI0/XI10/XI12/NET35_XI0/XI10/XI12/MM10_d
+ N_XI0/XI10/XI12/NET36_XI0/XI10/XI12/MM10_g N_VDD_XI0/XI10/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI12/MM11 N_XI0/XI10/XI12/NET36_XI0/XI10/XI12/MM11_d
+ N_XI0/XI10/XI12/NET35_XI0/XI10/XI12/MM11_g N_VDD_XI0/XI10/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI13/MM2 N_XI0/XI10/XI13/NET34_XI0/XI10/XI13/MM2_d
+ N_XI0/XI10/XI13/NET33_XI0/XI10/XI13/MM2_g N_VSS_XI0/XI10/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM3 N_XI0/XI10/XI13/NET33_XI0/XI10/XI13/MM3_d
+ N_WL<16>_XI0/XI10/XI13/MM3_g N_BLN<2>_XI0/XI10/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM0 N_XI0/XI10/XI13/NET34_XI0/XI10/XI13/MM0_d
+ N_WL<16>_XI0/XI10/XI13/MM0_g N_BL<2>_XI0/XI10/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM1 N_XI0/XI10/XI13/NET33_XI0/XI10/XI13/MM1_d
+ N_XI0/XI10/XI13/NET34_XI0/XI10/XI13/MM1_g N_VSS_XI0/XI10/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM9 N_XI0/XI10/XI13/NET36_XI0/XI10/XI13/MM9_d
+ N_WL<17>_XI0/XI10/XI13/MM9_g N_BL<2>_XI0/XI10/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM6 N_XI0/XI10/XI13/NET35_XI0/XI10/XI13/MM6_d
+ N_XI0/XI10/XI13/NET36_XI0/XI10/XI13/MM6_g N_VSS_XI0/XI10/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM7 N_XI0/XI10/XI13/NET36_XI0/XI10/XI13/MM7_d
+ N_XI0/XI10/XI13/NET35_XI0/XI10/XI13/MM7_g N_VSS_XI0/XI10/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM8 N_XI0/XI10/XI13/NET35_XI0/XI10/XI13/MM8_d
+ N_WL<17>_XI0/XI10/XI13/MM8_g N_BLN<2>_XI0/XI10/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI13/MM5 N_XI0/XI10/XI13/NET34_XI0/XI10/XI13/MM5_d
+ N_XI0/XI10/XI13/NET33_XI0/XI10/XI13/MM5_g N_VDD_XI0/XI10/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI13/MM4 N_XI0/XI10/XI13/NET33_XI0/XI10/XI13/MM4_d
+ N_XI0/XI10/XI13/NET34_XI0/XI10/XI13/MM4_g N_VDD_XI0/XI10/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI13/MM10 N_XI0/XI10/XI13/NET35_XI0/XI10/XI13/MM10_d
+ N_XI0/XI10/XI13/NET36_XI0/XI10/XI13/MM10_g N_VDD_XI0/XI10/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI13/MM11 N_XI0/XI10/XI13/NET36_XI0/XI10/XI13/MM11_d
+ N_XI0/XI10/XI13/NET35_XI0/XI10/XI13/MM11_g N_VDD_XI0/XI10/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI14/MM2 N_XI0/XI10/XI14/NET34_XI0/XI10/XI14/MM2_d
+ N_XI0/XI10/XI14/NET33_XI0/XI10/XI14/MM2_g N_VSS_XI0/XI10/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM3 N_XI0/XI10/XI14/NET33_XI0/XI10/XI14/MM3_d
+ N_WL<16>_XI0/XI10/XI14/MM3_g N_BLN<1>_XI0/XI10/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM0 N_XI0/XI10/XI14/NET34_XI0/XI10/XI14/MM0_d
+ N_WL<16>_XI0/XI10/XI14/MM0_g N_BL<1>_XI0/XI10/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM1 N_XI0/XI10/XI14/NET33_XI0/XI10/XI14/MM1_d
+ N_XI0/XI10/XI14/NET34_XI0/XI10/XI14/MM1_g N_VSS_XI0/XI10/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM9 N_XI0/XI10/XI14/NET36_XI0/XI10/XI14/MM9_d
+ N_WL<17>_XI0/XI10/XI14/MM9_g N_BL<1>_XI0/XI10/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM6 N_XI0/XI10/XI14/NET35_XI0/XI10/XI14/MM6_d
+ N_XI0/XI10/XI14/NET36_XI0/XI10/XI14/MM6_g N_VSS_XI0/XI10/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM7 N_XI0/XI10/XI14/NET36_XI0/XI10/XI14/MM7_d
+ N_XI0/XI10/XI14/NET35_XI0/XI10/XI14/MM7_g N_VSS_XI0/XI10/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM8 N_XI0/XI10/XI14/NET35_XI0/XI10/XI14/MM8_d
+ N_WL<17>_XI0/XI10/XI14/MM8_g N_BLN<1>_XI0/XI10/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI14/MM5 N_XI0/XI10/XI14/NET34_XI0/XI10/XI14/MM5_d
+ N_XI0/XI10/XI14/NET33_XI0/XI10/XI14/MM5_g N_VDD_XI0/XI10/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI14/MM4 N_XI0/XI10/XI14/NET33_XI0/XI10/XI14/MM4_d
+ N_XI0/XI10/XI14/NET34_XI0/XI10/XI14/MM4_g N_VDD_XI0/XI10/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI14/MM10 N_XI0/XI10/XI14/NET35_XI0/XI10/XI14/MM10_d
+ N_XI0/XI10/XI14/NET36_XI0/XI10/XI14/MM10_g N_VDD_XI0/XI10/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI14/MM11 N_XI0/XI10/XI14/NET36_XI0/XI10/XI14/MM11_d
+ N_XI0/XI10/XI14/NET35_XI0/XI10/XI14/MM11_g N_VDD_XI0/XI10/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI15/MM2 N_XI0/XI10/XI15/NET34_XI0/XI10/XI15/MM2_d
+ N_XI0/XI10/XI15/NET33_XI0/XI10/XI15/MM2_g N_VSS_XI0/XI10/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM3 N_XI0/XI10/XI15/NET33_XI0/XI10/XI15/MM3_d
+ N_WL<16>_XI0/XI10/XI15/MM3_g N_BLN<0>_XI0/XI10/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM0 N_XI0/XI10/XI15/NET34_XI0/XI10/XI15/MM0_d
+ N_WL<16>_XI0/XI10/XI15/MM0_g N_BL<0>_XI0/XI10/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM1 N_XI0/XI10/XI15/NET33_XI0/XI10/XI15/MM1_d
+ N_XI0/XI10/XI15/NET34_XI0/XI10/XI15/MM1_g N_VSS_XI0/XI10/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM9 N_XI0/XI10/XI15/NET36_XI0/XI10/XI15/MM9_d
+ N_WL<17>_XI0/XI10/XI15/MM9_g N_BL<0>_XI0/XI10/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM6 N_XI0/XI10/XI15/NET35_XI0/XI10/XI15/MM6_d
+ N_XI0/XI10/XI15/NET36_XI0/XI10/XI15/MM6_g N_VSS_XI0/XI10/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM7 N_XI0/XI10/XI15/NET36_XI0/XI10/XI15/MM7_d
+ N_XI0/XI10/XI15/NET35_XI0/XI10/XI15/MM7_g N_VSS_XI0/XI10/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM8 N_XI0/XI10/XI15/NET35_XI0/XI10/XI15/MM8_d
+ N_WL<17>_XI0/XI10/XI15/MM8_g N_BLN<0>_XI0/XI10/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/XI15/MM5 N_XI0/XI10/XI15/NET34_XI0/XI10/XI15/MM5_d
+ N_XI0/XI10/XI15/NET33_XI0/XI10/XI15/MM5_g N_VDD_XI0/XI10/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI15/MM4 N_XI0/XI10/XI15/NET33_XI0/XI10/XI15/MM4_d
+ N_XI0/XI10/XI15/NET34_XI0/XI10/XI15/MM4_g N_VDD_XI0/XI10/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI15/MM10 N_XI0/XI10/XI15/NET35_XI0/XI10/XI15/MM10_d
+ N_XI0/XI10/XI15/NET36_XI0/XI10/XI15/MM10_g N_VDD_XI0/XI10/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/XI15/MM11 N_XI0/XI10/XI15/NET36_XI0/XI10/XI15/MM11_d
+ N_XI0/XI10/XI15/NET35_XI0/XI10/XI15/MM11_g N_VDD_XI0/XI10/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI0/MM2 N_XI0/XI11/XI0/NET34_XI0/XI11/XI0/MM2_d
+ N_XI0/XI11/XI0/NET33_XI0/XI11/XI0/MM2_g N_VSS_XI0/XI11/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM3 N_XI0/XI11/XI0/NET33_XI0/XI11/XI0/MM3_d
+ N_WL<18>_XI0/XI11/XI0/MM3_g N_BLN<15>_XI0/XI11/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM0 N_XI0/XI11/XI0/NET34_XI0/XI11/XI0/MM0_d
+ N_WL<18>_XI0/XI11/XI0/MM0_g N_BL<15>_XI0/XI11/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM1 N_XI0/XI11/XI0/NET33_XI0/XI11/XI0/MM1_d
+ N_XI0/XI11/XI0/NET34_XI0/XI11/XI0/MM1_g N_VSS_XI0/XI11/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM9 N_XI0/XI11/XI0/NET36_XI0/XI11/XI0/MM9_d
+ N_WL<19>_XI0/XI11/XI0/MM9_g N_BL<15>_XI0/XI11/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM6 N_XI0/XI11/XI0/NET35_XI0/XI11/XI0/MM6_d
+ N_XI0/XI11/XI0/NET36_XI0/XI11/XI0/MM6_g N_VSS_XI0/XI11/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM7 N_XI0/XI11/XI0/NET36_XI0/XI11/XI0/MM7_d
+ N_XI0/XI11/XI0/NET35_XI0/XI11/XI0/MM7_g N_VSS_XI0/XI11/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM8 N_XI0/XI11/XI0/NET35_XI0/XI11/XI0/MM8_d
+ N_WL<19>_XI0/XI11/XI0/MM8_g N_BLN<15>_XI0/XI11/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI0/MM5 N_XI0/XI11/XI0/NET34_XI0/XI11/XI0/MM5_d
+ N_XI0/XI11/XI0/NET33_XI0/XI11/XI0/MM5_g N_VDD_XI0/XI11/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI0/MM4 N_XI0/XI11/XI0/NET33_XI0/XI11/XI0/MM4_d
+ N_XI0/XI11/XI0/NET34_XI0/XI11/XI0/MM4_g N_VDD_XI0/XI11/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI0/MM10 N_XI0/XI11/XI0/NET35_XI0/XI11/XI0/MM10_d
+ N_XI0/XI11/XI0/NET36_XI0/XI11/XI0/MM10_g N_VDD_XI0/XI11/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI0/MM11 N_XI0/XI11/XI0/NET36_XI0/XI11/XI0/MM11_d
+ N_XI0/XI11/XI0/NET35_XI0/XI11/XI0/MM11_g N_VDD_XI0/XI11/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI1/MM2 N_XI0/XI11/XI1/NET34_XI0/XI11/XI1/MM2_d
+ N_XI0/XI11/XI1/NET33_XI0/XI11/XI1/MM2_g N_VSS_XI0/XI11/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM3 N_XI0/XI11/XI1/NET33_XI0/XI11/XI1/MM3_d
+ N_WL<18>_XI0/XI11/XI1/MM3_g N_BLN<14>_XI0/XI11/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM0 N_XI0/XI11/XI1/NET34_XI0/XI11/XI1/MM0_d
+ N_WL<18>_XI0/XI11/XI1/MM0_g N_BL<14>_XI0/XI11/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM1 N_XI0/XI11/XI1/NET33_XI0/XI11/XI1/MM1_d
+ N_XI0/XI11/XI1/NET34_XI0/XI11/XI1/MM1_g N_VSS_XI0/XI11/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM9 N_XI0/XI11/XI1/NET36_XI0/XI11/XI1/MM9_d
+ N_WL<19>_XI0/XI11/XI1/MM9_g N_BL<14>_XI0/XI11/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM6 N_XI0/XI11/XI1/NET35_XI0/XI11/XI1/MM6_d
+ N_XI0/XI11/XI1/NET36_XI0/XI11/XI1/MM6_g N_VSS_XI0/XI11/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM7 N_XI0/XI11/XI1/NET36_XI0/XI11/XI1/MM7_d
+ N_XI0/XI11/XI1/NET35_XI0/XI11/XI1/MM7_g N_VSS_XI0/XI11/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM8 N_XI0/XI11/XI1/NET35_XI0/XI11/XI1/MM8_d
+ N_WL<19>_XI0/XI11/XI1/MM8_g N_BLN<14>_XI0/XI11/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI1/MM5 N_XI0/XI11/XI1/NET34_XI0/XI11/XI1/MM5_d
+ N_XI0/XI11/XI1/NET33_XI0/XI11/XI1/MM5_g N_VDD_XI0/XI11/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI1/MM4 N_XI0/XI11/XI1/NET33_XI0/XI11/XI1/MM4_d
+ N_XI0/XI11/XI1/NET34_XI0/XI11/XI1/MM4_g N_VDD_XI0/XI11/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI1/MM10 N_XI0/XI11/XI1/NET35_XI0/XI11/XI1/MM10_d
+ N_XI0/XI11/XI1/NET36_XI0/XI11/XI1/MM10_g N_VDD_XI0/XI11/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI1/MM11 N_XI0/XI11/XI1/NET36_XI0/XI11/XI1/MM11_d
+ N_XI0/XI11/XI1/NET35_XI0/XI11/XI1/MM11_g N_VDD_XI0/XI11/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI2/MM2 N_XI0/XI11/XI2/NET34_XI0/XI11/XI2/MM2_d
+ N_XI0/XI11/XI2/NET33_XI0/XI11/XI2/MM2_g N_VSS_XI0/XI11/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM3 N_XI0/XI11/XI2/NET33_XI0/XI11/XI2/MM3_d
+ N_WL<18>_XI0/XI11/XI2/MM3_g N_BLN<13>_XI0/XI11/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM0 N_XI0/XI11/XI2/NET34_XI0/XI11/XI2/MM0_d
+ N_WL<18>_XI0/XI11/XI2/MM0_g N_BL<13>_XI0/XI11/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM1 N_XI0/XI11/XI2/NET33_XI0/XI11/XI2/MM1_d
+ N_XI0/XI11/XI2/NET34_XI0/XI11/XI2/MM1_g N_VSS_XI0/XI11/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM9 N_XI0/XI11/XI2/NET36_XI0/XI11/XI2/MM9_d
+ N_WL<19>_XI0/XI11/XI2/MM9_g N_BL<13>_XI0/XI11/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM6 N_XI0/XI11/XI2/NET35_XI0/XI11/XI2/MM6_d
+ N_XI0/XI11/XI2/NET36_XI0/XI11/XI2/MM6_g N_VSS_XI0/XI11/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM7 N_XI0/XI11/XI2/NET36_XI0/XI11/XI2/MM7_d
+ N_XI0/XI11/XI2/NET35_XI0/XI11/XI2/MM7_g N_VSS_XI0/XI11/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM8 N_XI0/XI11/XI2/NET35_XI0/XI11/XI2/MM8_d
+ N_WL<19>_XI0/XI11/XI2/MM8_g N_BLN<13>_XI0/XI11/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI2/MM5 N_XI0/XI11/XI2/NET34_XI0/XI11/XI2/MM5_d
+ N_XI0/XI11/XI2/NET33_XI0/XI11/XI2/MM5_g N_VDD_XI0/XI11/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI2/MM4 N_XI0/XI11/XI2/NET33_XI0/XI11/XI2/MM4_d
+ N_XI0/XI11/XI2/NET34_XI0/XI11/XI2/MM4_g N_VDD_XI0/XI11/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI2/MM10 N_XI0/XI11/XI2/NET35_XI0/XI11/XI2/MM10_d
+ N_XI0/XI11/XI2/NET36_XI0/XI11/XI2/MM10_g N_VDD_XI0/XI11/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI2/MM11 N_XI0/XI11/XI2/NET36_XI0/XI11/XI2/MM11_d
+ N_XI0/XI11/XI2/NET35_XI0/XI11/XI2/MM11_g N_VDD_XI0/XI11/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI3/MM2 N_XI0/XI11/XI3/NET34_XI0/XI11/XI3/MM2_d
+ N_XI0/XI11/XI3/NET33_XI0/XI11/XI3/MM2_g N_VSS_XI0/XI11/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM3 N_XI0/XI11/XI3/NET33_XI0/XI11/XI3/MM3_d
+ N_WL<18>_XI0/XI11/XI3/MM3_g N_BLN<12>_XI0/XI11/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM0 N_XI0/XI11/XI3/NET34_XI0/XI11/XI3/MM0_d
+ N_WL<18>_XI0/XI11/XI3/MM0_g N_BL<12>_XI0/XI11/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM1 N_XI0/XI11/XI3/NET33_XI0/XI11/XI3/MM1_d
+ N_XI0/XI11/XI3/NET34_XI0/XI11/XI3/MM1_g N_VSS_XI0/XI11/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM9 N_XI0/XI11/XI3/NET36_XI0/XI11/XI3/MM9_d
+ N_WL<19>_XI0/XI11/XI3/MM9_g N_BL<12>_XI0/XI11/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM6 N_XI0/XI11/XI3/NET35_XI0/XI11/XI3/MM6_d
+ N_XI0/XI11/XI3/NET36_XI0/XI11/XI3/MM6_g N_VSS_XI0/XI11/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM7 N_XI0/XI11/XI3/NET36_XI0/XI11/XI3/MM7_d
+ N_XI0/XI11/XI3/NET35_XI0/XI11/XI3/MM7_g N_VSS_XI0/XI11/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM8 N_XI0/XI11/XI3/NET35_XI0/XI11/XI3/MM8_d
+ N_WL<19>_XI0/XI11/XI3/MM8_g N_BLN<12>_XI0/XI11/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI3/MM5 N_XI0/XI11/XI3/NET34_XI0/XI11/XI3/MM5_d
+ N_XI0/XI11/XI3/NET33_XI0/XI11/XI3/MM5_g N_VDD_XI0/XI11/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI3/MM4 N_XI0/XI11/XI3/NET33_XI0/XI11/XI3/MM4_d
+ N_XI0/XI11/XI3/NET34_XI0/XI11/XI3/MM4_g N_VDD_XI0/XI11/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI3/MM10 N_XI0/XI11/XI3/NET35_XI0/XI11/XI3/MM10_d
+ N_XI0/XI11/XI3/NET36_XI0/XI11/XI3/MM10_g N_VDD_XI0/XI11/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI3/MM11 N_XI0/XI11/XI3/NET36_XI0/XI11/XI3/MM11_d
+ N_XI0/XI11/XI3/NET35_XI0/XI11/XI3/MM11_g N_VDD_XI0/XI11/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI4/MM2 N_XI0/XI11/XI4/NET34_XI0/XI11/XI4/MM2_d
+ N_XI0/XI11/XI4/NET33_XI0/XI11/XI4/MM2_g N_VSS_XI0/XI11/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM3 N_XI0/XI11/XI4/NET33_XI0/XI11/XI4/MM3_d
+ N_WL<18>_XI0/XI11/XI4/MM3_g N_BLN<11>_XI0/XI11/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM0 N_XI0/XI11/XI4/NET34_XI0/XI11/XI4/MM0_d
+ N_WL<18>_XI0/XI11/XI4/MM0_g N_BL<11>_XI0/XI11/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM1 N_XI0/XI11/XI4/NET33_XI0/XI11/XI4/MM1_d
+ N_XI0/XI11/XI4/NET34_XI0/XI11/XI4/MM1_g N_VSS_XI0/XI11/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM9 N_XI0/XI11/XI4/NET36_XI0/XI11/XI4/MM9_d
+ N_WL<19>_XI0/XI11/XI4/MM9_g N_BL<11>_XI0/XI11/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM6 N_XI0/XI11/XI4/NET35_XI0/XI11/XI4/MM6_d
+ N_XI0/XI11/XI4/NET36_XI0/XI11/XI4/MM6_g N_VSS_XI0/XI11/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM7 N_XI0/XI11/XI4/NET36_XI0/XI11/XI4/MM7_d
+ N_XI0/XI11/XI4/NET35_XI0/XI11/XI4/MM7_g N_VSS_XI0/XI11/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM8 N_XI0/XI11/XI4/NET35_XI0/XI11/XI4/MM8_d
+ N_WL<19>_XI0/XI11/XI4/MM8_g N_BLN<11>_XI0/XI11/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI4/MM5 N_XI0/XI11/XI4/NET34_XI0/XI11/XI4/MM5_d
+ N_XI0/XI11/XI4/NET33_XI0/XI11/XI4/MM5_g N_VDD_XI0/XI11/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI4/MM4 N_XI0/XI11/XI4/NET33_XI0/XI11/XI4/MM4_d
+ N_XI0/XI11/XI4/NET34_XI0/XI11/XI4/MM4_g N_VDD_XI0/XI11/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI4/MM10 N_XI0/XI11/XI4/NET35_XI0/XI11/XI4/MM10_d
+ N_XI0/XI11/XI4/NET36_XI0/XI11/XI4/MM10_g N_VDD_XI0/XI11/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI4/MM11 N_XI0/XI11/XI4/NET36_XI0/XI11/XI4/MM11_d
+ N_XI0/XI11/XI4/NET35_XI0/XI11/XI4/MM11_g N_VDD_XI0/XI11/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI5/MM2 N_XI0/XI11/XI5/NET34_XI0/XI11/XI5/MM2_d
+ N_XI0/XI11/XI5/NET33_XI0/XI11/XI5/MM2_g N_VSS_XI0/XI11/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM3 N_XI0/XI11/XI5/NET33_XI0/XI11/XI5/MM3_d
+ N_WL<18>_XI0/XI11/XI5/MM3_g N_BLN<10>_XI0/XI11/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM0 N_XI0/XI11/XI5/NET34_XI0/XI11/XI5/MM0_d
+ N_WL<18>_XI0/XI11/XI5/MM0_g N_BL<10>_XI0/XI11/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM1 N_XI0/XI11/XI5/NET33_XI0/XI11/XI5/MM1_d
+ N_XI0/XI11/XI5/NET34_XI0/XI11/XI5/MM1_g N_VSS_XI0/XI11/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM9 N_XI0/XI11/XI5/NET36_XI0/XI11/XI5/MM9_d
+ N_WL<19>_XI0/XI11/XI5/MM9_g N_BL<10>_XI0/XI11/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM6 N_XI0/XI11/XI5/NET35_XI0/XI11/XI5/MM6_d
+ N_XI0/XI11/XI5/NET36_XI0/XI11/XI5/MM6_g N_VSS_XI0/XI11/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM7 N_XI0/XI11/XI5/NET36_XI0/XI11/XI5/MM7_d
+ N_XI0/XI11/XI5/NET35_XI0/XI11/XI5/MM7_g N_VSS_XI0/XI11/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM8 N_XI0/XI11/XI5/NET35_XI0/XI11/XI5/MM8_d
+ N_WL<19>_XI0/XI11/XI5/MM8_g N_BLN<10>_XI0/XI11/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI5/MM5 N_XI0/XI11/XI5/NET34_XI0/XI11/XI5/MM5_d
+ N_XI0/XI11/XI5/NET33_XI0/XI11/XI5/MM5_g N_VDD_XI0/XI11/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI5/MM4 N_XI0/XI11/XI5/NET33_XI0/XI11/XI5/MM4_d
+ N_XI0/XI11/XI5/NET34_XI0/XI11/XI5/MM4_g N_VDD_XI0/XI11/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI5/MM10 N_XI0/XI11/XI5/NET35_XI0/XI11/XI5/MM10_d
+ N_XI0/XI11/XI5/NET36_XI0/XI11/XI5/MM10_g N_VDD_XI0/XI11/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI5/MM11 N_XI0/XI11/XI5/NET36_XI0/XI11/XI5/MM11_d
+ N_XI0/XI11/XI5/NET35_XI0/XI11/XI5/MM11_g N_VDD_XI0/XI11/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI6/MM2 N_XI0/XI11/XI6/NET34_XI0/XI11/XI6/MM2_d
+ N_XI0/XI11/XI6/NET33_XI0/XI11/XI6/MM2_g N_VSS_XI0/XI11/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM3 N_XI0/XI11/XI6/NET33_XI0/XI11/XI6/MM3_d
+ N_WL<18>_XI0/XI11/XI6/MM3_g N_BLN<9>_XI0/XI11/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM0 N_XI0/XI11/XI6/NET34_XI0/XI11/XI6/MM0_d
+ N_WL<18>_XI0/XI11/XI6/MM0_g N_BL<9>_XI0/XI11/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM1 N_XI0/XI11/XI6/NET33_XI0/XI11/XI6/MM1_d
+ N_XI0/XI11/XI6/NET34_XI0/XI11/XI6/MM1_g N_VSS_XI0/XI11/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM9 N_XI0/XI11/XI6/NET36_XI0/XI11/XI6/MM9_d
+ N_WL<19>_XI0/XI11/XI6/MM9_g N_BL<9>_XI0/XI11/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM6 N_XI0/XI11/XI6/NET35_XI0/XI11/XI6/MM6_d
+ N_XI0/XI11/XI6/NET36_XI0/XI11/XI6/MM6_g N_VSS_XI0/XI11/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM7 N_XI0/XI11/XI6/NET36_XI0/XI11/XI6/MM7_d
+ N_XI0/XI11/XI6/NET35_XI0/XI11/XI6/MM7_g N_VSS_XI0/XI11/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM8 N_XI0/XI11/XI6/NET35_XI0/XI11/XI6/MM8_d
+ N_WL<19>_XI0/XI11/XI6/MM8_g N_BLN<9>_XI0/XI11/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI6/MM5 N_XI0/XI11/XI6/NET34_XI0/XI11/XI6/MM5_d
+ N_XI0/XI11/XI6/NET33_XI0/XI11/XI6/MM5_g N_VDD_XI0/XI11/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI6/MM4 N_XI0/XI11/XI6/NET33_XI0/XI11/XI6/MM4_d
+ N_XI0/XI11/XI6/NET34_XI0/XI11/XI6/MM4_g N_VDD_XI0/XI11/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI6/MM10 N_XI0/XI11/XI6/NET35_XI0/XI11/XI6/MM10_d
+ N_XI0/XI11/XI6/NET36_XI0/XI11/XI6/MM10_g N_VDD_XI0/XI11/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI6/MM11 N_XI0/XI11/XI6/NET36_XI0/XI11/XI6/MM11_d
+ N_XI0/XI11/XI6/NET35_XI0/XI11/XI6/MM11_g N_VDD_XI0/XI11/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI7/MM2 N_XI0/XI11/XI7/NET34_XI0/XI11/XI7/MM2_d
+ N_XI0/XI11/XI7/NET33_XI0/XI11/XI7/MM2_g N_VSS_XI0/XI11/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM3 N_XI0/XI11/XI7/NET33_XI0/XI11/XI7/MM3_d
+ N_WL<18>_XI0/XI11/XI7/MM3_g N_BLN<8>_XI0/XI11/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM0 N_XI0/XI11/XI7/NET34_XI0/XI11/XI7/MM0_d
+ N_WL<18>_XI0/XI11/XI7/MM0_g N_BL<8>_XI0/XI11/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM1 N_XI0/XI11/XI7/NET33_XI0/XI11/XI7/MM1_d
+ N_XI0/XI11/XI7/NET34_XI0/XI11/XI7/MM1_g N_VSS_XI0/XI11/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM9 N_XI0/XI11/XI7/NET36_XI0/XI11/XI7/MM9_d
+ N_WL<19>_XI0/XI11/XI7/MM9_g N_BL<8>_XI0/XI11/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM6 N_XI0/XI11/XI7/NET35_XI0/XI11/XI7/MM6_d
+ N_XI0/XI11/XI7/NET36_XI0/XI11/XI7/MM6_g N_VSS_XI0/XI11/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM7 N_XI0/XI11/XI7/NET36_XI0/XI11/XI7/MM7_d
+ N_XI0/XI11/XI7/NET35_XI0/XI11/XI7/MM7_g N_VSS_XI0/XI11/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM8 N_XI0/XI11/XI7/NET35_XI0/XI11/XI7/MM8_d
+ N_WL<19>_XI0/XI11/XI7/MM8_g N_BLN<8>_XI0/XI11/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI7/MM5 N_XI0/XI11/XI7/NET34_XI0/XI11/XI7/MM5_d
+ N_XI0/XI11/XI7/NET33_XI0/XI11/XI7/MM5_g N_VDD_XI0/XI11/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI7/MM4 N_XI0/XI11/XI7/NET33_XI0/XI11/XI7/MM4_d
+ N_XI0/XI11/XI7/NET34_XI0/XI11/XI7/MM4_g N_VDD_XI0/XI11/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI7/MM10 N_XI0/XI11/XI7/NET35_XI0/XI11/XI7/MM10_d
+ N_XI0/XI11/XI7/NET36_XI0/XI11/XI7/MM10_g N_VDD_XI0/XI11/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI7/MM11 N_XI0/XI11/XI7/NET36_XI0/XI11/XI7/MM11_d
+ N_XI0/XI11/XI7/NET35_XI0/XI11/XI7/MM11_g N_VDD_XI0/XI11/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI8/MM2 N_XI0/XI11/XI8/NET34_XI0/XI11/XI8/MM2_d
+ N_XI0/XI11/XI8/NET33_XI0/XI11/XI8/MM2_g N_VSS_XI0/XI11/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM3 N_XI0/XI11/XI8/NET33_XI0/XI11/XI8/MM3_d
+ N_WL<18>_XI0/XI11/XI8/MM3_g N_BLN<7>_XI0/XI11/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM0 N_XI0/XI11/XI8/NET34_XI0/XI11/XI8/MM0_d
+ N_WL<18>_XI0/XI11/XI8/MM0_g N_BL<7>_XI0/XI11/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM1 N_XI0/XI11/XI8/NET33_XI0/XI11/XI8/MM1_d
+ N_XI0/XI11/XI8/NET34_XI0/XI11/XI8/MM1_g N_VSS_XI0/XI11/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM9 N_XI0/XI11/XI8/NET36_XI0/XI11/XI8/MM9_d
+ N_WL<19>_XI0/XI11/XI8/MM9_g N_BL<7>_XI0/XI11/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM6 N_XI0/XI11/XI8/NET35_XI0/XI11/XI8/MM6_d
+ N_XI0/XI11/XI8/NET36_XI0/XI11/XI8/MM6_g N_VSS_XI0/XI11/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM7 N_XI0/XI11/XI8/NET36_XI0/XI11/XI8/MM7_d
+ N_XI0/XI11/XI8/NET35_XI0/XI11/XI8/MM7_g N_VSS_XI0/XI11/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM8 N_XI0/XI11/XI8/NET35_XI0/XI11/XI8/MM8_d
+ N_WL<19>_XI0/XI11/XI8/MM8_g N_BLN<7>_XI0/XI11/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI8/MM5 N_XI0/XI11/XI8/NET34_XI0/XI11/XI8/MM5_d
+ N_XI0/XI11/XI8/NET33_XI0/XI11/XI8/MM5_g N_VDD_XI0/XI11/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI8/MM4 N_XI0/XI11/XI8/NET33_XI0/XI11/XI8/MM4_d
+ N_XI0/XI11/XI8/NET34_XI0/XI11/XI8/MM4_g N_VDD_XI0/XI11/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI8/MM10 N_XI0/XI11/XI8/NET35_XI0/XI11/XI8/MM10_d
+ N_XI0/XI11/XI8/NET36_XI0/XI11/XI8/MM10_g N_VDD_XI0/XI11/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI8/MM11 N_XI0/XI11/XI8/NET36_XI0/XI11/XI8/MM11_d
+ N_XI0/XI11/XI8/NET35_XI0/XI11/XI8/MM11_g N_VDD_XI0/XI11/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI9/MM2 N_XI0/XI11/XI9/NET34_XI0/XI11/XI9/MM2_d
+ N_XI0/XI11/XI9/NET33_XI0/XI11/XI9/MM2_g N_VSS_XI0/XI11/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM3 N_XI0/XI11/XI9/NET33_XI0/XI11/XI9/MM3_d
+ N_WL<18>_XI0/XI11/XI9/MM3_g N_BLN<6>_XI0/XI11/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM0 N_XI0/XI11/XI9/NET34_XI0/XI11/XI9/MM0_d
+ N_WL<18>_XI0/XI11/XI9/MM0_g N_BL<6>_XI0/XI11/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM1 N_XI0/XI11/XI9/NET33_XI0/XI11/XI9/MM1_d
+ N_XI0/XI11/XI9/NET34_XI0/XI11/XI9/MM1_g N_VSS_XI0/XI11/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM9 N_XI0/XI11/XI9/NET36_XI0/XI11/XI9/MM9_d
+ N_WL<19>_XI0/XI11/XI9/MM9_g N_BL<6>_XI0/XI11/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM6 N_XI0/XI11/XI9/NET35_XI0/XI11/XI9/MM6_d
+ N_XI0/XI11/XI9/NET36_XI0/XI11/XI9/MM6_g N_VSS_XI0/XI11/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM7 N_XI0/XI11/XI9/NET36_XI0/XI11/XI9/MM7_d
+ N_XI0/XI11/XI9/NET35_XI0/XI11/XI9/MM7_g N_VSS_XI0/XI11/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM8 N_XI0/XI11/XI9/NET35_XI0/XI11/XI9/MM8_d
+ N_WL<19>_XI0/XI11/XI9/MM8_g N_BLN<6>_XI0/XI11/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI9/MM5 N_XI0/XI11/XI9/NET34_XI0/XI11/XI9/MM5_d
+ N_XI0/XI11/XI9/NET33_XI0/XI11/XI9/MM5_g N_VDD_XI0/XI11/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI9/MM4 N_XI0/XI11/XI9/NET33_XI0/XI11/XI9/MM4_d
+ N_XI0/XI11/XI9/NET34_XI0/XI11/XI9/MM4_g N_VDD_XI0/XI11/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI9/MM10 N_XI0/XI11/XI9/NET35_XI0/XI11/XI9/MM10_d
+ N_XI0/XI11/XI9/NET36_XI0/XI11/XI9/MM10_g N_VDD_XI0/XI11/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI9/MM11 N_XI0/XI11/XI9/NET36_XI0/XI11/XI9/MM11_d
+ N_XI0/XI11/XI9/NET35_XI0/XI11/XI9/MM11_g N_VDD_XI0/XI11/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI10/MM2 N_XI0/XI11/XI10/NET34_XI0/XI11/XI10/MM2_d
+ N_XI0/XI11/XI10/NET33_XI0/XI11/XI10/MM2_g N_VSS_XI0/XI11/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM3 N_XI0/XI11/XI10/NET33_XI0/XI11/XI10/MM3_d
+ N_WL<18>_XI0/XI11/XI10/MM3_g N_BLN<5>_XI0/XI11/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM0 N_XI0/XI11/XI10/NET34_XI0/XI11/XI10/MM0_d
+ N_WL<18>_XI0/XI11/XI10/MM0_g N_BL<5>_XI0/XI11/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM1 N_XI0/XI11/XI10/NET33_XI0/XI11/XI10/MM1_d
+ N_XI0/XI11/XI10/NET34_XI0/XI11/XI10/MM1_g N_VSS_XI0/XI11/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM9 N_XI0/XI11/XI10/NET36_XI0/XI11/XI10/MM9_d
+ N_WL<19>_XI0/XI11/XI10/MM9_g N_BL<5>_XI0/XI11/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM6 N_XI0/XI11/XI10/NET35_XI0/XI11/XI10/MM6_d
+ N_XI0/XI11/XI10/NET36_XI0/XI11/XI10/MM6_g N_VSS_XI0/XI11/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM7 N_XI0/XI11/XI10/NET36_XI0/XI11/XI10/MM7_d
+ N_XI0/XI11/XI10/NET35_XI0/XI11/XI10/MM7_g N_VSS_XI0/XI11/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM8 N_XI0/XI11/XI10/NET35_XI0/XI11/XI10/MM8_d
+ N_WL<19>_XI0/XI11/XI10/MM8_g N_BLN<5>_XI0/XI11/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI10/MM5 N_XI0/XI11/XI10/NET34_XI0/XI11/XI10/MM5_d
+ N_XI0/XI11/XI10/NET33_XI0/XI11/XI10/MM5_g N_VDD_XI0/XI11/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI10/MM4 N_XI0/XI11/XI10/NET33_XI0/XI11/XI10/MM4_d
+ N_XI0/XI11/XI10/NET34_XI0/XI11/XI10/MM4_g N_VDD_XI0/XI11/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI10/MM10 N_XI0/XI11/XI10/NET35_XI0/XI11/XI10/MM10_d
+ N_XI0/XI11/XI10/NET36_XI0/XI11/XI10/MM10_g N_VDD_XI0/XI11/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI10/MM11 N_XI0/XI11/XI10/NET36_XI0/XI11/XI10/MM11_d
+ N_XI0/XI11/XI10/NET35_XI0/XI11/XI10/MM11_g N_VDD_XI0/XI11/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI11/MM2 N_XI0/XI11/XI11/NET34_XI0/XI11/XI11/MM2_d
+ N_XI0/XI11/XI11/NET33_XI0/XI11/XI11/MM2_g N_VSS_XI0/XI11/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM3 N_XI0/XI11/XI11/NET33_XI0/XI11/XI11/MM3_d
+ N_WL<18>_XI0/XI11/XI11/MM3_g N_BLN<4>_XI0/XI11/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM0 N_XI0/XI11/XI11/NET34_XI0/XI11/XI11/MM0_d
+ N_WL<18>_XI0/XI11/XI11/MM0_g N_BL<4>_XI0/XI11/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM1 N_XI0/XI11/XI11/NET33_XI0/XI11/XI11/MM1_d
+ N_XI0/XI11/XI11/NET34_XI0/XI11/XI11/MM1_g N_VSS_XI0/XI11/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM9 N_XI0/XI11/XI11/NET36_XI0/XI11/XI11/MM9_d
+ N_WL<19>_XI0/XI11/XI11/MM9_g N_BL<4>_XI0/XI11/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM6 N_XI0/XI11/XI11/NET35_XI0/XI11/XI11/MM6_d
+ N_XI0/XI11/XI11/NET36_XI0/XI11/XI11/MM6_g N_VSS_XI0/XI11/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM7 N_XI0/XI11/XI11/NET36_XI0/XI11/XI11/MM7_d
+ N_XI0/XI11/XI11/NET35_XI0/XI11/XI11/MM7_g N_VSS_XI0/XI11/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM8 N_XI0/XI11/XI11/NET35_XI0/XI11/XI11/MM8_d
+ N_WL<19>_XI0/XI11/XI11/MM8_g N_BLN<4>_XI0/XI11/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI11/MM5 N_XI0/XI11/XI11/NET34_XI0/XI11/XI11/MM5_d
+ N_XI0/XI11/XI11/NET33_XI0/XI11/XI11/MM5_g N_VDD_XI0/XI11/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI11/MM4 N_XI0/XI11/XI11/NET33_XI0/XI11/XI11/MM4_d
+ N_XI0/XI11/XI11/NET34_XI0/XI11/XI11/MM4_g N_VDD_XI0/XI11/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI11/MM10 N_XI0/XI11/XI11/NET35_XI0/XI11/XI11/MM10_d
+ N_XI0/XI11/XI11/NET36_XI0/XI11/XI11/MM10_g N_VDD_XI0/XI11/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI11/MM11 N_XI0/XI11/XI11/NET36_XI0/XI11/XI11/MM11_d
+ N_XI0/XI11/XI11/NET35_XI0/XI11/XI11/MM11_g N_VDD_XI0/XI11/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI12/MM2 N_XI0/XI11/XI12/NET34_XI0/XI11/XI12/MM2_d
+ N_XI0/XI11/XI12/NET33_XI0/XI11/XI12/MM2_g N_VSS_XI0/XI11/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM3 N_XI0/XI11/XI12/NET33_XI0/XI11/XI12/MM3_d
+ N_WL<18>_XI0/XI11/XI12/MM3_g N_BLN<3>_XI0/XI11/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM0 N_XI0/XI11/XI12/NET34_XI0/XI11/XI12/MM0_d
+ N_WL<18>_XI0/XI11/XI12/MM0_g N_BL<3>_XI0/XI11/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM1 N_XI0/XI11/XI12/NET33_XI0/XI11/XI12/MM1_d
+ N_XI0/XI11/XI12/NET34_XI0/XI11/XI12/MM1_g N_VSS_XI0/XI11/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM9 N_XI0/XI11/XI12/NET36_XI0/XI11/XI12/MM9_d
+ N_WL<19>_XI0/XI11/XI12/MM9_g N_BL<3>_XI0/XI11/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM6 N_XI0/XI11/XI12/NET35_XI0/XI11/XI12/MM6_d
+ N_XI0/XI11/XI12/NET36_XI0/XI11/XI12/MM6_g N_VSS_XI0/XI11/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM7 N_XI0/XI11/XI12/NET36_XI0/XI11/XI12/MM7_d
+ N_XI0/XI11/XI12/NET35_XI0/XI11/XI12/MM7_g N_VSS_XI0/XI11/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM8 N_XI0/XI11/XI12/NET35_XI0/XI11/XI12/MM8_d
+ N_WL<19>_XI0/XI11/XI12/MM8_g N_BLN<3>_XI0/XI11/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI12/MM5 N_XI0/XI11/XI12/NET34_XI0/XI11/XI12/MM5_d
+ N_XI0/XI11/XI12/NET33_XI0/XI11/XI12/MM5_g N_VDD_XI0/XI11/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI12/MM4 N_XI0/XI11/XI12/NET33_XI0/XI11/XI12/MM4_d
+ N_XI0/XI11/XI12/NET34_XI0/XI11/XI12/MM4_g N_VDD_XI0/XI11/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI12/MM10 N_XI0/XI11/XI12/NET35_XI0/XI11/XI12/MM10_d
+ N_XI0/XI11/XI12/NET36_XI0/XI11/XI12/MM10_g N_VDD_XI0/XI11/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI12/MM11 N_XI0/XI11/XI12/NET36_XI0/XI11/XI12/MM11_d
+ N_XI0/XI11/XI12/NET35_XI0/XI11/XI12/MM11_g N_VDD_XI0/XI11/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI13/MM2 N_XI0/XI11/XI13/NET34_XI0/XI11/XI13/MM2_d
+ N_XI0/XI11/XI13/NET33_XI0/XI11/XI13/MM2_g N_VSS_XI0/XI11/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM3 N_XI0/XI11/XI13/NET33_XI0/XI11/XI13/MM3_d
+ N_WL<18>_XI0/XI11/XI13/MM3_g N_BLN<2>_XI0/XI11/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM0 N_XI0/XI11/XI13/NET34_XI0/XI11/XI13/MM0_d
+ N_WL<18>_XI0/XI11/XI13/MM0_g N_BL<2>_XI0/XI11/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM1 N_XI0/XI11/XI13/NET33_XI0/XI11/XI13/MM1_d
+ N_XI0/XI11/XI13/NET34_XI0/XI11/XI13/MM1_g N_VSS_XI0/XI11/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM9 N_XI0/XI11/XI13/NET36_XI0/XI11/XI13/MM9_d
+ N_WL<19>_XI0/XI11/XI13/MM9_g N_BL<2>_XI0/XI11/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM6 N_XI0/XI11/XI13/NET35_XI0/XI11/XI13/MM6_d
+ N_XI0/XI11/XI13/NET36_XI0/XI11/XI13/MM6_g N_VSS_XI0/XI11/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM7 N_XI0/XI11/XI13/NET36_XI0/XI11/XI13/MM7_d
+ N_XI0/XI11/XI13/NET35_XI0/XI11/XI13/MM7_g N_VSS_XI0/XI11/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM8 N_XI0/XI11/XI13/NET35_XI0/XI11/XI13/MM8_d
+ N_WL<19>_XI0/XI11/XI13/MM8_g N_BLN<2>_XI0/XI11/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI13/MM5 N_XI0/XI11/XI13/NET34_XI0/XI11/XI13/MM5_d
+ N_XI0/XI11/XI13/NET33_XI0/XI11/XI13/MM5_g N_VDD_XI0/XI11/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI13/MM4 N_XI0/XI11/XI13/NET33_XI0/XI11/XI13/MM4_d
+ N_XI0/XI11/XI13/NET34_XI0/XI11/XI13/MM4_g N_VDD_XI0/XI11/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI13/MM10 N_XI0/XI11/XI13/NET35_XI0/XI11/XI13/MM10_d
+ N_XI0/XI11/XI13/NET36_XI0/XI11/XI13/MM10_g N_VDD_XI0/XI11/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI13/MM11 N_XI0/XI11/XI13/NET36_XI0/XI11/XI13/MM11_d
+ N_XI0/XI11/XI13/NET35_XI0/XI11/XI13/MM11_g N_VDD_XI0/XI11/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI14/MM2 N_XI0/XI11/XI14/NET34_XI0/XI11/XI14/MM2_d
+ N_XI0/XI11/XI14/NET33_XI0/XI11/XI14/MM2_g N_VSS_XI0/XI11/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM3 N_XI0/XI11/XI14/NET33_XI0/XI11/XI14/MM3_d
+ N_WL<18>_XI0/XI11/XI14/MM3_g N_BLN<1>_XI0/XI11/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM0 N_XI0/XI11/XI14/NET34_XI0/XI11/XI14/MM0_d
+ N_WL<18>_XI0/XI11/XI14/MM0_g N_BL<1>_XI0/XI11/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM1 N_XI0/XI11/XI14/NET33_XI0/XI11/XI14/MM1_d
+ N_XI0/XI11/XI14/NET34_XI0/XI11/XI14/MM1_g N_VSS_XI0/XI11/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM9 N_XI0/XI11/XI14/NET36_XI0/XI11/XI14/MM9_d
+ N_WL<19>_XI0/XI11/XI14/MM9_g N_BL<1>_XI0/XI11/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM6 N_XI0/XI11/XI14/NET35_XI0/XI11/XI14/MM6_d
+ N_XI0/XI11/XI14/NET36_XI0/XI11/XI14/MM6_g N_VSS_XI0/XI11/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM7 N_XI0/XI11/XI14/NET36_XI0/XI11/XI14/MM7_d
+ N_XI0/XI11/XI14/NET35_XI0/XI11/XI14/MM7_g N_VSS_XI0/XI11/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM8 N_XI0/XI11/XI14/NET35_XI0/XI11/XI14/MM8_d
+ N_WL<19>_XI0/XI11/XI14/MM8_g N_BLN<1>_XI0/XI11/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI14/MM5 N_XI0/XI11/XI14/NET34_XI0/XI11/XI14/MM5_d
+ N_XI0/XI11/XI14/NET33_XI0/XI11/XI14/MM5_g N_VDD_XI0/XI11/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI14/MM4 N_XI0/XI11/XI14/NET33_XI0/XI11/XI14/MM4_d
+ N_XI0/XI11/XI14/NET34_XI0/XI11/XI14/MM4_g N_VDD_XI0/XI11/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI14/MM10 N_XI0/XI11/XI14/NET35_XI0/XI11/XI14/MM10_d
+ N_XI0/XI11/XI14/NET36_XI0/XI11/XI14/MM10_g N_VDD_XI0/XI11/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI14/MM11 N_XI0/XI11/XI14/NET36_XI0/XI11/XI14/MM11_d
+ N_XI0/XI11/XI14/NET35_XI0/XI11/XI14/MM11_g N_VDD_XI0/XI11/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI15/MM2 N_XI0/XI11/XI15/NET34_XI0/XI11/XI15/MM2_d
+ N_XI0/XI11/XI15/NET33_XI0/XI11/XI15/MM2_g N_VSS_XI0/XI11/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM3 N_XI0/XI11/XI15/NET33_XI0/XI11/XI15/MM3_d
+ N_WL<18>_XI0/XI11/XI15/MM3_g N_BLN<0>_XI0/XI11/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM0 N_XI0/XI11/XI15/NET34_XI0/XI11/XI15/MM0_d
+ N_WL<18>_XI0/XI11/XI15/MM0_g N_BL<0>_XI0/XI11/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM1 N_XI0/XI11/XI15/NET33_XI0/XI11/XI15/MM1_d
+ N_XI0/XI11/XI15/NET34_XI0/XI11/XI15/MM1_g N_VSS_XI0/XI11/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM9 N_XI0/XI11/XI15/NET36_XI0/XI11/XI15/MM9_d
+ N_WL<19>_XI0/XI11/XI15/MM9_g N_BL<0>_XI0/XI11/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM6 N_XI0/XI11/XI15/NET35_XI0/XI11/XI15/MM6_d
+ N_XI0/XI11/XI15/NET36_XI0/XI11/XI15/MM6_g N_VSS_XI0/XI11/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM7 N_XI0/XI11/XI15/NET36_XI0/XI11/XI15/MM7_d
+ N_XI0/XI11/XI15/NET35_XI0/XI11/XI15/MM7_g N_VSS_XI0/XI11/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM8 N_XI0/XI11/XI15/NET35_XI0/XI11/XI15/MM8_d
+ N_WL<19>_XI0/XI11/XI15/MM8_g N_BLN<0>_XI0/XI11/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/XI15/MM5 N_XI0/XI11/XI15/NET34_XI0/XI11/XI15/MM5_d
+ N_XI0/XI11/XI15/NET33_XI0/XI11/XI15/MM5_g N_VDD_XI0/XI11/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI15/MM4 N_XI0/XI11/XI15/NET33_XI0/XI11/XI15/MM4_d
+ N_XI0/XI11/XI15/NET34_XI0/XI11/XI15/MM4_g N_VDD_XI0/XI11/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI15/MM10 N_XI0/XI11/XI15/NET35_XI0/XI11/XI15/MM10_d
+ N_XI0/XI11/XI15/NET36_XI0/XI11/XI15/MM10_g N_VDD_XI0/XI11/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/XI15/MM11 N_XI0/XI11/XI15/NET36_XI0/XI11/XI15/MM11_d
+ N_XI0/XI11/XI15/NET35_XI0/XI11/XI15/MM11_g N_VDD_XI0/XI11/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI0/MM2 N_XI0/XI12/XI0/NET34_XI0/XI12/XI0/MM2_d
+ N_XI0/XI12/XI0/NET33_XI0/XI12/XI0/MM2_g N_VSS_XI0/XI12/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM3 N_XI0/XI12/XI0/NET33_XI0/XI12/XI0/MM3_d
+ N_WL<20>_XI0/XI12/XI0/MM3_g N_BLN<15>_XI0/XI12/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM0 N_XI0/XI12/XI0/NET34_XI0/XI12/XI0/MM0_d
+ N_WL<20>_XI0/XI12/XI0/MM0_g N_BL<15>_XI0/XI12/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM1 N_XI0/XI12/XI0/NET33_XI0/XI12/XI0/MM1_d
+ N_XI0/XI12/XI0/NET34_XI0/XI12/XI0/MM1_g N_VSS_XI0/XI12/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM9 N_XI0/XI12/XI0/NET36_XI0/XI12/XI0/MM9_d
+ N_WL<21>_XI0/XI12/XI0/MM9_g N_BL<15>_XI0/XI12/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM6 N_XI0/XI12/XI0/NET35_XI0/XI12/XI0/MM6_d
+ N_XI0/XI12/XI0/NET36_XI0/XI12/XI0/MM6_g N_VSS_XI0/XI12/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM7 N_XI0/XI12/XI0/NET36_XI0/XI12/XI0/MM7_d
+ N_XI0/XI12/XI0/NET35_XI0/XI12/XI0/MM7_g N_VSS_XI0/XI12/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM8 N_XI0/XI12/XI0/NET35_XI0/XI12/XI0/MM8_d
+ N_WL<21>_XI0/XI12/XI0/MM8_g N_BLN<15>_XI0/XI12/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI0/MM5 N_XI0/XI12/XI0/NET34_XI0/XI12/XI0/MM5_d
+ N_XI0/XI12/XI0/NET33_XI0/XI12/XI0/MM5_g N_VDD_XI0/XI12/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI0/MM4 N_XI0/XI12/XI0/NET33_XI0/XI12/XI0/MM4_d
+ N_XI0/XI12/XI0/NET34_XI0/XI12/XI0/MM4_g N_VDD_XI0/XI12/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI0/MM10 N_XI0/XI12/XI0/NET35_XI0/XI12/XI0/MM10_d
+ N_XI0/XI12/XI0/NET36_XI0/XI12/XI0/MM10_g N_VDD_XI0/XI12/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI0/MM11 N_XI0/XI12/XI0/NET36_XI0/XI12/XI0/MM11_d
+ N_XI0/XI12/XI0/NET35_XI0/XI12/XI0/MM11_g N_VDD_XI0/XI12/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI1/MM2 N_XI0/XI12/XI1/NET34_XI0/XI12/XI1/MM2_d
+ N_XI0/XI12/XI1/NET33_XI0/XI12/XI1/MM2_g N_VSS_XI0/XI12/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM3 N_XI0/XI12/XI1/NET33_XI0/XI12/XI1/MM3_d
+ N_WL<20>_XI0/XI12/XI1/MM3_g N_BLN<14>_XI0/XI12/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM0 N_XI0/XI12/XI1/NET34_XI0/XI12/XI1/MM0_d
+ N_WL<20>_XI0/XI12/XI1/MM0_g N_BL<14>_XI0/XI12/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM1 N_XI0/XI12/XI1/NET33_XI0/XI12/XI1/MM1_d
+ N_XI0/XI12/XI1/NET34_XI0/XI12/XI1/MM1_g N_VSS_XI0/XI12/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM9 N_XI0/XI12/XI1/NET36_XI0/XI12/XI1/MM9_d
+ N_WL<21>_XI0/XI12/XI1/MM9_g N_BL<14>_XI0/XI12/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM6 N_XI0/XI12/XI1/NET35_XI0/XI12/XI1/MM6_d
+ N_XI0/XI12/XI1/NET36_XI0/XI12/XI1/MM6_g N_VSS_XI0/XI12/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM7 N_XI0/XI12/XI1/NET36_XI0/XI12/XI1/MM7_d
+ N_XI0/XI12/XI1/NET35_XI0/XI12/XI1/MM7_g N_VSS_XI0/XI12/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM8 N_XI0/XI12/XI1/NET35_XI0/XI12/XI1/MM8_d
+ N_WL<21>_XI0/XI12/XI1/MM8_g N_BLN<14>_XI0/XI12/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI1/MM5 N_XI0/XI12/XI1/NET34_XI0/XI12/XI1/MM5_d
+ N_XI0/XI12/XI1/NET33_XI0/XI12/XI1/MM5_g N_VDD_XI0/XI12/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI1/MM4 N_XI0/XI12/XI1/NET33_XI0/XI12/XI1/MM4_d
+ N_XI0/XI12/XI1/NET34_XI0/XI12/XI1/MM4_g N_VDD_XI0/XI12/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI1/MM10 N_XI0/XI12/XI1/NET35_XI0/XI12/XI1/MM10_d
+ N_XI0/XI12/XI1/NET36_XI0/XI12/XI1/MM10_g N_VDD_XI0/XI12/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI1/MM11 N_XI0/XI12/XI1/NET36_XI0/XI12/XI1/MM11_d
+ N_XI0/XI12/XI1/NET35_XI0/XI12/XI1/MM11_g N_VDD_XI0/XI12/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI2/MM2 N_XI0/XI12/XI2/NET34_XI0/XI12/XI2/MM2_d
+ N_XI0/XI12/XI2/NET33_XI0/XI12/XI2/MM2_g N_VSS_XI0/XI12/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM3 N_XI0/XI12/XI2/NET33_XI0/XI12/XI2/MM3_d
+ N_WL<20>_XI0/XI12/XI2/MM3_g N_BLN<13>_XI0/XI12/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM0 N_XI0/XI12/XI2/NET34_XI0/XI12/XI2/MM0_d
+ N_WL<20>_XI0/XI12/XI2/MM0_g N_BL<13>_XI0/XI12/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM1 N_XI0/XI12/XI2/NET33_XI0/XI12/XI2/MM1_d
+ N_XI0/XI12/XI2/NET34_XI0/XI12/XI2/MM1_g N_VSS_XI0/XI12/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM9 N_XI0/XI12/XI2/NET36_XI0/XI12/XI2/MM9_d
+ N_WL<21>_XI0/XI12/XI2/MM9_g N_BL<13>_XI0/XI12/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM6 N_XI0/XI12/XI2/NET35_XI0/XI12/XI2/MM6_d
+ N_XI0/XI12/XI2/NET36_XI0/XI12/XI2/MM6_g N_VSS_XI0/XI12/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM7 N_XI0/XI12/XI2/NET36_XI0/XI12/XI2/MM7_d
+ N_XI0/XI12/XI2/NET35_XI0/XI12/XI2/MM7_g N_VSS_XI0/XI12/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM8 N_XI0/XI12/XI2/NET35_XI0/XI12/XI2/MM8_d
+ N_WL<21>_XI0/XI12/XI2/MM8_g N_BLN<13>_XI0/XI12/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI2/MM5 N_XI0/XI12/XI2/NET34_XI0/XI12/XI2/MM5_d
+ N_XI0/XI12/XI2/NET33_XI0/XI12/XI2/MM5_g N_VDD_XI0/XI12/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI2/MM4 N_XI0/XI12/XI2/NET33_XI0/XI12/XI2/MM4_d
+ N_XI0/XI12/XI2/NET34_XI0/XI12/XI2/MM4_g N_VDD_XI0/XI12/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI2/MM10 N_XI0/XI12/XI2/NET35_XI0/XI12/XI2/MM10_d
+ N_XI0/XI12/XI2/NET36_XI0/XI12/XI2/MM10_g N_VDD_XI0/XI12/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI2/MM11 N_XI0/XI12/XI2/NET36_XI0/XI12/XI2/MM11_d
+ N_XI0/XI12/XI2/NET35_XI0/XI12/XI2/MM11_g N_VDD_XI0/XI12/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI3/MM2 N_XI0/XI12/XI3/NET34_XI0/XI12/XI3/MM2_d
+ N_XI0/XI12/XI3/NET33_XI0/XI12/XI3/MM2_g N_VSS_XI0/XI12/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM3 N_XI0/XI12/XI3/NET33_XI0/XI12/XI3/MM3_d
+ N_WL<20>_XI0/XI12/XI3/MM3_g N_BLN<12>_XI0/XI12/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM0 N_XI0/XI12/XI3/NET34_XI0/XI12/XI3/MM0_d
+ N_WL<20>_XI0/XI12/XI3/MM0_g N_BL<12>_XI0/XI12/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM1 N_XI0/XI12/XI3/NET33_XI0/XI12/XI3/MM1_d
+ N_XI0/XI12/XI3/NET34_XI0/XI12/XI3/MM1_g N_VSS_XI0/XI12/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM9 N_XI0/XI12/XI3/NET36_XI0/XI12/XI3/MM9_d
+ N_WL<21>_XI0/XI12/XI3/MM9_g N_BL<12>_XI0/XI12/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM6 N_XI0/XI12/XI3/NET35_XI0/XI12/XI3/MM6_d
+ N_XI0/XI12/XI3/NET36_XI0/XI12/XI3/MM6_g N_VSS_XI0/XI12/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM7 N_XI0/XI12/XI3/NET36_XI0/XI12/XI3/MM7_d
+ N_XI0/XI12/XI3/NET35_XI0/XI12/XI3/MM7_g N_VSS_XI0/XI12/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM8 N_XI0/XI12/XI3/NET35_XI0/XI12/XI3/MM8_d
+ N_WL<21>_XI0/XI12/XI3/MM8_g N_BLN<12>_XI0/XI12/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI3/MM5 N_XI0/XI12/XI3/NET34_XI0/XI12/XI3/MM5_d
+ N_XI0/XI12/XI3/NET33_XI0/XI12/XI3/MM5_g N_VDD_XI0/XI12/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI3/MM4 N_XI0/XI12/XI3/NET33_XI0/XI12/XI3/MM4_d
+ N_XI0/XI12/XI3/NET34_XI0/XI12/XI3/MM4_g N_VDD_XI0/XI12/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI3/MM10 N_XI0/XI12/XI3/NET35_XI0/XI12/XI3/MM10_d
+ N_XI0/XI12/XI3/NET36_XI0/XI12/XI3/MM10_g N_VDD_XI0/XI12/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI3/MM11 N_XI0/XI12/XI3/NET36_XI0/XI12/XI3/MM11_d
+ N_XI0/XI12/XI3/NET35_XI0/XI12/XI3/MM11_g N_VDD_XI0/XI12/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI4/MM2 N_XI0/XI12/XI4/NET34_XI0/XI12/XI4/MM2_d
+ N_XI0/XI12/XI4/NET33_XI0/XI12/XI4/MM2_g N_VSS_XI0/XI12/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM3 N_XI0/XI12/XI4/NET33_XI0/XI12/XI4/MM3_d
+ N_WL<20>_XI0/XI12/XI4/MM3_g N_BLN<11>_XI0/XI12/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM0 N_XI0/XI12/XI4/NET34_XI0/XI12/XI4/MM0_d
+ N_WL<20>_XI0/XI12/XI4/MM0_g N_BL<11>_XI0/XI12/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM1 N_XI0/XI12/XI4/NET33_XI0/XI12/XI4/MM1_d
+ N_XI0/XI12/XI4/NET34_XI0/XI12/XI4/MM1_g N_VSS_XI0/XI12/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM9 N_XI0/XI12/XI4/NET36_XI0/XI12/XI4/MM9_d
+ N_WL<21>_XI0/XI12/XI4/MM9_g N_BL<11>_XI0/XI12/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM6 N_XI0/XI12/XI4/NET35_XI0/XI12/XI4/MM6_d
+ N_XI0/XI12/XI4/NET36_XI0/XI12/XI4/MM6_g N_VSS_XI0/XI12/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM7 N_XI0/XI12/XI4/NET36_XI0/XI12/XI4/MM7_d
+ N_XI0/XI12/XI4/NET35_XI0/XI12/XI4/MM7_g N_VSS_XI0/XI12/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM8 N_XI0/XI12/XI4/NET35_XI0/XI12/XI4/MM8_d
+ N_WL<21>_XI0/XI12/XI4/MM8_g N_BLN<11>_XI0/XI12/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI4/MM5 N_XI0/XI12/XI4/NET34_XI0/XI12/XI4/MM5_d
+ N_XI0/XI12/XI4/NET33_XI0/XI12/XI4/MM5_g N_VDD_XI0/XI12/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI4/MM4 N_XI0/XI12/XI4/NET33_XI0/XI12/XI4/MM4_d
+ N_XI0/XI12/XI4/NET34_XI0/XI12/XI4/MM4_g N_VDD_XI0/XI12/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI4/MM10 N_XI0/XI12/XI4/NET35_XI0/XI12/XI4/MM10_d
+ N_XI0/XI12/XI4/NET36_XI0/XI12/XI4/MM10_g N_VDD_XI0/XI12/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI4/MM11 N_XI0/XI12/XI4/NET36_XI0/XI12/XI4/MM11_d
+ N_XI0/XI12/XI4/NET35_XI0/XI12/XI4/MM11_g N_VDD_XI0/XI12/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI5/MM2 N_XI0/XI12/XI5/NET34_XI0/XI12/XI5/MM2_d
+ N_XI0/XI12/XI5/NET33_XI0/XI12/XI5/MM2_g N_VSS_XI0/XI12/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM3 N_XI0/XI12/XI5/NET33_XI0/XI12/XI5/MM3_d
+ N_WL<20>_XI0/XI12/XI5/MM3_g N_BLN<10>_XI0/XI12/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM0 N_XI0/XI12/XI5/NET34_XI0/XI12/XI5/MM0_d
+ N_WL<20>_XI0/XI12/XI5/MM0_g N_BL<10>_XI0/XI12/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM1 N_XI0/XI12/XI5/NET33_XI0/XI12/XI5/MM1_d
+ N_XI0/XI12/XI5/NET34_XI0/XI12/XI5/MM1_g N_VSS_XI0/XI12/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM9 N_XI0/XI12/XI5/NET36_XI0/XI12/XI5/MM9_d
+ N_WL<21>_XI0/XI12/XI5/MM9_g N_BL<10>_XI0/XI12/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM6 N_XI0/XI12/XI5/NET35_XI0/XI12/XI5/MM6_d
+ N_XI0/XI12/XI5/NET36_XI0/XI12/XI5/MM6_g N_VSS_XI0/XI12/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM7 N_XI0/XI12/XI5/NET36_XI0/XI12/XI5/MM7_d
+ N_XI0/XI12/XI5/NET35_XI0/XI12/XI5/MM7_g N_VSS_XI0/XI12/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM8 N_XI0/XI12/XI5/NET35_XI0/XI12/XI5/MM8_d
+ N_WL<21>_XI0/XI12/XI5/MM8_g N_BLN<10>_XI0/XI12/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI5/MM5 N_XI0/XI12/XI5/NET34_XI0/XI12/XI5/MM5_d
+ N_XI0/XI12/XI5/NET33_XI0/XI12/XI5/MM5_g N_VDD_XI0/XI12/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI5/MM4 N_XI0/XI12/XI5/NET33_XI0/XI12/XI5/MM4_d
+ N_XI0/XI12/XI5/NET34_XI0/XI12/XI5/MM4_g N_VDD_XI0/XI12/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI5/MM10 N_XI0/XI12/XI5/NET35_XI0/XI12/XI5/MM10_d
+ N_XI0/XI12/XI5/NET36_XI0/XI12/XI5/MM10_g N_VDD_XI0/XI12/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI5/MM11 N_XI0/XI12/XI5/NET36_XI0/XI12/XI5/MM11_d
+ N_XI0/XI12/XI5/NET35_XI0/XI12/XI5/MM11_g N_VDD_XI0/XI12/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI6/MM2 N_XI0/XI12/XI6/NET34_XI0/XI12/XI6/MM2_d
+ N_XI0/XI12/XI6/NET33_XI0/XI12/XI6/MM2_g N_VSS_XI0/XI12/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM3 N_XI0/XI12/XI6/NET33_XI0/XI12/XI6/MM3_d
+ N_WL<20>_XI0/XI12/XI6/MM3_g N_BLN<9>_XI0/XI12/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM0 N_XI0/XI12/XI6/NET34_XI0/XI12/XI6/MM0_d
+ N_WL<20>_XI0/XI12/XI6/MM0_g N_BL<9>_XI0/XI12/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM1 N_XI0/XI12/XI6/NET33_XI0/XI12/XI6/MM1_d
+ N_XI0/XI12/XI6/NET34_XI0/XI12/XI6/MM1_g N_VSS_XI0/XI12/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM9 N_XI0/XI12/XI6/NET36_XI0/XI12/XI6/MM9_d
+ N_WL<21>_XI0/XI12/XI6/MM9_g N_BL<9>_XI0/XI12/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM6 N_XI0/XI12/XI6/NET35_XI0/XI12/XI6/MM6_d
+ N_XI0/XI12/XI6/NET36_XI0/XI12/XI6/MM6_g N_VSS_XI0/XI12/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM7 N_XI0/XI12/XI6/NET36_XI0/XI12/XI6/MM7_d
+ N_XI0/XI12/XI6/NET35_XI0/XI12/XI6/MM7_g N_VSS_XI0/XI12/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM8 N_XI0/XI12/XI6/NET35_XI0/XI12/XI6/MM8_d
+ N_WL<21>_XI0/XI12/XI6/MM8_g N_BLN<9>_XI0/XI12/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI6/MM5 N_XI0/XI12/XI6/NET34_XI0/XI12/XI6/MM5_d
+ N_XI0/XI12/XI6/NET33_XI0/XI12/XI6/MM5_g N_VDD_XI0/XI12/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI6/MM4 N_XI0/XI12/XI6/NET33_XI0/XI12/XI6/MM4_d
+ N_XI0/XI12/XI6/NET34_XI0/XI12/XI6/MM4_g N_VDD_XI0/XI12/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI6/MM10 N_XI0/XI12/XI6/NET35_XI0/XI12/XI6/MM10_d
+ N_XI0/XI12/XI6/NET36_XI0/XI12/XI6/MM10_g N_VDD_XI0/XI12/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI6/MM11 N_XI0/XI12/XI6/NET36_XI0/XI12/XI6/MM11_d
+ N_XI0/XI12/XI6/NET35_XI0/XI12/XI6/MM11_g N_VDD_XI0/XI12/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI7/MM2 N_XI0/XI12/XI7/NET34_XI0/XI12/XI7/MM2_d
+ N_XI0/XI12/XI7/NET33_XI0/XI12/XI7/MM2_g N_VSS_XI0/XI12/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM3 N_XI0/XI12/XI7/NET33_XI0/XI12/XI7/MM3_d
+ N_WL<20>_XI0/XI12/XI7/MM3_g N_BLN<8>_XI0/XI12/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM0 N_XI0/XI12/XI7/NET34_XI0/XI12/XI7/MM0_d
+ N_WL<20>_XI0/XI12/XI7/MM0_g N_BL<8>_XI0/XI12/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM1 N_XI0/XI12/XI7/NET33_XI0/XI12/XI7/MM1_d
+ N_XI0/XI12/XI7/NET34_XI0/XI12/XI7/MM1_g N_VSS_XI0/XI12/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM9 N_XI0/XI12/XI7/NET36_XI0/XI12/XI7/MM9_d
+ N_WL<21>_XI0/XI12/XI7/MM9_g N_BL<8>_XI0/XI12/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM6 N_XI0/XI12/XI7/NET35_XI0/XI12/XI7/MM6_d
+ N_XI0/XI12/XI7/NET36_XI0/XI12/XI7/MM6_g N_VSS_XI0/XI12/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM7 N_XI0/XI12/XI7/NET36_XI0/XI12/XI7/MM7_d
+ N_XI0/XI12/XI7/NET35_XI0/XI12/XI7/MM7_g N_VSS_XI0/XI12/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM8 N_XI0/XI12/XI7/NET35_XI0/XI12/XI7/MM8_d
+ N_WL<21>_XI0/XI12/XI7/MM8_g N_BLN<8>_XI0/XI12/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI7/MM5 N_XI0/XI12/XI7/NET34_XI0/XI12/XI7/MM5_d
+ N_XI0/XI12/XI7/NET33_XI0/XI12/XI7/MM5_g N_VDD_XI0/XI12/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI7/MM4 N_XI0/XI12/XI7/NET33_XI0/XI12/XI7/MM4_d
+ N_XI0/XI12/XI7/NET34_XI0/XI12/XI7/MM4_g N_VDD_XI0/XI12/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI7/MM10 N_XI0/XI12/XI7/NET35_XI0/XI12/XI7/MM10_d
+ N_XI0/XI12/XI7/NET36_XI0/XI12/XI7/MM10_g N_VDD_XI0/XI12/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI7/MM11 N_XI0/XI12/XI7/NET36_XI0/XI12/XI7/MM11_d
+ N_XI0/XI12/XI7/NET35_XI0/XI12/XI7/MM11_g N_VDD_XI0/XI12/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI8/MM2 N_XI0/XI12/XI8/NET34_XI0/XI12/XI8/MM2_d
+ N_XI0/XI12/XI8/NET33_XI0/XI12/XI8/MM2_g N_VSS_XI0/XI12/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM3 N_XI0/XI12/XI8/NET33_XI0/XI12/XI8/MM3_d
+ N_WL<20>_XI0/XI12/XI8/MM3_g N_BLN<7>_XI0/XI12/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM0 N_XI0/XI12/XI8/NET34_XI0/XI12/XI8/MM0_d
+ N_WL<20>_XI0/XI12/XI8/MM0_g N_BL<7>_XI0/XI12/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM1 N_XI0/XI12/XI8/NET33_XI0/XI12/XI8/MM1_d
+ N_XI0/XI12/XI8/NET34_XI0/XI12/XI8/MM1_g N_VSS_XI0/XI12/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM9 N_XI0/XI12/XI8/NET36_XI0/XI12/XI8/MM9_d
+ N_WL<21>_XI0/XI12/XI8/MM9_g N_BL<7>_XI0/XI12/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM6 N_XI0/XI12/XI8/NET35_XI0/XI12/XI8/MM6_d
+ N_XI0/XI12/XI8/NET36_XI0/XI12/XI8/MM6_g N_VSS_XI0/XI12/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM7 N_XI0/XI12/XI8/NET36_XI0/XI12/XI8/MM7_d
+ N_XI0/XI12/XI8/NET35_XI0/XI12/XI8/MM7_g N_VSS_XI0/XI12/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM8 N_XI0/XI12/XI8/NET35_XI0/XI12/XI8/MM8_d
+ N_WL<21>_XI0/XI12/XI8/MM8_g N_BLN<7>_XI0/XI12/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI8/MM5 N_XI0/XI12/XI8/NET34_XI0/XI12/XI8/MM5_d
+ N_XI0/XI12/XI8/NET33_XI0/XI12/XI8/MM5_g N_VDD_XI0/XI12/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI8/MM4 N_XI0/XI12/XI8/NET33_XI0/XI12/XI8/MM4_d
+ N_XI0/XI12/XI8/NET34_XI0/XI12/XI8/MM4_g N_VDD_XI0/XI12/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI8/MM10 N_XI0/XI12/XI8/NET35_XI0/XI12/XI8/MM10_d
+ N_XI0/XI12/XI8/NET36_XI0/XI12/XI8/MM10_g N_VDD_XI0/XI12/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI8/MM11 N_XI0/XI12/XI8/NET36_XI0/XI12/XI8/MM11_d
+ N_XI0/XI12/XI8/NET35_XI0/XI12/XI8/MM11_g N_VDD_XI0/XI12/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI9/MM2 N_XI0/XI12/XI9/NET34_XI0/XI12/XI9/MM2_d
+ N_XI0/XI12/XI9/NET33_XI0/XI12/XI9/MM2_g N_VSS_XI0/XI12/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM3 N_XI0/XI12/XI9/NET33_XI0/XI12/XI9/MM3_d
+ N_WL<20>_XI0/XI12/XI9/MM3_g N_BLN<6>_XI0/XI12/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM0 N_XI0/XI12/XI9/NET34_XI0/XI12/XI9/MM0_d
+ N_WL<20>_XI0/XI12/XI9/MM0_g N_BL<6>_XI0/XI12/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM1 N_XI0/XI12/XI9/NET33_XI0/XI12/XI9/MM1_d
+ N_XI0/XI12/XI9/NET34_XI0/XI12/XI9/MM1_g N_VSS_XI0/XI12/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM9 N_XI0/XI12/XI9/NET36_XI0/XI12/XI9/MM9_d
+ N_WL<21>_XI0/XI12/XI9/MM9_g N_BL<6>_XI0/XI12/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM6 N_XI0/XI12/XI9/NET35_XI0/XI12/XI9/MM6_d
+ N_XI0/XI12/XI9/NET36_XI0/XI12/XI9/MM6_g N_VSS_XI0/XI12/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM7 N_XI0/XI12/XI9/NET36_XI0/XI12/XI9/MM7_d
+ N_XI0/XI12/XI9/NET35_XI0/XI12/XI9/MM7_g N_VSS_XI0/XI12/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM8 N_XI0/XI12/XI9/NET35_XI0/XI12/XI9/MM8_d
+ N_WL<21>_XI0/XI12/XI9/MM8_g N_BLN<6>_XI0/XI12/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI9/MM5 N_XI0/XI12/XI9/NET34_XI0/XI12/XI9/MM5_d
+ N_XI0/XI12/XI9/NET33_XI0/XI12/XI9/MM5_g N_VDD_XI0/XI12/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI9/MM4 N_XI0/XI12/XI9/NET33_XI0/XI12/XI9/MM4_d
+ N_XI0/XI12/XI9/NET34_XI0/XI12/XI9/MM4_g N_VDD_XI0/XI12/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI9/MM10 N_XI0/XI12/XI9/NET35_XI0/XI12/XI9/MM10_d
+ N_XI0/XI12/XI9/NET36_XI0/XI12/XI9/MM10_g N_VDD_XI0/XI12/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI9/MM11 N_XI0/XI12/XI9/NET36_XI0/XI12/XI9/MM11_d
+ N_XI0/XI12/XI9/NET35_XI0/XI12/XI9/MM11_g N_VDD_XI0/XI12/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI10/MM2 N_XI0/XI12/XI10/NET34_XI0/XI12/XI10/MM2_d
+ N_XI0/XI12/XI10/NET33_XI0/XI12/XI10/MM2_g N_VSS_XI0/XI12/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM3 N_XI0/XI12/XI10/NET33_XI0/XI12/XI10/MM3_d
+ N_WL<20>_XI0/XI12/XI10/MM3_g N_BLN<5>_XI0/XI12/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM0 N_XI0/XI12/XI10/NET34_XI0/XI12/XI10/MM0_d
+ N_WL<20>_XI0/XI12/XI10/MM0_g N_BL<5>_XI0/XI12/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM1 N_XI0/XI12/XI10/NET33_XI0/XI12/XI10/MM1_d
+ N_XI0/XI12/XI10/NET34_XI0/XI12/XI10/MM1_g N_VSS_XI0/XI12/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM9 N_XI0/XI12/XI10/NET36_XI0/XI12/XI10/MM9_d
+ N_WL<21>_XI0/XI12/XI10/MM9_g N_BL<5>_XI0/XI12/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM6 N_XI0/XI12/XI10/NET35_XI0/XI12/XI10/MM6_d
+ N_XI0/XI12/XI10/NET36_XI0/XI12/XI10/MM6_g N_VSS_XI0/XI12/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM7 N_XI0/XI12/XI10/NET36_XI0/XI12/XI10/MM7_d
+ N_XI0/XI12/XI10/NET35_XI0/XI12/XI10/MM7_g N_VSS_XI0/XI12/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM8 N_XI0/XI12/XI10/NET35_XI0/XI12/XI10/MM8_d
+ N_WL<21>_XI0/XI12/XI10/MM8_g N_BLN<5>_XI0/XI12/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI10/MM5 N_XI0/XI12/XI10/NET34_XI0/XI12/XI10/MM5_d
+ N_XI0/XI12/XI10/NET33_XI0/XI12/XI10/MM5_g N_VDD_XI0/XI12/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI10/MM4 N_XI0/XI12/XI10/NET33_XI0/XI12/XI10/MM4_d
+ N_XI0/XI12/XI10/NET34_XI0/XI12/XI10/MM4_g N_VDD_XI0/XI12/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI10/MM10 N_XI0/XI12/XI10/NET35_XI0/XI12/XI10/MM10_d
+ N_XI0/XI12/XI10/NET36_XI0/XI12/XI10/MM10_g N_VDD_XI0/XI12/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI10/MM11 N_XI0/XI12/XI10/NET36_XI0/XI12/XI10/MM11_d
+ N_XI0/XI12/XI10/NET35_XI0/XI12/XI10/MM11_g N_VDD_XI0/XI12/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI11/MM2 N_XI0/XI12/XI11/NET34_XI0/XI12/XI11/MM2_d
+ N_XI0/XI12/XI11/NET33_XI0/XI12/XI11/MM2_g N_VSS_XI0/XI12/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM3 N_XI0/XI12/XI11/NET33_XI0/XI12/XI11/MM3_d
+ N_WL<20>_XI0/XI12/XI11/MM3_g N_BLN<4>_XI0/XI12/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM0 N_XI0/XI12/XI11/NET34_XI0/XI12/XI11/MM0_d
+ N_WL<20>_XI0/XI12/XI11/MM0_g N_BL<4>_XI0/XI12/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM1 N_XI0/XI12/XI11/NET33_XI0/XI12/XI11/MM1_d
+ N_XI0/XI12/XI11/NET34_XI0/XI12/XI11/MM1_g N_VSS_XI0/XI12/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM9 N_XI0/XI12/XI11/NET36_XI0/XI12/XI11/MM9_d
+ N_WL<21>_XI0/XI12/XI11/MM9_g N_BL<4>_XI0/XI12/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM6 N_XI0/XI12/XI11/NET35_XI0/XI12/XI11/MM6_d
+ N_XI0/XI12/XI11/NET36_XI0/XI12/XI11/MM6_g N_VSS_XI0/XI12/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM7 N_XI0/XI12/XI11/NET36_XI0/XI12/XI11/MM7_d
+ N_XI0/XI12/XI11/NET35_XI0/XI12/XI11/MM7_g N_VSS_XI0/XI12/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM8 N_XI0/XI12/XI11/NET35_XI0/XI12/XI11/MM8_d
+ N_WL<21>_XI0/XI12/XI11/MM8_g N_BLN<4>_XI0/XI12/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI11/MM5 N_XI0/XI12/XI11/NET34_XI0/XI12/XI11/MM5_d
+ N_XI0/XI12/XI11/NET33_XI0/XI12/XI11/MM5_g N_VDD_XI0/XI12/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI11/MM4 N_XI0/XI12/XI11/NET33_XI0/XI12/XI11/MM4_d
+ N_XI0/XI12/XI11/NET34_XI0/XI12/XI11/MM4_g N_VDD_XI0/XI12/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI11/MM10 N_XI0/XI12/XI11/NET35_XI0/XI12/XI11/MM10_d
+ N_XI0/XI12/XI11/NET36_XI0/XI12/XI11/MM10_g N_VDD_XI0/XI12/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI11/MM11 N_XI0/XI12/XI11/NET36_XI0/XI12/XI11/MM11_d
+ N_XI0/XI12/XI11/NET35_XI0/XI12/XI11/MM11_g N_VDD_XI0/XI12/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI12/MM2 N_XI0/XI12/XI12/NET34_XI0/XI12/XI12/MM2_d
+ N_XI0/XI12/XI12/NET33_XI0/XI12/XI12/MM2_g N_VSS_XI0/XI12/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM3 N_XI0/XI12/XI12/NET33_XI0/XI12/XI12/MM3_d
+ N_WL<20>_XI0/XI12/XI12/MM3_g N_BLN<3>_XI0/XI12/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM0 N_XI0/XI12/XI12/NET34_XI0/XI12/XI12/MM0_d
+ N_WL<20>_XI0/XI12/XI12/MM0_g N_BL<3>_XI0/XI12/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM1 N_XI0/XI12/XI12/NET33_XI0/XI12/XI12/MM1_d
+ N_XI0/XI12/XI12/NET34_XI0/XI12/XI12/MM1_g N_VSS_XI0/XI12/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM9 N_XI0/XI12/XI12/NET36_XI0/XI12/XI12/MM9_d
+ N_WL<21>_XI0/XI12/XI12/MM9_g N_BL<3>_XI0/XI12/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM6 N_XI0/XI12/XI12/NET35_XI0/XI12/XI12/MM6_d
+ N_XI0/XI12/XI12/NET36_XI0/XI12/XI12/MM6_g N_VSS_XI0/XI12/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM7 N_XI0/XI12/XI12/NET36_XI0/XI12/XI12/MM7_d
+ N_XI0/XI12/XI12/NET35_XI0/XI12/XI12/MM7_g N_VSS_XI0/XI12/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM8 N_XI0/XI12/XI12/NET35_XI0/XI12/XI12/MM8_d
+ N_WL<21>_XI0/XI12/XI12/MM8_g N_BLN<3>_XI0/XI12/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI12/MM5 N_XI0/XI12/XI12/NET34_XI0/XI12/XI12/MM5_d
+ N_XI0/XI12/XI12/NET33_XI0/XI12/XI12/MM5_g N_VDD_XI0/XI12/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI12/MM4 N_XI0/XI12/XI12/NET33_XI0/XI12/XI12/MM4_d
+ N_XI0/XI12/XI12/NET34_XI0/XI12/XI12/MM4_g N_VDD_XI0/XI12/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI12/MM10 N_XI0/XI12/XI12/NET35_XI0/XI12/XI12/MM10_d
+ N_XI0/XI12/XI12/NET36_XI0/XI12/XI12/MM10_g N_VDD_XI0/XI12/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI12/MM11 N_XI0/XI12/XI12/NET36_XI0/XI12/XI12/MM11_d
+ N_XI0/XI12/XI12/NET35_XI0/XI12/XI12/MM11_g N_VDD_XI0/XI12/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI13/MM2 N_XI0/XI12/XI13/NET34_XI0/XI12/XI13/MM2_d
+ N_XI0/XI12/XI13/NET33_XI0/XI12/XI13/MM2_g N_VSS_XI0/XI12/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM3 N_XI0/XI12/XI13/NET33_XI0/XI12/XI13/MM3_d
+ N_WL<20>_XI0/XI12/XI13/MM3_g N_BLN<2>_XI0/XI12/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM0 N_XI0/XI12/XI13/NET34_XI0/XI12/XI13/MM0_d
+ N_WL<20>_XI0/XI12/XI13/MM0_g N_BL<2>_XI0/XI12/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM1 N_XI0/XI12/XI13/NET33_XI0/XI12/XI13/MM1_d
+ N_XI0/XI12/XI13/NET34_XI0/XI12/XI13/MM1_g N_VSS_XI0/XI12/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM9 N_XI0/XI12/XI13/NET36_XI0/XI12/XI13/MM9_d
+ N_WL<21>_XI0/XI12/XI13/MM9_g N_BL<2>_XI0/XI12/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM6 N_XI0/XI12/XI13/NET35_XI0/XI12/XI13/MM6_d
+ N_XI0/XI12/XI13/NET36_XI0/XI12/XI13/MM6_g N_VSS_XI0/XI12/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM7 N_XI0/XI12/XI13/NET36_XI0/XI12/XI13/MM7_d
+ N_XI0/XI12/XI13/NET35_XI0/XI12/XI13/MM7_g N_VSS_XI0/XI12/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM8 N_XI0/XI12/XI13/NET35_XI0/XI12/XI13/MM8_d
+ N_WL<21>_XI0/XI12/XI13/MM8_g N_BLN<2>_XI0/XI12/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI13/MM5 N_XI0/XI12/XI13/NET34_XI0/XI12/XI13/MM5_d
+ N_XI0/XI12/XI13/NET33_XI0/XI12/XI13/MM5_g N_VDD_XI0/XI12/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI13/MM4 N_XI0/XI12/XI13/NET33_XI0/XI12/XI13/MM4_d
+ N_XI0/XI12/XI13/NET34_XI0/XI12/XI13/MM4_g N_VDD_XI0/XI12/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI13/MM10 N_XI0/XI12/XI13/NET35_XI0/XI12/XI13/MM10_d
+ N_XI0/XI12/XI13/NET36_XI0/XI12/XI13/MM10_g N_VDD_XI0/XI12/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI13/MM11 N_XI0/XI12/XI13/NET36_XI0/XI12/XI13/MM11_d
+ N_XI0/XI12/XI13/NET35_XI0/XI12/XI13/MM11_g N_VDD_XI0/XI12/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI14/MM2 N_XI0/XI12/XI14/NET34_XI0/XI12/XI14/MM2_d
+ N_XI0/XI12/XI14/NET33_XI0/XI12/XI14/MM2_g N_VSS_XI0/XI12/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM3 N_XI0/XI12/XI14/NET33_XI0/XI12/XI14/MM3_d
+ N_WL<20>_XI0/XI12/XI14/MM3_g N_BLN<1>_XI0/XI12/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM0 N_XI0/XI12/XI14/NET34_XI0/XI12/XI14/MM0_d
+ N_WL<20>_XI0/XI12/XI14/MM0_g N_BL<1>_XI0/XI12/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM1 N_XI0/XI12/XI14/NET33_XI0/XI12/XI14/MM1_d
+ N_XI0/XI12/XI14/NET34_XI0/XI12/XI14/MM1_g N_VSS_XI0/XI12/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM9 N_XI0/XI12/XI14/NET36_XI0/XI12/XI14/MM9_d
+ N_WL<21>_XI0/XI12/XI14/MM9_g N_BL<1>_XI0/XI12/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM6 N_XI0/XI12/XI14/NET35_XI0/XI12/XI14/MM6_d
+ N_XI0/XI12/XI14/NET36_XI0/XI12/XI14/MM6_g N_VSS_XI0/XI12/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM7 N_XI0/XI12/XI14/NET36_XI0/XI12/XI14/MM7_d
+ N_XI0/XI12/XI14/NET35_XI0/XI12/XI14/MM7_g N_VSS_XI0/XI12/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM8 N_XI0/XI12/XI14/NET35_XI0/XI12/XI14/MM8_d
+ N_WL<21>_XI0/XI12/XI14/MM8_g N_BLN<1>_XI0/XI12/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI14/MM5 N_XI0/XI12/XI14/NET34_XI0/XI12/XI14/MM5_d
+ N_XI0/XI12/XI14/NET33_XI0/XI12/XI14/MM5_g N_VDD_XI0/XI12/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI14/MM4 N_XI0/XI12/XI14/NET33_XI0/XI12/XI14/MM4_d
+ N_XI0/XI12/XI14/NET34_XI0/XI12/XI14/MM4_g N_VDD_XI0/XI12/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI14/MM10 N_XI0/XI12/XI14/NET35_XI0/XI12/XI14/MM10_d
+ N_XI0/XI12/XI14/NET36_XI0/XI12/XI14/MM10_g N_VDD_XI0/XI12/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI14/MM11 N_XI0/XI12/XI14/NET36_XI0/XI12/XI14/MM11_d
+ N_XI0/XI12/XI14/NET35_XI0/XI12/XI14/MM11_g N_VDD_XI0/XI12/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI15/MM2 N_XI0/XI12/XI15/NET34_XI0/XI12/XI15/MM2_d
+ N_XI0/XI12/XI15/NET33_XI0/XI12/XI15/MM2_g N_VSS_XI0/XI12/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM3 N_XI0/XI12/XI15/NET33_XI0/XI12/XI15/MM3_d
+ N_WL<20>_XI0/XI12/XI15/MM3_g N_BLN<0>_XI0/XI12/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM0 N_XI0/XI12/XI15/NET34_XI0/XI12/XI15/MM0_d
+ N_WL<20>_XI0/XI12/XI15/MM0_g N_BL<0>_XI0/XI12/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM1 N_XI0/XI12/XI15/NET33_XI0/XI12/XI15/MM1_d
+ N_XI0/XI12/XI15/NET34_XI0/XI12/XI15/MM1_g N_VSS_XI0/XI12/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM9 N_XI0/XI12/XI15/NET36_XI0/XI12/XI15/MM9_d
+ N_WL<21>_XI0/XI12/XI15/MM9_g N_BL<0>_XI0/XI12/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM6 N_XI0/XI12/XI15/NET35_XI0/XI12/XI15/MM6_d
+ N_XI0/XI12/XI15/NET36_XI0/XI12/XI15/MM6_g N_VSS_XI0/XI12/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM7 N_XI0/XI12/XI15/NET36_XI0/XI12/XI15/MM7_d
+ N_XI0/XI12/XI15/NET35_XI0/XI12/XI15/MM7_g N_VSS_XI0/XI12/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM8 N_XI0/XI12/XI15/NET35_XI0/XI12/XI15/MM8_d
+ N_WL<21>_XI0/XI12/XI15/MM8_g N_BLN<0>_XI0/XI12/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/XI15/MM5 N_XI0/XI12/XI15/NET34_XI0/XI12/XI15/MM5_d
+ N_XI0/XI12/XI15/NET33_XI0/XI12/XI15/MM5_g N_VDD_XI0/XI12/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI15/MM4 N_XI0/XI12/XI15/NET33_XI0/XI12/XI15/MM4_d
+ N_XI0/XI12/XI15/NET34_XI0/XI12/XI15/MM4_g N_VDD_XI0/XI12/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI15/MM10 N_XI0/XI12/XI15/NET35_XI0/XI12/XI15/MM10_d
+ N_XI0/XI12/XI15/NET36_XI0/XI12/XI15/MM10_g N_VDD_XI0/XI12/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/XI15/MM11 N_XI0/XI12/XI15/NET36_XI0/XI12/XI15/MM11_d
+ N_XI0/XI12/XI15/NET35_XI0/XI12/XI15/MM11_g N_VDD_XI0/XI12/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI0/MM2 N_XI0/XI13/XI0/NET34_XI0/XI13/XI0/MM2_d
+ N_XI0/XI13/XI0/NET33_XI0/XI13/XI0/MM2_g N_VSS_XI0/XI13/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM3 N_XI0/XI13/XI0/NET33_XI0/XI13/XI0/MM3_d
+ N_WL<22>_XI0/XI13/XI0/MM3_g N_BLN<15>_XI0/XI13/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM0 N_XI0/XI13/XI0/NET34_XI0/XI13/XI0/MM0_d
+ N_WL<22>_XI0/XI13/XI0/MM0_g N_BL<15>_XI0/XI13/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM1 N_XI0/XI13/XI0/NET33_XI0/XI13/XI0/MM1_d
+ N_XI0/XI13/XI0/NET34_XI0/XI13/XI0/MM1_g N_VSS_XI0/XI13/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM9 N_XI0/XI13/XI0/NET36_XI0/XI13/XI0/MM9_d
+ N_WL<23>_XI0/XI13/XI0/MM9_g N_BL<15>_XI0/XI13/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM6 N_XI0/XI13/XI0/NET35_XI0/XI13/XI0/MM6_d
+ N_XI0/XI13/XI0/NET36_XI0/XI13/XI0/MM6_g N_VSS_XI0/XI13/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM7 N_XI0/XI13/XI0/NET36_XI0/XI13/XI0/MM7_d
+ N_XI0/XI13/XI0/NET35_XI0/XI13/XI0/MM7_g N_VSS_XI0/XI13/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM8 N_XI0/XI13/XI0/NET35_XI0/XI13/XI0/MM8_d
+ N_WL<23>_XI0/XI13/XI0/MM8_g N_BLN<15>_XI0/XI13/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI0/MM5 N_XI0/XI13/XI0/NET34_XI0/XI13/XI0/MM5_d
+ N_XI0/XI13/XI0/NET33_XI0/XI13/XI0/MM5_g N_VDD_XI0/XI13/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI0/MM4 N_XI0/XI13/XI0/NET33_XI0/XI13/XI0/MM4_d
+ N_XI0/XI13/XI0/NET34_XI0/XI13/XI0/MM4_g N_VDD_XI0/XI13/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI0/MM10 N_XI0/XI13/XI0/NET35_XI0/XI13/XI0/MM10_d
+ N_XI0/XI13/XI0/NET36_XI0/XI13/XI0/MM10_g N_VDD_XI0/XI13/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI0/MM11 N_XI0/XI13/XI0/NET36_XI0/XI13/XI0/MM11_d
+ N_XI0/XI13/XI0/NET35_XI0/XI13/XI0/MM11_g N_VDD_XI0/XI13/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI1/MM2 N_XI0/XI13/XI1/NET34_XI0/XI13/XI1/MM2_d
+ N_XI0/XI13/XI1/NET33_XI0/XI13/XI1/MM2_g N_VSS_XI0/XI13/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM3 N_XI0/XI13/XI1/NET33_XI0/XI13/XI1/MM3_d
+ N_WL<22>_XI0/XI13/XI1/MM3_g N_BLN<14>_XI0/XI13/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM0 N_XI0/XI13/XI1/NET34_XI0/XI13/XI1/MM0_d
+ N_WL<22>_XI0/XI13/XI1/MM0_g N_BL<14>_XI0/XI13/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM1 N_XI0/XI13/XI1/NET33_XI0/XI13/XI1/MM1_d
+ N_XI0/XI13/XI1/NET34_XI0/XI13/XI1/MM1_g N_VSS_XI0/XI13/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM9 N_XI0/XI13/XI1/NET36_XI0/XI13/XI1/MM9_d
+ N_WL<23>_XI0/XI13/XI1/MM9_g N_BL<14>_XI0/XI13/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM6 N_XI0/XI13/XI1/NET35_XI0/XI13/XI1/MM6_d
+ N_XI0/XI13/XI1/NET36_XI0/XI13/XI1/MM6_g N_VSS_XI0/XI13/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM7 N_XI0/XI13/XI1/NET36_XI0/XI13/XI1/MM7_d
+ N_XI0/XI13/XI1/NET35_XI0/XI13/XI1/MM7_g N_VSS_XI0/XI13/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM8 N_XI0/XI13/XI1/NET35_XI0/XI13/XI1/MM8_d
+ N_WL<23>_XI0/XI13/XI1/MM8_g N_BLN<14>_XI0/XI13/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI1/MM5 N_XI0/XI13/XI1/NET34_XI0/XI13/XI1/MM5_d
+ N_XI0/XI13/XI1/NET33_XI0/XI13/XI1/MM5_g N_VDD_XI0/XI13/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI1/MM4 N_XI0/XI13/XI1/NET33_XI0/XI13/XI1/MM4_d
+ N_XI0/XI13/XI1/NET34_XI0/XI13/XI1/MM4_g N_VDD_XI0/XI13/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI1/MM10 N_XI0/XI13/XI1/NET35_XI0/XI13/XI1/MM10_d
+ N_XI0/XI13/XI1/NET36_XI0/XI13/XI1/MM10_g N_VDD_XI0/XI13/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI1/MM11 N_XI0/XI13/XI1/NET36_XI0/XI13/XI1/MM11_d
+ N_XI0/XI13/XI1/NET35_XI0/XI13/XI1/MM11_g N_VDD_XI0/XI13/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI2/MM2 N_XI0/XI13/XI2/NET34_XI0/XI13/XI2/MM2_d
+ N_XI0/XI13/XI2/NET33_XI0/XI13/XI2/MM2_g N_VSS_XI0/XI13/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM3 N_XI0/XI13/XI2/NET33_XI0/XI13/XI2/MM3_d
+ N_WL<22>_XI0/XI13/XI2/MM3_g N_BLN<13>_XI0/XI13/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM0 N_XI0/XI13/XI2/NET34_XI0/XI13/XI2/MM0_d
+ N_WL<22>_XI0/XI13/XI2/MM0_g N_BL<13>_XI0/XI13/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM1 N_XI0/XI13/XI2/NET33_XI0/XI13/XI2/MM1_d
+ N_XI0/XI13/XI2/NET34_XI0/XI13/XI2/MM1_g N_VSS_XI0/XI13/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM9 N_XI0/XI13/XI2/NET36_XI0/XI13/XI2/MM9_d
+ N_WL<23>_XI0/XI13/XI2/MM9_g N_BL<13>_XI0/XI13/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM6 N_XI0/XI13/XI2/NET35_XI0/XI13/XI2/MM6_d
+ N_XI0/XI13/XI2/NET36_XI0/XI13/XI2/MM6_g N_VSS_XI0/XI13/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM7 N_XI0/XI13/XI2/NET36_XI0/XI13/XI2/MM7_d
+ N_XI0/XI13/XI2/NET35_XI0/XI13/XI2/MM7_g N_VSS_XI0/XI13/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM8 N_XI0/XI13/XI2/NET35_XI0/XI13/XI2/MM8_d
+ N_WL<23>_XI0/XI13/XI2/MM8_g N_BLN<13>_XI0/XI13/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI2/MM5 N_XI0/XI13/XI2/NET34_XI0/XI13/XI2/MM5_d
+ N_XI0/XI13/XI2/NET33_XI0/XI13/XI2/MM5_g N_VDD_XI0/XI13/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI2/MM4 N_XI0/XI13/XI2/NET33_XI0/XI13/XI2/MM4_d
+ N_XI0/XI13/XI2/NET34_XI0/XI13/XI2/MM4_g N_VDD_XI0/XI13/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI2/MM10 N_XI0/XI13/XI2/NET35_XI0/XI13/XI2/MM10_d
+ N_XI0/XI13/XI2/NET36_XI0/XI13/XI2/MM10_g N_VDD_XI0/XI13/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI2/MM11 N_XI0/XI13/XI2/NET36_XI0/XI13/XI2/MM11_d
+ N_XI0/XI13/XI2/NET35_XI0/XI13/XI2/MM11_g N_VDD_XI0/XI13/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI3/MM2 N_XI0/XI13/XI3/NET34_XI0/XI13/XI3/MM2_d
+ N_XI0/XI13/XI3/NET33_XI0/XI13/XI3/MM2_g N_VSS_XI0/XI13/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM3 N_XI0/XI13/XI3/NET33_XI0/XI13/XI3/MM3_d
+ N_WL<22>_XI0/XI13/XI3/MM3_g N_BLN<12>_XI0/XI13/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM0 N_XI0/XI13/XI3/NET34_XI0/XI13/XI3/MM0_d
+ N_WL<22>_XI0/XI13/XI3/MM0_g N_BL<12>_XI0/XI13/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM1 N_XI0/XI13/XI3/NET33_XI0/XI13/XI3/MM1_d
+ N_XI0/XI13/XI3/NET34_XI0/XI13/XI3/MM1_g N_VSS_XI0/XI13/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM9 N_XI0/XI13/XI3/NET36_XI0/XI13/XI3/MM9_d
+ N_WL<23>_XI0/XI13/XI3/MM9_g N_BL<12>_XI0/XI13/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM6 N_XI0/XI13/XI3/NET35_XI0/XI13/XI3/MM6_d
+ N_XI0/XI13/XI3/NET36_XI0/XI13/XI3/MM6_g N_VSS_XI0/XI13/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM7 N_XI0/XI13/XI3/NET36_XI0/XI13/XI3/MM7_d
+ N_XI0/XI13/XI3/NET35_XI0/XI13/XI3/MM7_g N_VSS_XI0/XI13/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM8 N_XI0/XI13/XI3/NET35_XI0/XI13/XI3/MM8_d
+ N_WL<23>_XI0/XI13/XI3/MM8_g N_BLN<12>_XI0/XI13/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI3/MM5 N_XI0/XI13/XI3/NET34_XI0/XI13/XI3/MM5_d
+ N_XI0/XI13/XI3/NET33_XI0/XI13/XI3/MM5_g N_VDD_XI0/XI13/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI3/MM4 N_XI0/XI13/XI3/NET33_XI0/XI13/XI3/MM4_d
+ N_XI0/XI13/XI3/NET34_XI0/XI13/XI3/MM4_g N_VDD_XI0/XI13/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI3/MM10 N_XI0/XI13/XI3/NET35_XI0/XI13/XI3/MM10_d
+ N_XI0/XI13/XI3/NET36_XI0/XI13/XI3/MM10_g N_VDD_XI0/XI13/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI3/MM11 N_XI0/XI13/XI3/NET36_XI0/XI13/XI3/MM11_d
+ N_XI0/XI13/XI3/NET35_XI0/XI13/XI3/MM11_g N_VDD_XI0/XI13/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI4/MM2 N_XI0/XI13/XI4/NET34_XI0/XI13/XI4/MM2_d
+ N_XI0/XI13/XI4/NET33_XI0/XI13/XI4/MM2_g N_VSS_XI0/XI13/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM3 N_XI0/XI13/XI4/NET33_XI0/XI13/XI4/MM3_d
+ N_WL<22>_XI0/XI13/XI4/MM3_g N_BLN<11>_XI0/XI13/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM0 N_XI0/XI13/XI4/NET34_XI0/XI13/XI4/MM0_d
+ N_WL<22>_XI0/XI13/XI4/MM0_g N_BL<11>_XI0/XI13/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM1 N_XI0/XI13/XI4/NET33_XI0/XI13/XI4/MM1_d
+ N_XI0/XI13/XI4/NET34_XI0/XI13/XI4/MM1_g N_VSS_XI0/XI13/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM9 N_XI0/XI13/XI4/NET36_XI0/XI13/XI4/MM9_d
+ N_WL<23>_XI0/XI13/XI4/MM9_g N_BL<11>_XI0/XI13/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM6 N_XI0/XI13/XI4/NET35_XI0/XI13/XI4/MM6_d
+ N_XI0/XI13/XI4/NET36_XI0/XI13/XI4/MM6_g N_VSS_XI0/XI13/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM7 N_XI0/XI13/XI4/NET36_XI0/XI13/XI4/MM7_d
+ N_XI0/XI13/XI4/NET35_XI0/XI13/XI4/MM7_g N_VSS_XI0/XI13/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM8 N_XI0/XI13/XI4/NET35_XI0/XI13/XI4/MM8_d
+ N_WL<23>_XI0/XI13/XI4/MM8_g N_BLN<11>_XI0/XI13/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI4/MM5 N_XI0/XI13/XI4/NET34_XI0/XI13/XI4/MM5_d
+ N_XI0/XI13/XI4/NET33_XI0/XI13/XI4/MM5_g N_VDD_XI0/XI13/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI4/MM4 N_XI0/XI13/XI4/NET33_XI0/XI13/XI4/MM4_d
+ N_XI0/XI13/XI4/NET34_XI0/XI13/XI4/MM4_g N_VDD_XI0/XI13/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI4/MM10 N_XI0/XI13/XI4/NET35_XI0/XI13/XI4/MM10_d
+ N_XI0/XI13/XI4/NET36_XI0/XI13/XI4/MM10_g N_VDD_XI0/XI13/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI4/MM11 N_XI0/XI13/XI4/NET36_XI0/XI13/XI4/MM11_d
+ N_XI0/XI13/XI4/NET35_XI0/XI13/XI4/MM11_g N_VDD_XI0/XI13/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI5/MM2 N_XI0/XI13/XI5/NET34_XI0/XI13/XI5/MM2_d
+ N_XI0/XI13/XI5/NET33_XI0/XI13/XI5/MM2_g N_VSS_XI0/XI13/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM3 N_XI0/XI13/XI5/NET33_XI0/XI13/XI5/MM3_d
+ N_WL<22>_XI0/XI13/XI5/MM3_g N_BLN<10>_XI0/XI13/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM0 N_XI0/XI13/XI5/NET34_XI0/XI13/XI5/MM0_d
+ N_WL<22>_XI0/XI13/XI5/MM0_g N_BL<10>_XI0/XI13/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM1 N_XI0/XI13/XI5/NET33_XI0/XI13/XI5/MM1_d
+ N_XI0/XI13/XI5/NET34_XI0/XI13/XI5/MM1_g N_VSS_XI0/XI13/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM9 N_XI0/XI13/XI5/NET36_XI0/XI13/XI5/MM9_d
+ N_WL<23>_XI0/XI13/XI5/MM9_g N_BL<10>_XI0/XI13/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM6 N_XI0/XI13/XI5/NET35_XI0/XI13/XI5/MM6_d
+ N_XI0/XI13/XI5/NET36_XI0/XI13/XI5/MM6_g N_VSS_XI0/XI13/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM7 N_XI0/XI13/XI5/NET36_XI0/XI13/XI5/MM7_d
+ N_XI0/XI13/XI5/NET35_XI0/XI13/XI5/MM7_g N_VSS_XI0/XI13/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM8 N_XI0/XI13/XI5/NET35_XI0/XI13/XI5/MM8_d
+ N_WL<23>_XI0/XI13/XI5/MM8_g N_BLN<10>_XI0/XI13/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI5/MM5 N_XI0/XI13/XI5/NET34_XI0/XI13/XI5/MM5_d
+ N_XI0/XI13/XI5/NET33_XI0/XI13/XI5/MM5_g N_VDD_XI0/XI13/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI5/MM4 N_XI0/XI13/XI5/NET33_XI0/XI13/XI5/MM4_d
+ N_XI0/XI13/XI5/NET34_XI0/XI13/XI5/MM4_g N_VDD_XI0/XI13/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI5/MM10 N_XI0/XI13/XI5/NET35_XI0/XI13/XI5/MM10_d
+ N_XI0/XI13/XI5/NET36_XI0/XI13/XI5/MM10_g N_VDD_XI0/XI13/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI5/MM11 N_XI0/XI13/XI5/NET36_XI0/XI13/XI5/MM11_d
+ N_XI0/XI13/XI5/NET35_XI0/XI13/XI5/MM11_g N_VDD_XI0/XI13/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI6/MM2 N_XI0/XI13/XI6/NET34_XI0/XI13/XI6/MM2_d
+ N_XI0/XI13/XI6/NET33_XI0/XI13/XI6/MM2_g N_VSS_XI0/XI13/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM3 N_XI0/XI13/XI6/NET33_XI0/XI13/XI6/MM3_d
+ N_WL<22>_XI0/XI13/XI6/MM3_g N_BLN<9>_XI0/XI13/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM0 N_XI0/XI13/XI6/NET34_XI0/XI13/XI6/MM0_d
+ N_WL<22>_XI0/XI13/XI6/MM0_g N_BL<9>_XI0/XI13/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM1 N_XI0/XI13/XI6/NET33_XI0/XI13/XI6/MM1_d
+ N_XI0/XI13/XI6/NET34_XI0/XI13/XI6/MM1_g N_VSS_XI0/XI13/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM9 N_XI0/XI13/XI6/NET36_XI0/XI13/XI6/MM9_d
+ N_WL<23>_XI0/XI13/XI6/MM9_g N_BL<9>_XI0/XI13/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM6 N_XI0/XI13/XI6/NET35_XI0/XI13/XI6/MM6_d
+ N_XI0/XI13/XI6/NET36_XI0/XI13/XI6/MM6_g N_VSS_XI0/XI13/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM7 N_XI0/XI13/XI6/NET36_XI0/XI13/XI6/MM7_d
+ N_XI0/XI13/XI6/NET35_XI0/XI13/XI6/MM7_g N_VSS_XI0/XI13/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM8 N_XI0/XI13/XI6/NET35_XI0/XI13/XI6/MM8_d
+ N_WL<23>_XI0/XI13/XI6/MM8_g N_BLN<9>_XI0/XI13/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI6/MM5 N_XI0/XI13/XI6/NET34_XI0/XI13/XI6/MM5_d
+ N_XI0/XI13/XI6/NET33_XI0/XI13/XI6/MM5_g N_VDD_XI0/XI13/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI6/MM4 N_XI0/XI13/XI6/NET33_XI0/XI13/XI6/MM4_d
+ N_XI0/XI13/XI6/NET34_XI0/XI13/XI6/MM4_g N_VDD_XI0/XI13/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI6/MM10 N_XI0/XI13/XI6/NET35_XI0/XI13/XI6/MM10_d
+ N_XI0/XI13/XI6/NET36_XI0/XI13/XI6/MM10_g N_VDD_XI0/XI13/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI6/MM11 N_XI0/XI13/XI6/NET36_XI0/XI13/XI6/MM11_d
+ N_XI0/XI13/XI6/NET35_XI0/XI13/XI6/MM11_g N_VDD_XI0/XI13/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI7/MM2 N_XI0/XI13/XI7/NET34_XI0/XI13/XI7/MM2_d
+ N_XI0/XI13/XI7/NET33_XI0/XI13/XI7/MM2_g N_VSS_XI0/XI13/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM3 N_XI0/XI13/XI7/NET33_XI0/XI13/XI7/MM3_d
+ N_WL<22>_XI0/XI13/XI7/MM3_g N_BLN<8>_XI0/XI13/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM0 N_XI0/XI13/XI7/NET34_XI0/XI13/XI7/MM0_d
+ N_WL<22>_XI0/XI13/XI7/MM0_g N_BL<8>_XI0/XI13/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM1 N_XI0/XI13/XI7/NET33_XI0/XI13/XI7/MM1_d
+ N_XI0/XI13/XI7/NET34_XI0/XI13/XI7/MM1_g N_VSS_XI0/XI13/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM9 N_XI0/XI13/XI7/NET36_XI0/XI13/XI7/MM9_d
+ N_WL<23>_XI0/XI13/XI7/MM9_g N_BL<8>_XI0/XI13/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM6 N_XI0/XI13/XI7/NET35_XI0/XI13/XI7/MM6_d
+ N_XI0/XI13/XI7/NET36_XI0/XI13/XI7/MM6_g N_VSS_XI0/XI13/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM7 N_XI0/XI13/XI7/NET36_XI0/XI13/XI7/MM7_d
+ N_XI0/XI13/XI7/NET35_XI0/XI13/XI7/MM7_g N_VSS_XI0/XI13/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM8 N_XI0/XI13/XI7/NET35_XI0/XI13/XI7/MM8_d
+ N_WL<23>_XI0/XI13/XI7/MM8_g N_BLN<8>_XI0/XI13/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI7/MM5 N_XI0/XI13/XI7/NET34_XI0/XI13/XI7/MM5_d
+ N_XI0/XI13/XI7/NET33_XI0/XI13/XI7/MM5_g N_VDD_XI0/XI13/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI7/MM4 N_XI0/XI13/XI7/NET33_XI0/XI13/XI7/MM4_d
+ N_XI0/XI13/XI7/NET34_XI0/XI13/XI7/MM4_g N_VDD_XI0/XI13/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI7/MM10 N_XI0/XI13/XI7/NET35_XI0/XI13/XI7/MM10_d
+ N_XI0/XI13/XI7/NET36_XI0/XI13/XI7/MM10_g N_VDD_XI0/XI13/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI7/MM11 N_XI0/XI13/XI7/NET36_XI0/XI13/XI7/MM11_d
+ N_XI0/XI13/XI7/NET35_XI0/XI13/XI7/MM11_g N_VDD_XI0/XI13/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI8/MM2 N_XI0/XI13/XI8/NET34_XI0/XI13/XI8/MM2_d
+ N_XI0/XI13/XI8/NET33_XI0/XI13/XI8/MM2_g N_VSS_XI0/XI13/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM3 N_XI0/XI13/XI8/NET33_XI0/XI13/XI8/MM3_d
+ N_WL<22>_XI0/XI13/XI8/MM3_g N_BLN<7>_XI0/XI13/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM0 N_XI0/XI13/XI8/NET34_XI0/XI13/XI8/MM0_d
+ N_WL<22>_XI0/XI13/XI8/MM0_g N_BL<7>_XI0/XI13/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM1 N_XI0/XI13/XI8/NET33_XI0/XI13/XI8/MM1_d
+ N_XI0/XI13/XI8/NET34_XI0/XI13/XI8/MM1_g N_VSS_XI0/XI13/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM9 N_XI0/XI13/XI8/NET36_XI0/XI13/XI8/MM9_d
+ N_WL<23>_XI0/XI13/XI8/MM9_g N_BL<7>_XI0/XI13/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM6 N_XI0/XI13/XI8/NET35_XI0/XI13/XI8/MM6_d
+ N_XI0/XI13/XI8/NET36_XI0/XI13/XI8/MM6_g N_VSS_XI0/XI13/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM7 N_XI0/XI13/XI8/NET36_XI0/XI13/XI8/MM7_d
+ N_XI0/XI13/XI8/NET35_XI0/XI13/XI8/MM7_g N_VSS_XI0/XI13/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM8 N_XI0/XI13/XI8/NET35_XI0/XI13/XI8/MM8_d
+ N_WL<23>_XI0/XI13/XI8/MM8_g N_BLN<7>_XI0/XI13/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI8/MM5 N_XI0/XI13/XI8/NET34_XI0/XI13/XI8/MM5_d
+ N_XI0/XI13/XI8/NET33_XI0/XI13/XI8/MM5_g N_VDD_XI0/XI13/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI8/MM4 N_XI0/XI13/XI8/NET33_XI0/XI13/XI8/MM4_d
+ N_XI0/XI13/XI8/NET34_XI0/XI13/XI8/MM4_g N_VDD_XI0/XI13/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI8/MM10 N_XI0/XI13/XI8/NET35_XI0/XI13/XI8/MM10_d
+ N_XI0/XI13/XI8/NET36_XI0/XI13/XI8/MM10_g N_VDD_XI0/XI13/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI8/MM11 N_XI0/XI13/XI8/NET36_XI0/XI13/XI8/MM11_d
+ N_XI0/XI13/XI8/NET35_XI0/XI13/XI8/MM11_g N_VDD_XI0/XI13/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI9/MM2 N_XI0/XI13/XI9/NET34_XI0/XI13/XI9/MM2_d
+ N_XI0/XI13/XI9/NET33_XI0/XI13/XI9/MM2_g N_VSS_XI0/XI13/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM3 N_XI0/XI13/XI9/NET33_XI0/XI13/XI9/MM3_d
+ N_WL<22>_XI0/XI13/XI9/MM3_g N_BLN<6>_XI0/XI13/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM0 N_XI0/XI13/XI9/NET34_XI0/XI13/XI9/MM0_d
+ N_WL<22>_XI0/XI13/XI9/MM0_g N_BL<6>_XI0/XI13/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM1 N_XI0/XI13/XI9/NET33_XI0/XI13/XI9/MM1_d
+ N_XI0/XI13/XI9/NET34_XI0/XI13/XI9/MM1_g N_VSS_XI0/XI13/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM9 N_XI0/XI13/XI9/NET36_XI0/XI13/XI9/MM9_d
+ N_WL<23>_XI0/XI13/XI9/MM9_g N_BL<6>_XI0/XI13/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM6 N_XI0/XI13/XI9/NET35_XI0/XI13/XI9/MM6_d
+ N_XI0/XI13/XI9/NET36_XI0/XI13/XI9/MM6_g N_VSS_XI0/XI13/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM7 N_XI0/XI13/XI9/NET36_XI0/XI13/XI9/MM7_d
+ N_XI0/XI13/XI9/NET35_XI0/XI13/XI9/MM7_g N_VSS_XI0/XI13/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM8 N_XI0/XI13/XI9/NET35_XI0/XI13/XI9/MM8_d
+ N_WL<23>_XI0/XI13/XI9/MM8_g N_BLN<6>_XI0/XI13/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI9/MM5 N_XI0/XI13/XI9/NET34_XI0/XI13/XI9/MM5_d
+ N_XI0/XI13/XI9/NET33_XI0/XI13/XI9/MM5_g N_VDD_XI0/XI13/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI9/MM4 N_XI0/XI13/XI9/NET33_XI0/XI13/XI9/MM4_d
+ N_XI0/XI13/XI9/NET34_XI0/XI13/XI9/MM4_g N_VDD_XI0/XI13/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI9/MM10 N_XI0/XI13/XI9/NET35_XI0/XI13/XI9/MM10_d
+ N_XI0/XI13/XI9/NET36_XI0/XI13/XI9/MM10_g N_VDD_XI0/XI13/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI9/MM11 N_XI0/XI13/XI9/NET36_XI0/XI13/XI9/MM11_d
+ N_XI0/XI13/XI9/NET35_XI0/XI13/XI9/MM11_g N_VDD_XI0/XI13/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI10/MM2 N_XI0/XI13/XI10/NET34_XI0/XI13/XI10/MM2_d
+ N_XI0/XI13/XI10/NET33_XI0/XI13/XI10/MM2_g N_VSS_XI0/XI13/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM3 N_XI0/XI13/XI10/NET33_XI0/XI13/XI10/MM3_d
+ N_WL<22>_XI0/XI13/XI10/MM3_g N_BLN<5>_XI0/XI13/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM0 N_XI0/XI13/XI10/NET34_XI0/XI13/XI10/MM0_d
+ N_WL<22>_XI0/XI13/XI10/MM0_g N_BL<5>_XI0/XI13/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM1 N_XI0/XI13/XI10/NET33_XI0/XI13/XI10/MM1_d
+ N_XI0/XI13/XI10/NET34_XI0/XI13/XI10/MM1_g N_VSS_XI0/XI13/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM9 N_XI0/XI13/XI10/NET36_XI0/XI13/XI10/MM9_d
+ N_WL<23>_XI0/XI13/XI10/MM9_g N_BL<5>_XI0/XI13/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM6 N_XI0/XI13/XI10/NET35_XI0/XI13/XI10/MM6_d
+ N_XI0/XI13/XI10/NET36_XI0/XI13/XI10/MM6_g N_VSS_XI0/XI13/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM7 N_XI0/XI13/XI10/NET36_XI0/XI13/XI10/MM7_d
+ N_XI0/XI13/XI10/NET35_XI0/XI13/XI10/MM7_g N_VSS_XI0/XI13/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM8 N_XI0/XI13/XI10/NET35_XI0/XI13/XI10/MM8_d
+ N_WL<23>_XI0/XI13/XI10/MM8_g N_BLN<5>_XI0/XI13/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI10/MM5 N_XI0/XI13/XI10/NET34_XI0/XI13/XI10/MM5_d
+ N_XI0/XI13/XI10/NET33_XI0/XI13/XI10/MM5_g N_VDD_XI0/XI13/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI10/MM4 N_XI0/XI13/XI10/NET33_XI0/XI13/XI10/MM4_d
+ N_XI0/XI13/XI10/NET34_XI0/XI13/XI10/MM4_g N_VDD_XI0/XI13/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI10/MM10 N_XI0/XI13/XI10/NET35_XI0/XI13/XI10/MM10_d
+ N_XI0/XI13/XI10/NET36_XI0/XI13/XI10/MM10_g N_VDD_XI0/XI13/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI10/MM11 N_XI0/XI13/XI10/NET36_XI0/XI13/XI10/MM11_d
+ N_XI0/XI13/XI10/NET35_XI0/XI13/XI10/MM11_g N_VDD_XI0/XI13/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI11/MM2 N_XI0/XI13/XI11/NET34_XI0/XI13/XI11/MM2_d
+ N_XI0/XI13/XI11/NET33_XI0/XI13/XI11/MM2_g N_VSS_XI0/XI13/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM3 N_XI0/XI13/XI11/NET33_XI0/XI13/XI11/MM3_d
+ N_WL<22>_XI0/XI13/XI11/MM3_g N_BLN<4>_XI0/XI13/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM0 N_XI0/XI13/XI11/NET34_XI0/XI13/XI11/MM0_d
+ N_WL<22>_XI0/XI13/XI11/MM0_g N_BL<4>_XI0/XI13/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM1 N_XI0/XI13/XI11/NET33_XI0/XI13/XI11/MM1_d
+ N_XI0/XI13/XI11/NET34_XI0/XI13/XI11/MM1_g N_VSS_XI0/XI13/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM9 N_XI0/XI13/XI11/NET36_XI0/XI13/XI11/MM9_d
+ N_WL<23>_XI0/XI13/XI11/MM9_g N_BL<4>_XI0/XI13/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM6 N_XI0/XI13/XI11/NET35_XI0/XI13/XI11/MM6_d
+ N_XI0/XI13/XI11/NET36_XI0/XI13/XI11/MM6_g N_VSS_XI0/XI13/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM7 N_XI0/XI13/XI11/NET36_XI0/XI13/XI11/MM7_d
+ N_XI0/XI13/XI11/NET35_XI0/XI13/XI11/MM7_g N_VSS_XI0/XI13/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM8 N_XI0/XI13/XI11/NET35_XI0/XI13/XI11/MM8_d
+ N_WL<23>_XI0/XI13/XI11/MM8_g N_BLN<4>_XI0/XI13/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI11/MM5 N_XI0/XI13/XI11/NET34_XI0/XI13/XI11/MM5_d
+ N_XI0/XI13/XI11/NET33_XI0/XI13/XI11/MM5_g N_VDD_XI0/XI13/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI11/MM4 N_XI0/XI13/XI11/NET33_XI0/XI13/XI11/MM4_d
+ N_XI0/XI13/XI11/NET34_XI0/XI13/XI11/MM4_g N_VDD_XI0/XI13/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI11/MM10 N_XI0/XI13/XI11/NET35_XI0/XI13/XI11/MM10_d
+ N_XI0/XI13/XI11/NET36_XI0/XI13/XI11/MM10_g N_VDD_XI0/XI13/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI11/MM11 N_XI0/XI13/XI11/NET36_XI0/XI13/XI11/MM11_d
+ N_XI0/XI13/XI11/NET35_XI0/XI13/XI11/MM11_g N_VDD_XI0/XI13/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI12/MM2 N_XI0/XI13/XI12/NET34_XI0/XI13/XI12/MM2_d
+ N_XI0/XI13/XI12/NET33_XI0/XI13/XI12/MM2_g N_VSS_XI0/XI13/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM3 N_XI0/XI13/XI12/NET33_XI0/XI13/XI12/MM3_d
+ N_WL<22>_XI0/XI13/XI12/MM3_g N_BLN<3>_XI0/XI13/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM0 N_XI0/XI13/XI12/NET34_XI0/XI13/XI12/MM0_d
+ N_WL<22>_XI0/XI13/XI12/MM0_g N_BL<3>_XI0/XI13/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM1 N_XI0/XI13/XI12/NET33_XI0/XI13/XI12/MM1_d
+ N_XI0/XI13/XI12/NET34_XI0/XI13/XI12/MM1_g N_VSS_XI0/XI13/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM9 N_XI0/XI13/XI12/NET36_XI0/XI13/XI12/MM9_d
+ N_WL<23>_XI0/XI13/XI12/MM9_g N_BL<3>_XI0/XI13/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM6 N_XI0/XI13/XI12/NET35_XI0/XI13/XI12/MM6_d
+ N_XI0/XI13/XI12/NET36_XI0/XI13/XI12/MM6_g N_VSS_XI0/XI13/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM7 N_XI0/XI13/XI12/NET36_XI0/XI13/XI12/MM7_d
+ N_XI0/XI13/XI12/NET35_XI0/XI13/XI12/MM7_g N_VSS_XI0/XI13/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM8 N_XI0/XI13/XI12/NET35_XI0/XI13/XI12/MM8_d
+ N_WL<23>_XI0/XI13/XI12/MM8_g N_BLN<3>_XI0/XI13/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI12/MM5 N_XI0/XI13/XI12/NET34_XI0/XI13/XI12/MM5_d
+ N_XI0/XI13/XI12/NET33_XI0/XI13/XI12/MM5_g N_VDD_XI0/XI13/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI12/MM4 N_XI0/XI13/XI12/NET33_XI0/XI13/XI12/MM4_d
+ N_XI0/XI13/XI12/NET34_XI0/XI13/XI12/MM4_g N_VDD_XI0/XI13/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI12/MM10 N_XI0/XI13/XI12/NET35_XI0/XI13/XI12/MM10_d
+ N_XI0/XI13/XI12/NET36_XI0/XI13/XI12/MM10_g N_VDD_XI0/XI13/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI12/MM11 N_XI0/XI13/XI12/NET36_XI0/XI13/XI12/MM11_d
+ N_XI0/XI13/XI12/NET35_XI0/XI13/XI12/MM11_g N_VDD_XI0/XI13/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI13/MM2 N_XI0/XI13/XI13/NET34_XI0/XI13/XI13/MM2_d
+ N_XI0/XI13/XI13/NET33_XI0/XI13/XI13/MM2_g N_VSS_XI0/XI13/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM3 N_XI0/XI13/XI13/NET33_XI0/XI13/XI13/MM3_d
+ N_WL<22>_XI0/XI13/XI13/MM3_g N_BLN<2>_XI0/XI13/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM0 N_XI0/XI13/XI13/NET34_XI0/XI13/XI13/MM0_d
+ N_WL<22>_XI0/XI13/XI13/MM0_g N_BL<2>_XI0/XI13/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM1 N_XI0/XI13/XI13/NET33_XI0/XI13/XI13/MM1_d
+ N_XI0/XI13/XI13/NET34_XI0/XI13/XI13/MM1_g N_VSS_XI0/XI13/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM9 N_XI0/XI13/XI13/NET36_XI0/XI13/XI13/MM9_d
+ N_WL<23>_XI0/XI13/XI13/MM9_g N_BL<2>_XI0/XI13/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM6 N_XI0/XI13/XI13/NET35_XI0/XI13/XI13/MM6_d
+ N_XI0/XI13/XI13/NET36_XI0/XI13/XI13/MM6_g N_VSS_XI0/XI13/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM7 N_XI0/XI13/XI13/NET36_XI0/XI13/XI13/MM7_d
+ N_XI0/XI13/XI13/NET35_XI0/XI13/XI13/MM7_g N_VSS_XI0/XI13/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM8 N_XI0/XI13/XI13/NET35_XI0/XI13/XI13/MM8_d
+ N_WL<23>_XI0/XI13/XI13/MM8_g N_BLN<2>_XI0/XI13/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI13/MM5 N_XI0/XI13/XI13/NET34_XI0/XI13/XI13/MM5_d
+ N_XI0/XI13/XI13/NET33_XI0/XI13/XI13/MM5_g N_VDD_XI0/XI13/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI13/MM4 N_XI0/XI13/XI13/NET33_XI0/XI13/XI13/MM4_d
+ N_XI0/XI13/XI13/NET34_XI0/XI13/XI13/MM4_g N_VDD_XI0/XI13/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI13/MM10 N_XI0/XI13/XI13/NET35_XI0/XI13/XI13/MM10_d
+ N_XI0/XI13/XI13/NET36_XI0/XI13/XI13/MM10_g N_VDD_XI0/XI13/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI13/MM11 N_XI0/XI13/XI13/NET36_XI0/XI13/XI13/MM11_d
+ N_XI0/XI13/XI13/NET35_XI0/XI13/XI13/MM11_g N_VDD_XI0/XI13/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI14/MM2 N_XI0/XI13/XI14/NET34_XI0/XI13/XI14/MM2_d
+ N_XI0/XI13/XI14/NET33_XI0/XI13/XI14/MM2_g N_VSS_XI0/XI13/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM3 N_XI0/XI13/XI14/NET33_XI0/XI13/XI14/MM3_d
+ N_WL<22>_XI0/XI13/XI14/MM3_g N_BLN<1>_XI0/XI13/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM0 N_XI0/XI13/XI14/NET34_XI0/XI13/XI14/MM0_d
+ N_WL<22>_XI0/XI13/XI14/MM0_g N_BL<1>_XI0/XI13/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM1 N_XI0/XI13/XI14/NET33_XI0/XI13/XI14/MM1_d
+ N_XI0/XI13/XI14/NET34_XI0/XI13/XI14/MM1_g N_VSS_XI0/XI13/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM9 N_XI0/XI13/XI14/NET36_XI0/XI13/XI14/MM9_d
+ N_WL<23>_XI0/XI13/XI14/MM9_g N_BL<1>_XI0/XI13/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM6 N_XI0/XI13/XI14/NET35_XI0/XI13/XI14/MM6_d
+ N_XI0/XI13/XI14/NET36_XI0/XI13/XI14/MM6_g N_VSS_XI0/XI13/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM7 N_XI0/XI13/XI14/NET36_XI0/XI13/XI14/MM7_d
+ N_XI0/XI13/XI14/NET35_XI0/XI13/XI14/MM7_g N_VSS_XI0/XI13/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM8 N_XI0/XI13/XI14/NET35_XI0/XI13/XI14/MM8_d
+ N_WL<23>_XI0/XI13/XI14/MM8_g N_BLN<1>_XI0/XI13/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI14/MM5 N_XI0/XI13/XI14/NET34_XI0/XI13/XI14/MM5_d
+ N_XI0/XI13/XI14/NET33_XI0/XI13/XI14/MM5_g N_VDD_XI0/XI13/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI14/MM4 N_XI0/XI13/XI14/NET33_XI0/XI13/XI14/MM4_d
+ N_XI0/XI13/XI14/NET34_XI0/XI13/XI14/MM4_g N_VDD_XI0/XI13/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI14/MM10 N_XI0/XI13/XI14/NET35_XI0/XI13/XI14/MM10_d
+ N_XI0/XI13/XI14/NET36_XI0/XI13/XI14/MM10_g N_VDD_XI0/XI13/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI14/MM11 N_XI0/XI13/XI14/NET36_XI0/XI13/XI14/MM11_d
+ N_XI0/XI13/XI14/NET35_XI0/XI13/XI14/MM11_g N_VDD_XI0/XI13/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI15/MM2 N_XI0/XI13/XI15/NET34_XI0/XI13/XI15/MM2_d
+ N_XI0/XI13/XI15/NET33_XI0/XI13/XI15/MM2_g N_VSS_XI0/XI13/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM3 N_XI0/XI13/XI15/NET33_XI0/XI13/XI15/MM3_d
+ N_WL<22>_XI0/XI13/XI15/MM3_g N_BLN<0>_XI0/XI13/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM0 N_XI0/XI13/XI15/NET34_XI0/XI13/XI15/MM0_d
+ N_WL<22>_XI0/XI13/XI15/MM0_g N_BL<0>_XI0/XI13/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM1 N_XI0/XI13/XI15/NET33_XI0/XI13/XI15/MM1_d
+ N_XI0/XI13/XI15/NET34_XI0/XI13/XI15/MM1_g N_VSS_XI0/XI13/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM9 N_XI0/XI13/XI15/NET36_XI0/XI13/XI15/MM9_d
+ N_WL<23>_XI0/XI13/XI15/MM9_g N_BL<0>_XI0/XI13/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM6 N_XI0/XI13/XI15/NET35_XI0/XI13/XI15/MM6_d
+ N_XI0/XI13/XI15/NET36_XI0/XI13/XI15/MM6_g N_VSS_XI0/XI13/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM7 N_XI0/XI13/XI15/NET36_XI0/XI13/XI15/MM7_d
+ N_XI0/XI13/XI15/NET35_XI0/XI13/XI15/MM7_g N_VSS_XI0/XI13/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM8 N_XI0/XI13/XI15/NET35_XI0/XI13/XI15/MM8_d
+ N_WL<23>_XI0/XI13/XI15/MM8_g N_BLN<0>_XI0/XI13/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/XI15/MM5 N_XI0/XI13/XI15/NET34_XI0/XI13/XI15/MM5_d
+ N_XI0/XI13/XI15/NET33_XI0/XI13/XI15/MM5_g N_VDD_XI0/XI13/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI15/MM4 N_XI0/XI13/XI15/NET33_XI0/XI13/XI15/MM4_d
+ N_XI0/XI13/XI15/NET34_XI0/XI13/XI15/MM4_g N_VDD_XI0/XI13/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI15/MM10 N_XI0/XI13/XI15/NET35_XI0/XI13/XI15/MM10_d
+ N_XI0/XI13/XI15/NET36_XI0/XI13/XI15/MM10_g N_VDD_XI0/XI13/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/XI15/MM11 N_XI0/XI13/XI15/NET36_XI0/XI13/XI15/MM11_d
+ N_XI0/XI13/XI15/NET35_XI0/XI13/XI15/MM11_g N_VDD_XI0/XI13/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI0/MM2 N_XI0/XI14/XI0/NET34_XI0/XI14/XI0/MM2_d
+ N_XI0/XI14/XI0/NET33_XI0/XI14/XI0/MM2_g N_VSS_XI0/XI14/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM3 N_XI0/XI14/XI0/NET33_XI0/XI14/XI0/MM3_d
+ N_WL<24>_XI0/XI14/XI0/MM3_g N_BLN<15>_XI0/XI14/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM0 N_XI0/XI14/XI0/NET34_XI0/XI14/XI0/MM0_d
+ N_WL<24>_XI0/XI14/XI0/MM0_g N_BL<15>_XI0/XI14/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM1 N_XI0/XI14/XI0/NET33_XI0/XI14/XI0/MM1_d
+ N_XI0/XI14/XI0/NET34_XI0/XI14/XI0/MM1_g N_VSS_XI0/XI14/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM9 N_XI0/XI14/XI0/NET36_XI0/XI14/XI0/MM9_d
+ N_WL<25>_XI0/XI14/XI0/MM9_g N_BL<15>_XI0/XI14/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM6 N_XI0/XI14/XI0/NET35_XI0/XI14/XI0/MM6_d
+ N_XI0/XI14/XI0/NET36_XI0/XI14/XI0/MM6_g N_VSS_XI0/XI14/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM7 N_XI0/XI14/XI0/NET36_XI0/XI14/XI0/MM7_d
+ N_XI0/XI14/XI0/NET35_XI0/XI14/XI0/MM7_g N_VSS_XI0/XI14/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM8 N_XI0/XI14/XI0/NET35_XI0/XI14/XI0/MM8_d
+ N_WL<25>_XI0/XI14/XI0/MM8_g N_BLN<15>_XI0/XI14/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI0/MM5 N_XI0/XI14/XI0/NET34_XI0/XI14/XI0/MM5_d
+ N_XI0/XI14/XI0/NET33_XI0/XI14/XI0/MM5_g N_VDD_XI0/XI14/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI0/MM4 N_XI0/XI14/XI0/NET33_XI0/XI14/XI0/MM4_d
+ N_XI0/XI14/XI0/NET34_XI0/XI14/XI0/MM4_g N_VDD_XI0/XI14/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI0/MM10 N_XI0/XI14/XI0/NET35_XI0/XI14/XI0/MM10_d
+ N_XI0/XI14/XI0/NET36_XI0/XI14/XI0/MM10_g N_VDD_XI0/XI14/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI0/MM11 N_XI0/XI14/XI0/NET36_XI0/XI14/XI0/MM11_d
+ N_XI0/XI14/XI0/NET35_XI0/XI14/XI0/MM11_g N_VDD_XI0/XI14/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI1/MM2 N_XI0/XI14/XI1/NET34_XI0/XI14/XI1/MM2_d
+ N_XI0/XI14/XI1/NET33_XI0/XI14/XI1/MM2_g N_VSS_XI0/XI14/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM3 N_XI0/XI14/XI1/NET33_XI0/XI14/XI1/MM3_d
+ N_WL<24>_XI0/XI14/XI1/MM3_g N_BLN<14>_XI0/XI14/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM0 N_XI0/XI14/XI1/NET34_XI0/XI14/XI1/MM0_d
+ N_WL<24>_XI0/XI14/XI1/MM0_g N_BL<14>_XI0/XI14/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM1 N_XI0/XI14/XI1/NET33_XI0/XI14/XI1/MM1_d
+ N_XI0/XI14/XI1/NET34_XI0/XI14/XI1/MM1_g N_VSS_XI0/XI14/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM9 N_XI0/XI14/XI1/NET36_XI0/XI14/XI1/MM9_d
+ N_WL<25>_XI0/XI14/XI1/MM9_g N_BL<14>_XI0/XI14/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM6 N_XI0/XI14/XI1/NET35_XI0/XI14/XI1/MM6_d
+ N_XI0/XI14/XI1/NET36_XI0/XI14/XI1/MM6_g N_VSS_XI0/XI14/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM7 N_XI0/XI14/XI1/NET36_XI0/XI14/XI1/MM7_d
+ N_XI0/XI14/XI1/NET35_XI0/XI14/XI1/MM7_g N_VSS_XI0/XI14/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM8 N_XI0/XI14/XI1/NET35_XI0/XI14/XI1/MM8_d
+ N_WL<25>_XI0/XI14/XI1/MM8_g N_BLN<14>_XI0/XI14/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI1/MM5 N_XI0/XI14/XI1/NET34_XI0/XI14/XI1/MM5_d
+ N_XI0/XI14/XI1/NET33_XI0/XI14/XI1/MM5_g N_VDD_XI0/XI14/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI1/MM4 N_XI0/XI14/XI1/NET33_XI0/XI14/XI1/MM4_d
+ N_XI0/XI14/XI1/NET34_XI0/XI14/XI1/MM4_g N_VDD_XI0/XI14/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI1/MM10 N_XI0/XI14/XI1/NET35_XI0/XI14/XI1/MM10_d
+ N_XI0/XI14/XI1/NET36_XI0/XI14/XI1/MM10_g N_VDD_XI0/XI14/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI1/MM11 N_XI0/XI14/XI1/NET36_XI0/XI14/XI1/MM11_d
+ N_XI0/XI14/XI1/NET35_XI0/XI14/XI1/MM11_g N_VDD_XI0/XI14/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI2/MM2 N_XI0/XI14/XI2/NET34_XI0/XI14/XI2/MM2_d
+ N_XI0/XI14/XI2/NET33_XI0/XI14/XI2/MM2_g N_VSS_XI0/XI14/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM3 N_XI0/XI14/XI2/NET33_XI0/XI14/XI2/MM3_d
+ N_WL<24>_XI0/XI14/XI2/MM3_g N_BLN<13>_XI0/XI14/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM0 N_XI0/XI14/XI2/NET34_XI0/XI14/XI2/MM0_d
+ N_WL<24>_XI0/XI14/XI2/MM0_g N_BL<13>_XI0/XI14/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM1 N_XI0/XI14/XI2/NET33_XI0/XI14/XI2/MM1_d
+ N_XI0/XI14/XI2/NET34_XI0/XI14/XI2/MM1_g N_VSS_XI0/XI14/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM9 N_XI0/XI14/XI2/NET36_XI0/XI14/XI2/MM9_d
+ N_WL<25>_XI0/XI14/XI2/MM9_g N_BL<13>_XI0/XI14/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM6 N_XI0/XI14/XI2/NET35_XI0/XI14/XI2/MM6_d
+ N_XI0/XI14/XI2/NET36_XI0/XI14/XI2/MM6_g N_VSS_XI0/XI14/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM7 N_XI0/XI14/XI2/NET36_XI0/XI14/XI2/MM7_d
+ N_XI0/XI14/XI2/NET35_XI0/XI14/XI2/MM7_g N_VSS_XI0/XI14/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM8 N_XI0/XI14/XI2/NET35_XI0/XI14/XI2/MM8_d
+ N_WL<25>_XI0/XI14/XI2/MM8_g N_BLN<13>_XI0/XI14/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI2/MM5 N_XI0/XI14/XI2/NET34_XI0/XI14/XI2/MM5_d
+ N_XI0/XI14/XI2/NET33_XI0/XI14/XI2/MM5_g N_VDD_XI0/XI14/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI2/MM4 N_XI0/XI14/XI2/NET33_XI0/XI14/XI2/MM4_d
+ N_XI0/XI14/XI2/NET34_XI0/XI14/XI2/MM4_g N_VDD_XI0/XI14/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI2/MM10 N_XI0/XI14/XI2/NET35_XI0/XI14/XI2/MM10_d
+ N_XI0/XI14/XI2/NET36_XI0/XI14/XI2/MM10_g N_VDD_XI0/XI14/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI2/MM11 N_XI0/XI14/XI2/NET36_XI0/XI14/XI2/MM11_d
+ N_XI0/XI14/XI2/NET35_XI0/XI14/XI2/MM11_g N_VDD_XI0/XI14/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI3/MM2 N_XI0/XI14/XI3/NET34_XI0/XI14/XI3/MM2_d
+ N_XI0/XI14/XI3/NET33_XI0/XI14/XI3/MM2_g N_VSS_XI0/XI14/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM3 N_XI0/XI14/XI3/NET33_XI0/XI14/XI3/MM3_d
+ N_WL<24>_XI0/XI14/XI3/MM3_g N_BLN<12>_XI0/XI14/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM0 N_XI0/XI14/XI3/NET34_XI0/XI14/XI3/MM0_d
+ N_WL<24>_XI0/XI14/XI3/MM0_g N_BL<12>_XI0/XI14/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM1 N_XI0/XI14/XI3/NET33_XI0/XI14/XI3/MM1_d
+ N_XI0/XI14/XI3/NET34_XI0/XI14/XI3/MM1_g N_VSS_XI0/XI14/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM9 N_XI0/XI14/XI3/NET36_XI0/XI14/XI3/MM9_d
+ N_WL<25>_XI0/XI14/XI3/MM9_g N_BL<12>_XI0/XI14/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM6 N_XI0/XI14/XI3/NET35_XI0/XI14/XI3/MM6_d
+ N_XI0/XI14/XI3/NET36_XI0/XI14/XI3/MM6_g N_VSS_XI0/XI14/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM7 N_XI0/XI14/XI3/NET36_XI0/XI14/XI3/MM7_d
+ N_XI0/XI14/XI3/NET35_XI0/XI14/XI3/MM7_g N_VSS_XI0/XI14/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM8 N_XI0/XI14/XI3/NET35_XI0/XI14/XI3/MM8_d
+ N_WL<25>_XI0/XI14/XI3/MM8_g N_BLN<12>_XI0/XI14/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI3/MM5 N_XI0/XI14/XI3/NET34_XI0/XI14/XI3/MM5_d
+ N_XI0/XI14/XI3/NET33_XI0/XI14/XI3/MM5_g N_VDD_XI0/XI14/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI3/MM4 N_XI0/XI14/XI3/NET33_XI0/XI14/XI3/MM4_d
+ N_XI0/XI14/XI3/NET34_XI0/XI14/XI3/MM4_g N_VDD_XI0/XI14/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI3/MM10 N_XI0/XI14/XI3/NET35_XI0/XI14/XI3/MM10_d
+ N_XI0/XI14/XI3/NET36_XI0/XI14/XI3/MM10_g N_VDD_XI0/XI14/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI3/MM11 N_XI0/XI14/XI3/NET36_XI0/XI14/XI3/MM11_d
+ N_XI0/XI14/XI3/NET35_XI0/XI14/XI3/MM11_g N_VDD_XI0/XI14/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI4/MM2 N_XI0/XI14/XI4/NET34_XI0/XI14/XI4/MM2_d
+ N_XI0/XI14/XI4/NET33_XI0/XI14/XI4/MM2_g N_VSS_XI0/XI14/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM3 N_XI0/XI14/XI4/NET33_XI0/XI14/XI4/MM3_d
+ N_WL<24>_XI0/XI14/XI4/MM3_g N_BLN<11>_XI0/XI14/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM0 N_XI0/XI14/XI4/NET34_XI0/XI14/XI4/MM0_d
+ N_WL<24>_XI0/XI14/XI4/MM0_g N_BL<11>_XI0/XI14/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM1 N_XI0/XI14/XI4/NET33_XI0/XI14/XI4/MM1_d
+ N_XI0/XI14/XI4/NET34_XI0/XI14/XI4/MM1_g N_VSS_XI0/XI14/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM9 N_XI0/XI14/XI4/NET36_XI0/XI14/XI4/MM9_d
+ N_WL<25>_XI0/XI14/XI4/MM9_g N_BL<11>_XI0/XI14/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM6 N_XI0/XI14/XI4/NET35_XI0/XI14/XI4/MM6_d
+ N_XI0/XI14/XI4/NET36_XI0/XI14/XI4/MM6_g N_VSS_XI0/XI14/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM7 N_XI0/XI14/XI4/NET36_XI0/XI14/XI4/MM7_d
+ N_XI0/XI14/XI4/NET35_XI0/XI14/XI4/MM7_g N_VSS_XI0/XI14/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM8 N_XI0/XI14/XI4/NET35_XI0/XI14/XI4/MM8_d
+ N_WL<25>_XI0/XI14/XI4/MM8_g N_BLN<11>_XI0/XI14/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI4/MM5 N_XI0/XI14/XI4/NET34_XI0/XI14/XI4/MM5_d
+ N_XI0/XI14/XI4/NET33_XI0/XI14/XI4/MM5_g N_VDD_XI0/XI14/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI4/MM4 N_XI0/XI14/XI4/NET33_XI0/XI14/XI4/MM4_d
+ N_XI0/XI14/XI4/NET34_XI0/XI14/XI4/MM4_g N_VDD_XI0/XI14/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI4/MM10 N_XI0/XI14/XI4/NET35_XI0/XI14/XI4/MM10_d
+ N_XI0/XI14/XI4/NET36_XI0/XI14/XI4/MM10_g N_VDD_XI0/XI14/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI4/MM11 N_XI0/XI14/XI4/NET36_XI0/XI14/XI4/MM11_d
+ N_XI0/XI14/XI4/NET35_XI0/XI14/XI4/MM11_g N_VDD_XI0/XI14/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI5/MM2 N_XI0/XI14/XI5/NET34_XI0/XI14/XI5/MM2_d
+ N_XI0/XI14/XI5/NET33_XI0/XI14/XI5/MM2_g N_VSS_XI0/XI14/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM3 N_XI0/XI14/XI5/NET33_XI0/XI14/XI5/MM3_d
+ N_WL<24>_XI0/XI14/XI5/MM3_g N_BLN<10>_XI0/XI14/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM0 N_XI0/XI14/XI5/NET34_XI0/XI14/XI5/MM0_d
+ N_WL<24>_XI0/XI14/XI5/MM0_g N_BL<10>_XI0/XI14/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM1 N_XI0/XI14/XI5/NET33_XI0/XI14/XI5/MM1_d
+ N_XI0/XI14/XI5/NET34_XI0/XI14/XI5/MM1_g N_VSS_XI0/XI14/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM9 N_XI0/XI14/XI5/NET36_XI0/XI14/XI5/MM9_d
+ N_WL<25>_XI0/XI14/XI5/MM9_g N_BL<10>_XI0/XI14/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM6 N_XI0/XI14/XI5/NET35_XI0/XI14/XI5/MM6_d
+ N_XI0/XI14/XI5/NET36_XI0/XI14/XI5/MM6_g N_VSS_XI0/XI14/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM7 N_XI0/XI14/XI5/NET36_XI0/XI14/XI5/MM7_d
+ N_XI0/XI14/XI5/NET35_XI0/XI14/XI5/MM7_g N_VSS_XI0/XI14/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM8 N_XI0/XI14/XI5/NET35_XI0/XI14/XI5/MM8_d
+ N_WL<25>_XI0/XI14/XI5/MM8_g N_BLN<10>_XI0/XI14/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI5/MM5 N_XI0/XI14/XI5/NET34_XI0/XI14/XI5/MM5_d
+ N_XI0/XI14/XI5/NET33_XI0/XI14/XI5/MM5_g N_VDD_XI0/XI14/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI5/MM4 N_XI0/XI14/XI5/NET33_XI0/XI14/XI5/MM4_d
+ N_XI0/XI14/XI5/NET34_XI0/XI14/XI5/MM4_g N_VDD_XI0/XI14/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI5/MM10 N_XI0/XI14/XI5/NET35_XI0/XI14/XI5/MM10_d
+ N_XI0/XI14/XI5/NET36_XI0/XI14/XI5/MM10_g N_VDD_XI0/XI14/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI5/MM11 N_XI0/XI14/XI5/NET36_XI0/XI14/XI5/MM11_d
+ N_XI0/XI14/XI5/NET35_XI0/XI14/XI5/MM11_g N_VDD_XI0/XI14/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI6/MM2 N_XI0/XI14/XI6/NET34_XI0/XI14/XI6/MM2_d
+ N_XI0/XI14/XI6/NET33_XI0/XI14/XI6/MM2_g N_VSS_XI0/XI14/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM3 N_XI0/XI14/XI6/NET33_XI0/XI14/XI6/MM3_d
+ N_WL<24>_XI0/XI14/XI6/MM3_g N_BLN<9>_XI0/XI14/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM0 N_XI0/XI14/XI6/NET34_XI0/XI14/XI6/MM0_d
+ N_WL<24>_XI0/XI14/XI6/MM0_g N_BL<9>_XI0/XI14/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM1 N_XI0/XI14/XI6/NET33_XI0/XI14/XI6/MM1_d
+ N_XI0/XI14/XI6/NET34_XI0/XI14/XI6/MM1_g N_VSS_XI0/XI14/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM9 N_XI0/XI14/XI6/NET36_XI0/XI14/XI6/MM9_d
+ N_WL<25>_XI0/XI14/XI6/MM9_g N_BL<9>_XI0/XI14/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM6 N_XI0/XI14/XI6/NET35_XI0/XI14/XI6/MM6_d
+ N_XI0/XI14/XI6/NET36_XI0/XI14/XI6/MM6_g N_VSS_XI0/XI14/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM7 N_XI0/XI14/XI6/NET36_XI0/XI14/XI6/MM7_d
+ N_XI0/XI14/XI6/NET35_XI0/XI14/XI6/MM7_g N_VSS_XI0/XI14/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM8 N_XI0/XI14/XI6/NET35_XI0/XI14/XI6/MM8_d
+ N_WL<25>_XI0/XI14/XI6/MM8_g N_BLN<9>_XI0/XI14/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI6/MM5 N_XI0/XI14/XI6/NET34_XI0/XI14/XI6/MM5_d
+ N_XI0/XI14/XI6/NET33_XI0/XI14/XI6/MM5_g N_VDD_XI0/XI14/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI6/MM4 N_XI0/XI14/XI6/NET33_XI0/XI14/XI6/MM4_d
+ N_XI0/XI14/XI6/NET34_XI0/XI14/XI6/MM4_g N_VDD_XI0/XI14/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI6/MM10 N_XI0/XI14/XI6/NET35_XI0/XI14/XI6/MM10_d
+ N_XI0/XI14/XI6/NET36_XI0/XI14/XI6/MM10_g N_VDD_XI0/XI14/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI6/MM11 N_XI0/XI14/XI6/NET36_XI0/XI14/XI6/MM11_d
+ N_XI0/XI14/XI6/NET35_XI0/XI14/XI6/MM11_g N_VDD_XI0/XI14/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI7/MM2 N_XI0/XI14/XI7/NET34_XI0/XI14/XI7/MM2_d
+ N_XI0/XI14/XI7/NET33_XI0/XI14/XI7/MM2_g N_VSS_XI0/XI14/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM3 N_XI0/XI14/XI7/NET33_XI0/XI14/XI7/MM3_d
+ N_WL<24>_XI0/XI14/XI7/MM3_g N_BLN<8>_XI0/XI14/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM0 N_XI0/XI14/XI7/NET34_XI0/XI14/XI7/MM0_d
+ N_WL<24>_XI0/XI14/XI7/MM0_g N_BL<8>_XI0/XI14/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM1 N_XI0/XI14/XI7/NET33_XI0/XI14/XI7/MM1_d
+ N_XI0/XI14/XI7/NET34_XI0/XI14/XI7/MM1_g N_VSS_XI0/XI14/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM9 N_XI0/XI14/XI7/NET36_XI0/XI14/XI7/MM9_d
+ N_WL<25>_XI0/XI14/XI7/MM9_g N_BL<8>_XI0/XI14/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM6 N_XI0/XI14/XI7/NET35_XI0/XI14/XI7/MM6_d
+ N_XI0/XI14/XI7/NET36_XI0/XI14/XI7/MM6_g N_VSS_XI0/XI14/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM7 N_XI0/XI14/XI7/NET36_XI0/XI14/XI7/MM7_d
+ N_XI0/XI14/XI7/NET35_XI0/XI14/XI7/MM7_g N_VSS_XI0/XI14/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM8 N_XI0/XI14/XI7/NET35_XI0/XI14/XI7/MM8_d
+ N_WL<25>_XI0/XI14/XI7/MM8_g N_BLN<8>_XI0/XI14/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI7/MM5 N_XI0/XI14/XI7/NET34_XI0/XI14/XI7/MM5_d
+ N_XI0/XI14/XI7/NET33_XI0/XI14/XI7/MM5_g N_VDD_XI0/XI14/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI7/MM4 N_XI0/XI14/XI7/NET33_XI0/XI14/XI7/MM4_d
+ N_XI0/XI14/XI7/NET34_XI0/XI14/XI7/MM4_g N_VDD_XI0/XI14/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI7/MM10 N_XI0/XI14/XI7/NET35_XI0/XI14/XI7/MM10_d
+ N_XI0/XI14/XI7/NET36_XI0/XI14/XI7/MM10_g N_VDD_XI0/XI14/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI7/MM11 N_XI0/XI14/XI7/NET36_XI0/XI14/XI7/MM11_d
+ N_XI0/XI14/XI7/NET35_XI0/XI14/XI7/MM11_g N_VDD_XI0/XI14/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI8/MM2 N_XI0/XI14/XI8/NET34_XI0/XI14/XI8/MM2_d
+ N_XI0/XI14/XI8/NET33_XI0/XI14/XI8/MM2_g N_VSS_XI0/XI14/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM3 N_XI0/XI14/XI8/NET33_XI0/XI14/XI8/MM3_d
+ N_WL<24>_XI0/XI14/XI8/MM3_g N_BLN<7>_XI0/XI14/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM0 N_XI0/XI14/XI8/NET34_XI0/XI14/XI8/MM0_d
+ N_WL<24>_XI0/XI14/XI8/MM0_g N_BL<7>_XI0/XI14/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM1 N_XI0/XI14/XI8/NET33_XI0/XI14/XI8/MM1_d
+ N_XI0/XI14/XI8/NET34_XI0/XI14/XI8/MM1_g N_VSS_XI0/XI14/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM9 N_XI0/XI14/XI8/NET36_XI0/XI14/XI8/MM9_d
+ N_WL<25>_XI0/XI14/XI8/MM9_g N_BL<7>_XI0/XI14/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM6 N_XI0/XI14/XI8/NET35_XI0/XI14/XI8/MM6_d
+ N_XI0/XI14/XI8/NET36_XI0/XI14/XI8/MM6_g N_VSS_XI0/XI14/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM7 N_XI0/XI14/XI8/NET36_XI0/XI14/XI8/MM7_d
+ N_XI0/XI14/XI8/NET35_XI0/XI14/XI8/MM7_g N_VSS_XI0/XI14/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM8 N_XI0/XI14/XI8/NET35_XI0/XI14/XI8/MM8_d
+ N_WL<25>_XI0/XI14/XI8/MM8_g N_BLN<7>_XI0/XI14/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI8/MM5 N_XI0/XI14/XI8/NET34_XI0/XI14/XI8/MM5_d
+ N_XI0/XI14/XI8/NET33_XI0/XI14/XI8/MM5_g N_VDD_XI0/XI14/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI8/MM4 N_XI0/XI14/XI8/NET33_XI0/XI14/XI8/MM4_d
+ N_XI0/XI14/XI8/NET34_XI0/XI14/XI8/MM4_g N_VDD_XI0/XI14/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI8/MM10 N_XI0/XI14/XI8/NET35_XI0/XI14/XI8/MM10_d
+ N_XI0/XI14/XI8/NET36_XI0/XI14/XI8/MM10_g N_VDD_XI0/XI14/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI8/MM11 N_XI0/XI14/XI8/NET36_XI0/XI14/XI8/MM11_d
+ N_XI0/XI14/XI8/NET35_XI0/XI14/XI8/MM11_g N_VDD_XI0/XI14/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI9/MM2 N_XI0/XI14/XI9/NET34_XI0/XI14/XI9/MM2_d
+ N_XI0/XI14/XI9/NET33_XI0/XI14/XI9/MM2_g N_VSS_XI0/XI14/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM3 N_XI0/XI14/XI9/NET33_XI0/XI14/XI9/MM3_d
+ N_WL<24>_XI0/XI14/XI9/MM3_g N_BLN<6>_XI0/XI14/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM0 N_XI0/XI14/XI9/NET34_XI0/XI14/XI9/MM0_d
+ N_WL<24>_XI0/XI14/XI9/MM0_g N_BL<6>_XI0/XI14/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM1 N_XI0/XI14/XI9/NET33_XI0/XI14/XI9/MM1_d
+ N_XI0/XI14/XI9/NET34_XI0/XI14/XI9/MM1_g N_VSS_XI0/XI14/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM9 N_XI0/XI14/XI9/NET36_XI0/XI14/XI9/MM9_d
+ N_WL<25>_XI0/XI14/XI9/MM9_g N_BL<6>_XI0/XI14/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM6 N_XI0/XI14/XI9/NET35_XI0/XI14/XI9/MM6_d
+ N_XI0/XI14/XI9/NET36_XI0/XI14/XI9/MM6_g N_VSS_XI0/XI14/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM7 N_XI0/XI14/XI9/NET36_XI0/XI14/XI9/MM7_d
+ N_XI0/XI14/XI9/NET35_XI0/XI14/XI9/MM7_g N_VSS_XI0/XI14/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM8 N_XI0/XI14/XI9/NET35_XI0/XI14/XI9/MM8_d
+ N_WL<25>_XI0/XI14/XI9/MM8_g N_BLN<6>_XI0/XI14/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI9/MM5 N_XI0/XI14/XI9/NET34_XI0/XI14/XI9/MM5_d
+ N_XI0/XI14/XI9/NET33_XI0/XI14/XI9/MM5_g N_VDD_XI0/XI14/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI9/MM4 N_XI0/XI14/XI9/NET33_XI0/XI14/XI9/MM4_d
+ N_XI0/XI14/XI9/NET34_XI0/XI14/XI9/MM4_g N_VDD_XI0/XI14/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI9/MM10 N_XI0/XI14/XI9/NET35_XI0/XI14/XI9/MM10_d
+ N_XI0/XI14/XI9/NET36_XI0/XI14/XI9/MM10_g N_VDD_XI0/XI14/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI9/MM11 N_XI0/XI14/XI9/NET36_XI0/XI14/XI9/MM11_d
+ N_XI0/XI14/XI9/NET35_XI0/XI14/XI9/MM11_g N_VDD_XI0/XI14/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI10/MM2 N_XI0/XI14/XI10/NET34_XI0/XI14/XI10/MM2_d
+ N_XI0/XI14/XI10/NET33_XI0/XI14/XI10/MM2_g N_VSS_XI0/XI14/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM3 N_XI0/XI14/XI10/NET33_XI0/XI14/XI10/MM3_d
+ N_WL<24>_XI0/XI14/XI10/MM3_g N_BLN<5>_XI0/XI14/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM0 N_XI0/XI14/XI10/NET34_XI0/XI14/XI10/MM0_d
+ N_WL<24>_XI0/XI14/XI10/MM0_g N_BL<5>_XI0/XI14/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM1 N_XI0/XI14/XI10/NET33_XI0/XI14/XI10/MM1_d
+ N_XI0/XI14/XI10/NET34_XI0/XI14/XI10/MM1_g N_VSS_XI0/XI14/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM9 N_XI0/XI14/XI10/NET36_XI0/XI14/XI10/MM9_d
+ N_WL<25>_XI0/XI14/XI10/MM9_g N_BL<5>_XI0/XI14/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM6 N_XI0/XI14/XI10/NET35_XI0/XI14/XI10/MM6_d
+ N_XI0/XI14/XI10/NET36_XI0/XI14/XI10/MM6_g N_VSS_XI0/XI14/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM7 N_XI0/XI14/XI10/NET36_XI0/XI14/XI10/MM7_d
+ N_XI0/XI14/XI10/NET35_XI0/XI14/XI10/MM7_g N_VSS_XI0/XI14/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM8 N_XI0/XI14/XI10/NET35_XI0/XI14/XI10/MM8_d
+ N_WL<25>_XI0/XI14/XI10/MM8_g N_BLN<5>_XI0/XI14/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI10/MM5 N_XI0/XI14/XI10/NET34_XI0/XI14/XI10/MM5_d
+ N_XI0/XI14/XI10/NET33_XI0/XI14/XI10/MM5_g N_VDD_XI0/XI14/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI10/MM4 N_XI0/XI14/XI10/NET33_XI0/XI14/XI10/MM4_d
+ N_XI0/XI14/XI10/NET34_XI0/XI14/XI10/MM4_g N_VDD_XI0/XI14/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI10/MM10 N_XI0/XI14/XI10/NET35_XI0/XI14/XI10/MM10_d
+ N_XI0/XI14/XI10/NET36_XI0/XI14/XI10/MM10_g N_VDD_XI0/XI14/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI10/MM11 N_XI0/XI14/XI10/NET36_XI0/XI14/XI10/MM11_d
+ N_XI0/XI14/XI10/NET35_XI0/XI14/XI10/MM11_g N_VDD_XI0/XI14/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI11/MM2 N_XI0/XI14/XI11/NET34_XI0/XI14/XI11/MM2_d
+ N_XI0/XI14/XI11/NET33_XI0/XI14/XI11/MM2_g N_VSS_XI0/XI14/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM3 N_XI0/XI14/XI11/NET33_XI0/XI14/XI11/MM3_d
+ N_WL<24>_XI0/XI14/XI11/MM3_g N_BLN<4>_XI0/XI14/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM0 N_XI0/XI14/XI11/NET34_XI0/XI14/XI11/MM0_d
+ N_WL<24>_XI0/XI14/XI11/MM0_g N_BL<4>_XI0/XI14/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM1 N_XI0/XI14/XI11/NET33_XI0/XI14/XI11/MM1_d
+ N_XI0/XI14/XI11/NET34_XI0/XI14/XI11/MM1_g N_VSS_XI0/XI14/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM9 N_XI0/XI14/XI11/NET36_XI0/XI14/XI11/MM9_d
+ N_WL<25>_XI0/XI14/XI11/MM9_g N_BL<4>_XI0/XI14/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM6 N_XI0/XI14/XI11/NET35_XI0/XI14/XI11/MM6_d
+ N_XI0/XI14/XI11/NET36_XI0/XI14/XI11/MM6_g N_VSS_XI0/XI14/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM7 N_XI0/XI14/XI11/NET36_XI0/XI14/XI11/MM7_d
+ N_XI0/XI14/XI11/NET35_XI0/XI14/XI11/MM7_g N_VSS_XI0/XI14/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM8 N_XI0/XI14/XI11/NET35_XI0/XI14/XI11/MM8_d
+ N_WL<25>_XI0/XI14/XI11/MM8_g N_BLN<4>_XI0/XI14/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI11/MM5 N_XI0/XI14/XI11/NET34_XI0/XI14/XI11/MM5_d
+ N_XI0/XI14/XI11/NET33_XI0/XI14/XI11/MM5_g N_VDD_XI0/XI14/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI11/MM4 N_XI0/XI14/XI11/NET33_XI0/XI14/XI11/MM4_d
+ N_XI0/XI14/XI11/NET34_XI0/XI14/XI11/MM4_g N_VDD_XI0/XI14/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI11/MM10 N_XI0/XI14/XI11/NET35_XI0/XI14/XI11/MM10_d
+ N_XI0/XI14/XI11/NET36_XI0/XI14/XI11/MM10_g N_VDD_XI0/XI14/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI11/MM11 N_XI0/XI14/XI11/NET36_XI0/XI14/XI11/MM11_d
+ N_XI0/XI14/XI11/NET35_XI0/XI14/XI11/MM11_g N_VDD_XI0/XI14/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI12/MM2 N_XI0/XI14/XI12/NET34_XI0/XI14/XI12/MM2_d
+ N_XI0/XI14/XI12/NET33_XI0/XI14/XI12/MM2_g N_VSS_XI0/XI14/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM3 N_XI0/XI14/XI12/NET33_XI0/XI14/XI12/MM3_d
+ N_WL<24>_XI0/XI14/XI12/MM3_g N_BLN<3>_XI0/XI14/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM0 N_XI0/XI14/XI12/NET34_XI0/XI14/XI12/MM0_d
+ N_WL<24>_XI0/XI14/XI12/MM0_g N_BL<3>_XI0/XI14/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM1 N_XI0/XI14/XI12/NET33_XI0/XI14/XI12/MM1_d
+ N_XI0/XI14/XI12/NET34_XI0/XI14/XI12/MM1_g N_VSS_XI0/XI14/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM9 N_XI0/XI14/XI12/NET36_XI0/XI14/XI12/MM9_d
+ N_WL<25>_XI0/XI14/XI12/MM9_g N_BL<3>_XI0/XI14/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM6 N_XI0/XI14/XI12/NET35_XI0/XI14/XI12/MM6_d
+ N_XI0/XI14/XI12/NET36_XI0/XI14/XI12/MM6_g N_VSS_XI0/XI14/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM7 N_XI0/XI14/XI12/NET36_XI0/XI14/XI12/MM7_d
+ N_XI0/XI14/XI12/NET35_XI0/XI14/XI12/MM7_g N_VSS_XI0/XI14/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM8 N_XI0/XI14/XI12/NET35_XI0/XI14/XI12/MM8_d
+ N_WL<25>_XI0/XI14/XI12/MM8_g N_BLN<3>_XI0/XI14/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI12/MM5 N_XI0/XI14/XI12/NET34_XI0/XI14/XI12/MM5_d
+ N_XI0/XI14/XI12/NET33_XI0/XI14/XI12/MM5_g N_VDD_XI0/XI14/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI12/MM4 N_XI0/XI14/XI12/NET33_XI0/XI14/XI12/MM4_d
+ N_XI0/XI14/XI12/NET34_XI0/XI14/XI12/MM4_g N_VDD_XI0/XI14/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI12/MM10 N_XI0/XI14/XI12/NET35_XI0/XI14/XI12/MM10_d
+ N_XI0/XI14/XI12/NET36_XI0/XI14/XI12/MM10_g N_VDD_XI0/XI14/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI12/MM11 N_XI0/XI14/XI12/NET36_XI0/XI14/XI12/MM11_d
+ N_XI0/XI14/XI12/NET35_XI0/XI14/XI12/MM11_g N_VDD_XI0/XI14/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI13/MM2 N_XI0/XI14/XI13/NET34_XI0/XI14/XI13/MM2_d
+ N_XI0/XI14/XI13/NET33_XI0/XI14/XI13/MM2_g N_VSS_XI0/XI14/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM3 N_XI0/XI14/XI13/NET33_XI0/XI14/XI13/MM3_d
+ N_WL<24>_XI0/XI14/XI13/MM3_g N_BLN<2>_XI0/XI14/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM0 N_XI0/XI14/XI13/NET34_XI0/XI14/XI13/MM0_d
+ N_WL<24>_XI0/XI14/XI13/MM0_g N_BL<2>_XI0/XI14/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM1 N_XI0/XI14/XI13/NET33_XI0/XI14/XI13/MM1_d
+ N_XI0/XI14/XI13/NET34_XI0/XI14/XI13/MM1_g N_VSS_XI0/XI14/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM9 N_XI0/XI14/XI13/NET36_XI0/XI14/XI13/MM9_d
+ N_WL<25>_XI0/XI14/XI13/MM9_g N_BL<2>_XI0/XI14/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM6 N_XI0/XI14/XI13/NET35_XI0/XI14/XI13/MM6_d
+ N_XI0/XI14/XI13/NET36_XI0/XI14/XI13/MM6_g N_VSS_XI0/XI14/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM7 N_XI0/XI14/XI13/NET36_XI0/XI14/XI13/MM7_d
+ N_XI0/XI14/XI13/NET35_XI0/XI14/XI13/MM7_g N_VSS_XI0/XI14/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM8 N_XI0/XI14/XI13/NET35_XI0/XI14/XI13/MM8_d
+ N_WL<25>_XI0/XI14/XI13/MM8_g N_BLN<2>_XI0/XI14/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI13/MM5 N_XI0/XI14/XI13/NET34_XI0/XI14/XI13/MM5_d
+ N_XI0/XI14/XI13/NET33_XI0/XI14/XI13/MM5_g N_VDD_XI0/XI14/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI13/MM4 N_XI0/XI14/XI13/NET33_XI0/XI14/XI13/MM4_d
+ N_XI0/XI14/XI13/NET34_XI0/XI14/XI13/MM4_g N_VDD_XI0/XI14/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI13/MM10 N_XI0/XI14/XI13/NET35_XI0/XI14/XI13/MM10_d
+ N_XI0/XI14/XI13/NET36_XI0/XI14/XI13/MM10_g N_VDD_XI0/XI14/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI13/MM11 N_XI0/XI14/XI13/NET36_XI0/XI14/XI13/MM11_d
+ N_XI0/XI14/XI13/NET35_XI0/XI14/XI13/MM11_g N_VDD_XI0/XI14/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI14/MM2 N_XI0/XI14/XI14/NET34_XI0/XI14/XI14/MM2_d
+ N_XI0/XI14/XI14/NET33_XI0/XI14/XI14/MM2_g N_VSS_XI0/XI14/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM3 N_XI0/XI14/XI14/NET33_XI0/XI14/XI14/MM3_d
+ N_WL<24>_XI0/XI14/XI14/MM3_g N_BLN<1>_XI0/XI14/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM0 N_XI0/XI14/XI14/NET34_XI0/XI14/XI14/MM0_d
+ N_WL<24>_XI0/XI14/XI14/MM0_g N_BL<1>_XI0/XI14/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM1 N_XI0/XI14/XI14/NET33_XI0/XI14/XI14/MM1_d
+ N_XI0/XI14/XI14/NET34_XI0/XI14/XI14/MM1_g N_VSS_XI0/XI14/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM9 N_XI0/XI14/XI14/NET36_XI0/XI14/XI14/MM9_d
+ N_WL<25>_XI0/XI14/XI14/MM9_g N_BL<1>_XI0/XI14/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM6 N_XI0/XI14/XI14/NET35_XI0/XI14/XI14/MM6_d
+ N_XI0/XI14/XI14/NET36_XI0/XI14/XI14/MM6_g N_VSS_XI0/XI14/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM7 N_XI0/XI14/XI14/NET36_XI0/XI14/XI14/MM7_d
+ N_XI0/XI14/XI14/NET35_XI0/XI14/XI14/MM7_g N_VSS_XI0/XI14/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM8 N_XI0/XI14/XI14/NET35_XI0/XI14/XI14/MM8_d
+ N_WL<25>_XI0/XI14/XI14/MM8_g N_BLN<1>_XI0/XI14/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI14/MM5 N_XI0/XI14/XI14/NET34_XI0/XI14/XI14/MM5_d
+ N_XI0/XI14/XI14/NET33_XI0/XI14/XI14/MM5_g N_VDD_XI0/XI14/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI14/MM4 N_XI0/XI14/XI14/NET33_XI0/XI14/XI14/MM4_d
+ N_XI0/XI14/XI14/NET34_XI0/XI14/XI14/MM4_g N_VDD_XI0/XI14/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI14/MM10 N_XI0/XI14/XI14/NET35_XI0/XI14/XI14/MM10_d
+ N_XI0/XI14/XI14/NET36_XI0/XI14/XI14/MM10_g N_VDD_XI0/XI14/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI14/MM11 N_XI0/XI14/XI14/NET36_XI0/XI14/XI14/MM11_d
+ N_XI0/XI14/XI14/NET35_XI0/XI14/XI14/MM11_g N_VDD_XI0/XI14/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI15/MM2 N_XI0/XI14/XI15/NET34_XI0/XI14/XI15/MM2_d
+ N_XI0/XI14/XI15/NET33_XI0/XI14/XI15/MM2_g N_VSS_XI0/XI14/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM3 N_XI0/XI14/XI15/NET33_XI0/XI14/XI15/MM3_d
+ N_WL<24>_XI0/XI14/XI15/MM3_g N_BLN<0>_XI0/XI14/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM0 N_XI0/XI14/XI15/NET34_XI0/XI14/XI15/MM0_d
+ N_WL<24>_XI0/XI14/XI15/MM0_g N_BL<0>_XI0/XI14/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM1 N_XI0/XI14/XI15/NET33_XI0/XI14/XI15/MM1_d
+ N_XI0/XI14/XI15/NET34_XI0/XI14/XI15/MM1_g N_VSS_XI0/XI14/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM9 N_XI0/XI14/XI15/NET36_XI0/XI14/XI15/MM9_d
+ N_WL<25>_XI0/XI14/XI15/MM9_g N_BL<0>_XI0/XI14/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM6 N_XI0/XI14/XI15/NET35_XI0/XI14/XI15/MM6_d
+ N_XI0/XI14/XI15/NET36_XI0/XI14/XI15/MM6_g N_VSS_XI0/XI14/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM7 N_XI0/XI14/XI15/NET36_XI0/XI14/XI15/MM7_d
+ N_XI0/XI14/XI15/NET35_XI0/XI14/XI15/MM7_g N_VSS_XI0/XI14/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM8 N_XI0/XI14/XI15/NET35_XI0/XI14/XI15/MM8_d
+ N_WL<25>_XI0/XI14/XI15/MM8_g N_BLN<0>_XI0/XI14/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/XI15/MM5 N_XI0/XI14/XI15/NET34_XI0/XI14/XI15/MM5_d
+ N_XI0/XI14/XI15/NET33_XI0/XI14/XI15/MM5_g N_VDD_XI0/XI14/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI15/MM4 N_XI0/XI14/XI15/NET33_XI0/XI14/XI15/MM4_d
+ N_XI0/XI14/XI15/NET34_XI0/XI14/XI15/MM4_g N_VDD_XI0/XI14/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI15/MM10 N_XI0/XI14/XI15/NET35_XI0/XI14/XI15/MM10_d
+ N_XI0/XI14/XI15/NET36_XI0/XI14/XI15/MM10_g N_VDD_XI0/XI14/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/XI15/MM11 N_XI0/XI14/XI15/NET36_XI0/XI14/XI15/MM11_d
+ N_XI0/XI14/XI15/NET35_XI0/XI14/XI15/MM11_g N_VDD_XI0/XI14/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI0/MM2 N_XI0/XI15/XI0/NET34_XI0/XI15/XI0/MM2_d
+ N_XI0/XI15/XI0/NET33_XI0/XI15/XI0/MM2_g N_VSS_XI0/XI15/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM3 N_XI0/XI15/XI0/NET33_XI0/XI15/XI0/MM3_d
+ N_WL<26>_XI0/XI15/XI0/MM3_g N_BLN<15>_XI0/XI15/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM0 N_XI0/XI15/XI0/NET34_XI0/XI15/XI0/MM0_d
+ N_WL<26>_XI0/XI15/XI0/MM0_g N_BL<15>_XI0/XI15/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM1 N_XI0/XI15/XI0/NET33_XI0/XI15/XI0/MM1_d
+ N_XI0/XI15/XI0/NET34_XI0/XI15/XI0/MM1_g N_VSS_XI0/XI15/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM9 N_XI0/XI15/XI0/NET36_XI0/XI15/XI0/MM9_d
+ N_WL<27>_XI0/XI15/XI0/MM9_g N_BL<15>_XI0/XI15/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM6 N_XI0/XI15/XI0/NET35_XI0/XI15/XI0/MM6_d
+ N_XI0/XI15/XI0/NET36_XI0/XI15/XI0/MM6_g N_VSS_XI0/XI15/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM7 N_XI0/XI15/XI0/NET36_XI0/XI15/XI0/MM7_d
+ N_XI0/XI15/XI0/NET35_XI0/XI15/XI0/MM7_g N_VSS_XI0/XI15/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM8 N_XI0/XI15/XI0/NET35_XI0/XI15/XI0/MM8_d
+ N_WL<27>_XI0/XI15/XI0/MM8_g N_BLN<15>_XI0/XI15/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI0/MM5 N_XI0/XI15/XI0/NET34_XI0/XI15/XI0/MM5_d
+ N_XI0/XI15/XI0/NET33_XI0/XI15/XI0/MM5_g N_VDD_XI0/XI15/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI0/MM4 N_XI0/XI15/XI0/NET33_XI0/XI15/XI0/MM4_d
+ N_XI0/XI15/XI0/NET34_XI0/XI15/XI0/MM4_g N_VDD_XI0/XI15/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI0/MM10 N_XI0/XI15/XI0/NET35_XI0/XI15/XI0/MM10_d
+ N_XI0/XI15/XI0/NET36_XI0/XI15/XI0/MM10_g N_VDD_XI0/XI15/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI0/MM11 N_XI0/XI15/XI0/NET36_XI0/XI15/XI0/MM11_d
+ N_XI0/XI15/XI0/NET35_XI0/XI15/XI0/MM11_g N_VDD_XI0/XI15/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI1/MM2 N_XI0/XI15/XI1/NET34_XI0/XI15/XI1/MM2_d
+ N_XI0/XI15/XI1/NET33_XI0/XI15/XI1/MM2_g N_VSS_XI0/XI15/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM3 N_XI0/XI15/XI1/NET33_XI0/XI15/XI1/MM3_d
+ N_WL<26>_XI0/XI15/XI1/MM3_g N_BLN<14>_XI0/XI15/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM0 N_XI0/XI15/XI1/NET34_XI0/XI15/XI1/MM0_d
+ N_WL<26>_XI0/XI15/XI1/MM0_g N_BL<14>_XI0/XI15/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM1 N_XI0/XI15/XI1/NET33_XI0/XI15/XI1/MM1_d
+ N_XI0/XI15/XI1/NET34_XI0/XI15/XI1/MM1_g N_VSS_XI0/XI15/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM9 N_XI0/XI15/XI1/NET36_XI0/XI15/XI1/MM9_d
+ N_WL<27>_XI0/XI15/XI1/MM9_g N_BL<14>_XI0/XI15/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM6 N_XI0/XI15/XI1/NET35_XI0/XI15/XI1/MM6_d
+ N_XI0/XI15/XI1/NET36_XI0/XI15/XI1/MM6_g N_VSS_XI0/XI15/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM7 N_XI0/XI15/XI1/NET36_XI0/XI15/XI1/MM7_d
+ N_XI0/XI15/XI1/NET35_XI0/XI15/XI1/MM7_g N_VSS_XI0/XI15/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM8 N_XI0/XI15/XI1/NET35_XI0/XI15/XI1/MM8_d
+ N_WL<27>_XI0/XI15/XI1/MM8_g N_BLN<14>_XI0/XI15/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI1/MM5 N_XI0/XI15/XI1/NET34_XI0/XI15/XI1/MM5_d
+ N_XI0/XI15/XI1/NET33_XI0/XI15/XI1/MM5_g N_VDD_XI0/XI15/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI1/MM4 N_XI0/XI15/XI1/NET33_XI0/XI15/XI1/MM4_d
+ N_XI0/XI15/XI1/NET34_XI0/XI15/XI1/MM4_g N_VDD_XI0/XI15/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI1/MM10 N_XI0/XI15/XI1/NET35_XI0/XI15/XI1/MM10_d
+ N_XI0/XI15/XI1/NET36_XI0/XI15/XI1/MM10_g N_VDD_XI0/XI15/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI1/MM11 N_XI0/XI15/XI1/NET36_XI0/XI15/XI1/MM11_d
+ N_XI0/XI15/XI1/NET35_XI0/XI15/XI1/MM11_g N_VDD_XI0/XI15/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI2/MM2 N_XI0/XI15/XI2/NET34_XI0/XI15/XI2/MM2_d
+ N_XI0/XI15/XI2/NET33_XI0/XI15/XI2/MM2_g N_VSS_XI0/XI15/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM3 N_XI0/XI15/XI2/NET33_XI0/XI15/XI2/MM3_d
+ N_WL<26>_XI0/XI15/XI2/MM3_g N_BLN<13>_XI0/XI15/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM0 N_XI0/XI15/XI2/NET34_XI0/XI15/XI2/MM0_d
+ N_WL<26>_XI0/XI15/XI2/MM0_g N_BL<13>_XI0/XI15/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM1 N_XI0/XI15/XI2/NET33_XI0/XI15/XI2/MM1_d
+ N_XI0/XI15/XI2/NET34_XI0/XI15/XI2/MM1_g N_VSS_XI0/XI15/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM9 N_XI0/XI15/XI2/NET36_XI0/XI15/XI2/MM9_d
+ N_WL<27>_XI0/XI15/XI2/MM9_g N_BL<13>_XI0/XI15/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM6 N_XI0/XI15/XI2/NET35_XI0/XI15/XI2/MM6_d
+ N_XI0/XI15/XI2/NET36_XI0/XI15/XI2/MM6_g N_VSS_XI0/XI15/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM7 N_XI0/XI15/XI2/NET36_XI0/XI15/XI2/MM7_d
+ N_XI0/XI15/XI2/NET35_XI0/XI15/XI2/MM7_g N_VSS_XI0/XI15/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM8 N_XI0/XI15/XI2/NET35_XI0/XI15/XI2/MM8_d
+ N_WL<27>_XI0/XI15/XI2/MM8_g N_BLN<13>_XI0/XI15/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI2/MM5 N_XI0/XI15/XI2/NET34_XI0/XI15/XI2/MM5_d
+ N_XI0/XI15/XI2/NET33_XI0/XI15/XI2/MM5_g N_VDD_XI0/XI15/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI2/MM4 N_XI0/XI15/XI2/NET33_XI0/XI15/XI2/MM4_d
+ N_XI0/XI15/XI2/NET34_XI0/XI15/XI2/MM4_g N_VDD_XI0/XI15/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI2/MM10 N_XI0/XI15/XI2/NET35_XI0/XI15/XI2/MM10_d
+ N_XI0/XI15/XI2/NET36_XI0/XI15/XI2/MM10_g N_VDD_XI0/XI15/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI2/MM11 N_XI0/XI15/XI2/NET36_XI0/XI15/XI2/MM11_d
+ N_XI0/XI15/XI2/NET35_XI0/XI15/XI2/MM11_g N_VDD_XI0/XI15/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI3/MM2 N_XI0/XI15/XI3/NET34_XI0/XI15/XI3/MM2_d
+ N_XI0/XI15/XI3/NET33_XI0/XI15/XI3/MM2_g N_VSS_XI0/XI15/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM3 N_XI0/XI15/XI3/NET33_XI0/XI15/XI3/MM3_d
+ N_WL<26>_XI0/XI15/XI3/MM3_g N_BLN<12>_XI0/XI15/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM0 N_XI0/XI15/XI3/NET34_XI0/XI15/XI3/MM0_d
+ N_WL<26>_XI0/XI15/XI3/MM0_g N_BL<12>_XI0/XI15/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM1 N_XI0/XI15/XI3/NET33_XI0/XI15/XI3/MM1_d
+ N_XI0/XI15/XI3/NET34_XI0/XI15/XI3/MM1_g N_VSS_XI0/XI15/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM9 N_XI0/XI15/XI3/NET36_XI0/XI15/XI3/MM9_d
+ N_WL<27>_XI0/XI15/XI3/MM9_g N_BL<12>_XI0/XI15/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM6 N_XI0/XI15/XI3/NET35_XI0/XI15/XI3/MM6_d
+ N_XI0/XI15/XI3/NET36_XI0/XI15/XI3/MM6_g N_VSS_XI0/XI15/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM7 N_XI0/XI15/XI3/NET36_XI0/XI15/XI3/MM7_d
+ N_XI0/XI15/XI3/NET35_XI0/XI15/XI3/MM7_g N_VSS_XI0/XI15/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM8 N_XI0/XI15/XI3/NET35_XI0/XI15/XI3/MM8_d
+ N_WL<27>_XI0/XI15/XI3/MM8_g N_BLN<12>_XI0/XI15/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI3/MM5 N_XI0/XI15/XI3/NET34_XI0/XI15/XI3/MM5_d
+ N_XI0/XI15/XI3/NET33_XI0/XI15/XI3/MM5_g N_VDD_XI0/XI15/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI3/MM4 N_XI0/XI15/XI3/NET33_XI0/XI15/XI3/MM4_d
+ N_XI0/XI15/XI3/NET34_XI0/XI15/XI3/MM4_g N_VDD_XI0/XI15/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI3/MM10 N_XI0/XI15/XI3/NET35_XI0/XI15/XI3/MM10_d
+ N_XI0/XI15/XI3/NET36_XI0/XI15/XI3/MM10_g N_VDD_XI0/XI15/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI3/MM11 N_XI0/XI15/XI3/NET36_XI0/XI15/XI3/MM11_d
+ N_XI0/XI15/XI3/NET35_XI0/XI15/XI3/MM11_g N_VDD_XI0/XI15/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI4/MM2 N_XI0/XI15/XI4/NET34_XI0/XI15/XI4/MM2_d
+ N_XI0/XI15/XI4/NET33_XI0/XI15/XI4/MM2_g N_VSS_XI0/XI15/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM3 N_XI0/XI15/XI4/NET33_XI0/XI15/XI4/MM3_d
+ N_WL<26>_XI0/XI15/XI4/MM3_g N_BLN<11>_XI0/XI15/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM0 N_XI0/XI15/XI4/NET34_XI0/XI15/XI4/MM0_d
+ N_WL<26>_XI0/XI15/XI4/MM0_g N_BL<11>_XI0/XI15/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM1 N_XI0/XI15/XI4/NET33_XI0/XI15/XI4/MM1_d
+ N_XI0/XI15/XI4/NET34_XI0/XI15/XI4/MM1_g N_VSS_XI0/XI15/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM9 N_XI0/XI15/XI4/NET36_XI0/XI15/XI4/MM9_d
+ N_WL<27>_XI0/XI15/XI4/MM9_g N_BL<11>_XI0/XI15/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM6 N_XI0/XI15/XI4/NET35_XI0/XI15/XI4/MM6_d
+ N_XI0/XI15/XI4/NET36_XI0/XI15/XI4/MM6_g N_VSS_XI0/XI15/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM7 N_XI0/XI15/XI4/NET36_XI0/XI15/XI4/MM7_d
+ N_XI0/XI15/XI4/NET35_XI0/XI15/XI4/MM7_g N_VSS_XI0/XI15/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM8 N_XI0/XI15/XI4/NET35_XI0/XI15/XI4/MM8_d
+ N_WL<27>_XI0/XI15/XI4/MM8_g N_BLN<11>_XI0/XI15/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI4/MM5 N_XI0/XI15/XI4/NET34_XI0/XI15/XI4/MM5_d
+ N_XI0/XI15/XI4/NET33_XI0/XI15/XI4/MM5_g N_VDD_XI0/XI15/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI4/MM4 N_XI0/XI15/XI4/NET33_XI0/XI15/XI4/MM4_d
+ N_XI0/XI15/XI4/NET34_XI0/XI15/XI4/MM4_g N_VDD_XI0/XI15/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI4/MM10 N_XI0/XI15/XI4/NET35_XI0/XI15/XI4/MM10_d
+ N_XI0/XI15/XI4/NET36_XI0/XI15/XI4/MM10_g N_VDD_XI0/XI15/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI4/MM11 N_XI0/XI15/XI4/NET36_XI0/XI15/XI4/MM11_d
+ N_XI0/XI15/XI4/NET35_XI0/XI15/XI4/MM11_g N_VDD_XI0/XI15/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI5/MM2 N_XI0/XI15/XI5/NET34_XI0/XI15/XI5/MM2_d
+ N_XI0/XI15/XI5/NET33_XI0/XI15/XI5/MM2_g N_VSS_XI0/XI15/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM3 N_XI0/XI15/XI5/NET33_XI0/XI15/XI5/MM3_d
+ N_WL<26>_XI0/XI15/XI5/MM3_g N_BLN<10>_XI0/XI15/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM0 N_XI0/XI15/XI5/NET34_XI0/XI15/XI5/MM0_d
+ N_WL<26>_XI0/XI15/XI5/MM0_g N_BL<10>_XI0/XI15/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM1 N_XI0/XI15/XI5/NET33_XI0/XI15/XI5/MM1_d
+ N_XI0/XI15/XI5/NET34_XI0/XI15/XI5/MM1_g N_VSS_XI0/XI15/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM9 N_XI0/XI15/XI5/NET36_XI0/XI15/XI5/MM9_d
+ N_WL<27>_XI0/XI15/XI5/MM9_g N_BL<10>_XI0/XI15/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM6 N_XI0/XI15/XI5/NET35_XI0/XI15/XI5/MM6_d
+ N_XI0/XI15/XI5/NET36_XI0/XI15/XI5/MM6_g N_VSS_XI0/XI15/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM7 N_XI0/XI15/XI5/NET36_XI0/XI15/XI5/MM7_d
+ N_XI0/XI15/XI5/NET35_XI0/XI15/XI5/MM7_g N_VSS_XI0/XI15/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM8 N_XI0/XI15/XI5/NET35_XI0/XI15/XI5/MM8_d
+ N_WL<27>_XI0/XI15/XI5/MM8_g N_BLN<10>_XI0/XI15/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI5/MM5 N_XI0/XI15/XI5/NET34_XI0/XI15/XI5/MM5_d
+ N_XI0/XI15/XI5/NET33_XI0/XI15/XI5/MM5_g N_VDD_XI0/XI15/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI5/MM4 N_XI0/XI15/XI5/NET33_XI0/XI15/XI5/MM4_d
+ N_XI0/XI15/XI5/NET34_XI0/XI15/XI5/MM4_g N_VDD_XI0/XI15/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI5/MM10 N_XI0/XI15/XI5/NET35_XI0/XI15/XI5/MM10_d
+ N_XI0/XI15/XI5/NET36_XI0/XI15/XI5/MM10_g N_VDD_XI0/XI15/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI5/MM11 N_XI0/XI15/XI5/NET36_XI0/XI15/XI5/MM11_d
+ N_XI0/XI15/XI5/NET35_XI0/XI15/XI5/MM11_g N_VDD_XI0/XI15/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI6/MM2 N_XI0/XI15/XI6/NET34_XI0/XI15/XI6/MM2_d
+ N_XI0/XI15/XI6/NET33_XI0/XI15/XI6/MM2_g N_VSS_XI0/XI15/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM3 N_XI0/XI15/XI6/NET33_XI0/XI15/XI6/MM3_d
+ N_WL<26>_XI0/XI15/XI6/MM3_g N_BLN<9>_XI0/XI15/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM0 N_XI0/XI15/XI6/NET34_XI0/XI15/XI6/MM0_d
+ N_WL<26>_XI0/XI15/XI6/MM0_g N_BL<9>_XI0/XI15/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM1 N_XI0/XI15/XI6/NET33_XI0/XI15/XI6/MM1_d
+ N_XI0/XI15/XI6/NET34_XI0/XI15/XI6/MM1_g N_VSS_XI0/XI15/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM9 N_XI0/XI15/XI6/NET36_XI0/XI15/XI6/MM9_d
+ N_WL<27>_XI0/XI15/XI6/MM9_g N_BL<9>_XI0/XI15/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM6 N_XI0/XI15/XI6/NET35_XI0/XI15/XI6/MM6_d
+ N_XI0/XI15/XI6/NET36_XI0/XI15/XI6/MM6_g N_VSS_XI0/XI15/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM7 N_XI0/XI15/XI6/NET36_XI0/XI15/XI6/MM7_d
+ N_XI0/XI15/XI6/NET35_XI0/XI15/XI6/MM7_g N_VSS_XI0/XI15/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM8 N_XI0/XI15/XI6/NET35_XI0/XI15/XI6/MM8_d
+ N_WL<27>_XI0/XI15/XI6/MM8_g N_BLN<9>_XI0/XI15/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI6/MM5 N_XI0/XI15/XI6/NET34_XI0/XI15/XI6/MM5_d
+ N_XI0/XI15/XI6/NET33_XI0/XI15/XI6/MM5_g N_VDD_XI0/XI15/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI6/MM4 N_XI0/XI15/XI6/NET33_XI0/XI15/XI6/MM4_d
+ N_XI0/XI15/XI6/NET34_XI0/XI15/XI6/MM4_g N_VDD_XI0/XI15/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI6/MM10 N_XI0/XI15/XI6/NET35_XI0/XI15/XI6/MM10_d
+ N_XI0/XI15/XI6/NET36_XI0/XI15/XI6/MM10_g N_VDD_XI0/XI15/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI6/MM11 N_XI0/XI15/XI6/NET36_XI0/XI15/XI6/MM11_d
+ N_XI0/XI15/XI6/NET35_XI0/XI15/XI6/MM11_g N_VDD_XI0/XI15/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI7/MM2 N_XI0/XI15/XI7/NET34_XI0/XI15/XI7/MM2_d
+ N_XI0/XI15/XI7/NET33_XI0/XI15/XI7/MM2_g N_VSS_XI0/XI15/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM3 N_XI0/XI15/XI7/NET33_XI0/XI15/XI7/MM3_d
+ N_WL<26>_XI0/XI15/XI7/MM3_g N_BLN<8>_XI0/XI15/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM0 N_XI0/XI15/XI7/NET34_XI0/XI15/XI7/MM0_d
+ N_WL<26>_XI0/XI15/XI7/MM0_g N_BL<8>_XI0/XI15/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM1 N_XI0/XI15/XI7/NET33_XI0/XI15/XI7/MM1_d
+ N_XI0/XI15/XI7/NET34_XI0/XI15/XI7/MM1_g N_VSS_XI0/XI15/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM9 N_XI0/XI15/XI7/NET36_XI0/XI15/XI7/MM9_d
+ N_WL<27>_XI0/XI15/XI7/MM9_g N_BL<8>_XI0/XI15/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM6 N_XI0/XI15/XI7/NET35_XI0/XI15/XI7/MM6_d
+ N_XI0/XI15/XI7/NET36_XI0/XI15/XI7/MM6_g N_VSS_XI0/XI15/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM7 N_XI0/XI15/XI7/NET36_XI0/XI15/XI7/MM7_d
+ N_XI0/XI15/XI7/NET35_XI0/XI15/XI7/MM7_g N_VSS_XI0/XI15/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM8 N_XI0/XI15/XI7/NET35_XI0/XI15/XI7/MM8_d
+ N_WL<27>_XI0/XI15/XI7/MM8_g N_BLN<8>_XI0/XI15/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI7/MM5 N_XI0/XI15/XI7/NET34_XI0/XI15/XI7/MM5_d
+ N_XI0/XI15/XI7/NET33_XI0/XI15/XI7/MM5_g N_VDD_XI0/XI15/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI7/MM4 N_XI0/XI15/XI7/NET33_XI0/XI15/XI7/MM4_d
+ N_XI0/XI15/XI7/NET34_XI0/XI15/XI7/MM4_g N_VDD_XI0/XI15/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI7/MM10 N_XI0/XI15/XI7/NET35_XI0/XI15/XI7/MM10_d
+ N_XI0/XI15/XI7/NET36_XI0/XI15/XI7/MM10_g N_VDD_XI0/XI15/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI7/MM11 N_XI0/XI15/XI7/NET36_XI0/XI15/XI7/MM11_d
+ N_XI0/XI15/XI7/NET35_XI0/XI15/XI7/MM11_g N_VDD_XI0/XI15/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI8/MM2 N_XI0/XI15/XI8/NET34_XI0/XI15/XI8/MM2_d
+ N_XI0/XI15/XI8/NET33_XI0/XI15/XI8/MM2_g N_VSS_XI0/XI15/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM3 N_XI0/XI15/XI8/NET33_XI0/XI15/XI8/MM3_d
+ N_WL<26>_XI0/XI15/XI8/MM3_g N_BLN<7>_XI0/XI15/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM0 N_XI0/XI15/XI8/NET34_XI0/XI15/XI8/MM0_d
+ N_WL<26>_XI0/XI15/XI8/MM0_g N_BL<7>_XI0/XI15/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM1 N_XI0/XI15/XI8/NET33_XI0/XI15/XI8/MM1_d
+ N_XI0/XI15/XI8/NET34_XI0/XI15/XI8/MM1_g N_VSS_XI0/XI15/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM9 N_XI0/XI15/XI8/NET36_XI0/XI15/XI8/MM9_d
+ N_WL<27>_XI0/XI15/XI8/MM9_g N_BL<7>_XI0/XI15/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM6 N_XI0/XI15/XI8/NET35_XI0/XI15/XI8/MM6_d
+ N_XI0/XI15/XI8/NET36_XI0/XI15/XI8/MM6_g N_VSS_XI0/XI15/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM7 N_XI0/XI15/XI8/NET36_XI0/XI15/XI8/MM7_d
+ N_XI0/XI15/XI8/NET35_XI0/XI15/XI8/MM7_g N_VSS_XI0/XI15/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM8 N_XI0/XI15/XI8/NET35_XI0/XI15/XI8/MM8_d
+ N_WL<27>_XI0/XI15/XI8/MM8_g N_BLN<7>_XI0/XI15/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI8/MM5 N_XI0/XI15/XI8/NET34_XI0/XI15/XI8/MM5_d
+ N_XI0/XI15/XI8/NET33_XI0/XI15/XI8/MM5_g N_VDD_XI0/XI15/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI8/MM4 N_XI0/XI15/XI8/NET33_XI0/XI15/XI8/MM4_d
+ N_XI0/XI15/XI8/NET34_XI0/XI15/XI8/MM4_g N_VDD_XI0/XI15/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI8/MM10 N_XI0/XI15/XI8/NET35_XI0/XI15/XI8/MM10_d
+ N_XI0/XI15/XI8/NET36_XI0/XI15/XI8/MM10_g N_VDD_XI0/XI15/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI8/MM11 N_XI0/XI15/XI8/NET36_XI0/XI15/XI8/MM11_d
+ N_XI0/XI15/XI8/NET35_XI0/XI15/XI8/MM11_g N_VDD_XI0/XI15/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI9/MM2 N_XI0/XI15/XI9/NET34_XI0/XI15/XI9/MM2_d
+ N_XI0/XI15/XI9/NET33_XI0/XI15/XI9/MM2_g N_VSS_XI0/XI15/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM3 N_XI0/XI15/XI9/NET33_XI0/XI15/XI9/MM3_d
+ N_WL<26>_XI0/XI15/XI9/MM3_g N_BLN<6>_XI0/XI15/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM0 N_XI0/XI15/XI9/NET34_XI0/XI15/XI9/MM0_d
+ N_WL<26>_XI0/XI15/XI9/MM0_g N_BL<6>_XI0/XI15/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM1 N_XI0/XI15/XI9/NET33_XI0/XI15/XI9/MM1_d
+ N_XI0/XI15/XI9/NET34_XI0/XI15/XI9/MM1_g N_VSS_XI0/XI15/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM9 N_XI0/XI15/XI9/NET36_XI0/XI15/XI9/MM9_d
+ N_WL<27>_XI0/XI15/XI9/MM9_g N_BL<6>_XI0/XI15/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM6 N_XI0/XI15/XI9/NET35_XI0/XI15/XI9/MM6_d
+ N_XI0/XI15/XI9/NET36_XI0/XI15/XI9/MM6_g N_VSS_XI0/XI15/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM7 N_XI0/XI15/XI9/NET36_XI0/XI15/XI9/MM7_d
+ N_XI0/XI15/XI9/NET35_XI0/XI15/XI9/MM7_g N_VSS_XI0/XI15/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM8 N_XI0/XI15/XI9/NET35_XI0/XI15/XI9/MM8_d
+ N_WL<27>_XI0/XI15/XI9/MM8_g N_BLN<6>_XI0/XI15/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI9/MM5 N_XI0/XI15/XI9/NET34_XI0/XI15/XI9/MM5_d
+ N_XI0/XI15/XI9/NET33_XI0/XI15/XI9/MM5_g N_VDD_XI0/XI15/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI9/MM4 N_XI0/XI15/XI9/NET33_XI0/XI15/XI9/MM4_d
+ N_XI0/XI15/XI9/NET34_XI0/XI15/XI9/MM4_g N_VDD_XI0/XI15/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI9/MM10 N_XI0/XI15/XI9/NET35_XI0/XI15/XI9/MM10_d
+ N_XI0/XI15/XI9/NET36_XI0/XI15/XI9/MM10_g N_VDD_XI0/XI15/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI9/MM11 N_XI0/XI15/XI9/NET36_XI0/XI15/XI9/MM11_d
+ N_XI0/XI15/XI9/NET35_XI0/XI15/XI9/MM11_g N_VDD_XI0/XI15/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI10/MM2 N_XI0/XI15/XI10/NET34_XI0/XI15/XI10/MM2_d
+ N_XI0/XI15/XI10/NET33_XI0/XI15/XI10/MM2_g N_VSS_XI0/XI15/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM3 N_XI0/XI15/XI10/NET33_XI0/XI15/XI10/MM3_d
+ N_WL<26>_XI0/XI15/XI10/MM3_g N_BLN<5>_XI0/XI15/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM0 N_XI0/XI15/XI10/NET34_XI0/XI15/XI10/MM0_d
+ N_WL<26>_XI0/XI15/XI10/MM0_g N_BL<5>_XI0/XI15/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM1 N_XI0/XI15/XI10/NET33_XI0/XI15/XI10/MM1_d
+ N_XI0/XI15/XI10/NET34_XI0/XI15/XI10/MM1_g N_VSS_XI0/XI15/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM9 N_XI0/XI15/XI10/NET36_XI0/XI15/XI10/MM9_d
+ N_WL<27>_XI0/XI15/XI10/MM9_g N_BL<5>_XI0/XI15/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM6 N_XI0/XI15/XI10/NET35_XI0/XI15/XI10/MM6_d
+ N_XI0/XI15/XI10/NET36_XI0/XI15/XI10/MM6_g N_VSS_XI0/XI15/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM7 N_XI0/XI15/XI10/NET36_XI0/XI15/XI10/MM7_d
+ N_XI0/XI15/XI10/NET35_XI0/XI15/XI10/MM7_g N_VSS_XI0/XI15/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM8 N_XI0/XI15/XI10/NET35_XI0/XI15/XI10/MM8_d
+ N_WL<27>_XI0/XI15/XI10/MM8_g N_BLN<5>_XI0/XI15/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI10/MM5 N_XI0/XI15/XI10/NET34_XI0/XI15/XI10/MM5_d
+ N_XI0/XI15/XI10/NET33_XI0/XI15/XI10/MM5_g N_VDD_XI0/XI15/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI10/MM4 N_XI0/XI15/XI10/NET33_XI0/XI15/XI10/MM4_d
+ N_XI0/XI15/XI10/NET34_XI0/XI15/XI10/MM4_g N_VDD_XI0/XI15/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI10/MM10 N_XI0/XI15/XI10/NET35_XI0/XI15/XI10/MM10_d
+ N_XI0/XI15/XI10/NET36_XI0/XI15/XI10/MM10_g N_VDD_XI0/XI15/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI10/MM11 N_XI0/XI15/XI10/NET36_XI0/XI15/XI10/MM11_d
+ N_XI0/XI15/XI10/NET35_XI0/XI15/XI10/MM11_g N_VDD_XI0/XI15/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI11/MM2 N_XI0/XI15/XI11/NET34_XI0/XI15/XI11/MM2_d
+ N_XI0/XI15/XI11/NET33_XI0/XI15/XI11/MM2_g N_VSS_XI0/XI15/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM3 N_XI0/XI15/XI11/NET33_XI0/XI15/XI11/MM3_d
+ N_WL<26>_XI0/XI15/XI11/MM3_g N_BLN<4>_XI0/XI15/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM0 N_XI0/XI15/XI11/NET34_XI0/XI15/XI11/MM0_d
+ N_WL<26>_XI0/XI15/XI11/MM0_g N_BL<4>_XI0/XI15/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM1 N_XI0/XI15/XI11/NET33_XI0/XI15/XI11/MM1_d
+ N_XI0/XI15/XI11/NET34_XI0/XI15/XI11/MM1_g N_VSS_XI0/XI15/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM9 N_XI0/XI15/XI11/NET36_XI0/XI15/XI11/MM9_d
+ N_WL<27>_XI0/XI15/XI11/MM9_g N_BL<4>_XI0/XI15/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM6 N_XI0/XI15/XI11/NET35_XI0/XI15/XI11/MM6_d
+ N_XI0/XI15/XI11/NET36_XI0/XI15/XI11/MM6_g N_VSS_XI0/XI15/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM7 N_XI0/XI15/XI11/NET36_XI0/XI15/XI11/MM7_d
+ N_XI0/XI15/XI11/NET35_XI0/XI15/XI11/MM7_g N_VSS_XI0/XI15/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM8 N_XI0/XI15/XI11/NET35_XI0/XI15/XI11/MM8_d
+ N_WL<27>_XI0/XI15/XI11/MM8_g N_BLN<4>_XI0/XI15/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI11/MM5 N_XI0/XI15/XI11/NET34_XI0/XI15/XI11/MM5_d
+ N_XI0/XI15/XI11/NET33_XI0/XI15/XI11/MM5_g N_VDD_XI0/XI15/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI11/MM4 N_XI0/XI15/XI11/NET33_XI0/XI15/XI11/MM4_d
+ N_XI0/XI15/XI11/NET34_XI0/XI15/XI11/MM4_g N_VDD_XI0/XI15/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI11/MM10 N_XI0/XI15/XI11/NET35_XI0/XI15/XI11/MM10_d
+ N_XI0/XI15/XI11/NET36_XI0/XI15/XI11/MM10_g N_VDD_XI0/XI15/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI11/MM11 N_XI0/XI15/XI11/NET36_XI0/XI15/XI11/MM11_d
+ N_XI0/XI15/XI11/NET35_XI0/XI15/XI11/MM11_g N_VDD_XI0/XI15/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI12/MM2 N_XI0/XI15/XI12/NET34_XI0/XI15/XI12/MM2_d
+ N_XI0/XI15/XI12/NET33_XI0/XI15/XI12/MM2_g N_VSS_XI0/XI15/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM3 N_XI0/XI15/XI12/NET33_XI0/XI15/XI12/MM3_d
+ N_WL<26>_XI0/XI15/XI12/MM3_g N_BLN<3>_XI0/XI15/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM0 N_XI0/XI15/XI12/NET34_XI0/XI15/XI12/MM0_d
+ N_WL<26>_XI0/XI15/XI12/MM0_g N_BL<3>_XI0/XI15/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM1 N_XI0/XI15/XI12/NET33_XI0/XI15/XI12/MM1_d
+ N_XI0/XI15/XI12/NET34_XI0/XI15/XI12/MM1_g N_VSS_XI0/XI15/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM9 N_XI0/XI15/XI12/NET36_XI0/XI15/XI12/MM9_d
+ N_WL<27>_XI0/XI15/XI12/MM9_g N_BL<3>_XI0/XI15/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM6 N_XI0/XI15/XI12/NET35_XI0/XI15/XI12/MM6_d
+ N_XI0/XI15/XI12/NET36_XI0/XI15/XI12/MM6_g N_VSS_XI0/XI15/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM7 N_XI0/XI15/XI12/NET36_XI0/XI15/XI12/MM7_d
+ N_XI0/XI15/XI12/NET35_XI0/XI15/XI12/MM7_g N_VSS_XI0/XI15/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM8 N_XI0/XI15/XI12/NET35_XI0/XI15/XI12/MM8_d
+ N_WL<27>_XI0/XI15/XI12/MM8_g N_BLN<3>_XI0/XI15/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI12/MM5 N_XI0/XI15/XI12/NET34_XI0/XI15/XI12/MM5_d
+ N_XI0/XI15/XI12/NET33_XI0/XI15/XI12/MM5_g N_VDD_XI0/XI15/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI12/MM4 N_XI0/XI15/XI12/NET33_XI0/XI15/XI12/MM4_d
+ N_XI0/XI15/XI12/NET34_XI0/XI15/XI12/MM4_g N_VDD_XI0/XI15/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI12/MM10 N_XI0/XI15/XI12/NET35_XI0/XI15/XI12/MM10_d
+ N_XI0/XI15/XI12/NET36_XI0/XI15/XI12/MM10_g N_VDD_XI0/XI15/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI12/MM11 N_XI0/XI15/XI12/NET36_XI0/XI15/XI12/MM11_d
+ N_XI0/XI15/XI12/NET35_XI0/XI15/XI12/MM11_g N_VDD_XI0/XI15/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI13/MM2 N_XI0/XI15/XI13/NET34_XI0/XI15/XI13/MM2_d
+ N_XI0/XI15/XI13/NET33_XI0/XI15/XI13/MM2_g N_VSS_XI0/XI15/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM3 N_XI0/XI15/XI13/NET33_XI0/XI15/XI13/MM3_d
+ N_WL<26>_XI0/XI15/XI13/MM3_g N_BLN<2>_XI0/XI15/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM0 N_XI0/XI15/XI13/NET34_XI0/XI15/XI13/MM0_d
+ N_WL<26>_XI0/XI15/XI13/MM0_g N_BL<2>_XI0/XI15/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM1 N_XI0/XI15/XI13/NET33_XI0/XI15/XI13/MM1_d
+ N_XI0/XI15/XI13/NET34_XI0/XI15/XI13/MM1_g N_VSS_XI0/XI15/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM9 N_XI0/XI15/XI13/NET36_XI0/XI15/XI13/MM9_d
+ N_WL<27>_XI0/XI15/XI13/MM9_g N_BL<2>_XI0/XI15/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM6 N_XI0/XI15/XI13/NET35_XI0/XI15/XI13/MM6_d
+ N_XI0/XI15/XI13/NET36_XI0/XI15/XI13/MM6_g N_VSS_XI0/XI15/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM7 N_XI0/XI15/XI13/NET36_XI0/XI15/XI13/MM7_d
+ N_XI0/XI15/XI13/NET35_XI0/XI15/XI13/MM7_g N_VSS_XI0/XI15/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM8 N_XI0/XI15/XI13/NET35_XI0/XI15/XI13/MM8_d
+ N_WL<27>_XI0/XI15/XI13/MM8_g N_BLN<2>_XI0/XI15/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI13/MM5 N_XI0/XI15/XI13/NET34_XI0/XI15/XI13/MM5_d
+ N_XI0/XI15/XI13/NET33_XI0/XI15/XI13/MM5_g N_VDD_XI0/XI15/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI13/MM4 N_XI0/XI15/XI13/NET33_XI0/XI15/XI13/MM4_d
+ N_XI0/XI15/XI13/NET34_XI0/XI15/XI13/MM4_g N_VDD_XI0/XI15/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI13/MM10 N_XI0/XI15/XI13/NET35_XI0/XI15/XI13/MM10_d
+ N_XI0/XI15/XI13/NET36_XI0/XI15/XI13/MM10_g N_VDD_XI0/XI15/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI13/MM11 N_XI0/XI15/XI13/NET36_XI0/XI15/XI13/MM11_d
+ N_XI0/XI15/XI13/NET35_XI0/XI15/XI13/MM11_g N_VDD_XI0/XI15/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI14/MM2 N_XI0/XI15/XI14/NET34_XI0/XI15/XI14/MM2_d
+ N_XI0/XI15/XI14/NET33_XI0/XI15/XI14/MM2_g N_VSS_XI0/XI15/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM3 N_XI0/XI15/XI14/NET33_XI0/XI15/XI14/MM3_d
+ N_WL<26>_XI0/XI15/XI14/MM3_g N_BLN<1>_XI0/XI15/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM0 N_XI0/XI15/XI14/NET34_XI0/XI15/XI14/MM0_d
+ N_WL<26>_XI0/XI15/XI14/MM0_g N_BL<1>_XI0/XI15/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM1 N_XI0/XI15/XI14/NET33_XI0/XI15/XI14/MM1_d
+ N_XI0/XI15/XI14/NET34_XI0/XI15/XI14/MM1_g N_VSS_XI0/XI15/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM9 N_XI0/XI15/XI14/NET36_XI0/XI15/XI14/MM9_d
+ N_WL<27>_XI0/XI15/XI14/MM9_g N_BL<1>_XI0/XI15/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM6 N_XI0/XI15/XI14/NET35_XI0/XI15/XI14/MM6_d
+ N_XI0/XI15/XI14/NET36_XI0/XI15/XI14/MM6_g N_VSS_XI0/XI15/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM7 N_XI0/XI15/XI14/NET36_XI0/XI15/XI14/MM7_d
+ N_XI0/XI15/XI14/NET35_XI0/XI15/XI14/MM7_g N_VSS_XI0/XI15/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM8 N_XI0/XI15/XI14/NET35_XI0/XI15/XI14/MM8_d
+ N_WL<27>_XI0/XI15/XI14/MM8_g N_BLN<1>_XI0/XI15/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI14/MM5 N_XI0/XI15/XI14/NET34_XI0/XI15/XI14/MM5_d
+ N_XI0/XI15/XI14/NET33_XI0/XI15/XI14/MM5_g N_VDD_XI0/XI15/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI14/MM4 N_XI0/XI15/XI14/NET33_XI0/XI15/XI14/MM4_d
+ N_XI0/XI15/XI14/NET34_XI0/XI15/XI14/MM4_g N_VDD_XI0/XI15/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI14/MM10 N_XI0/XI15/XI14/NET35_XI0/XI15/XI14/MM10_d
+ N_XI0/XI15/XI14/NET36_XI0/XI15/XI14/MM10_g N_VDD_XI0/XI15/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI14/MM11 N_XI0/XI15/XI14/NET36_XI0/XI15/XI14/MM11_d
+ N_XI0/XI15/XI14/NET35_XI0/XI15/XI14/MM11_g N_VDD_XI0/XI15/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI15/MM2 N_XI0/XI15/XI15/NET34_XI0/XI15/XI15/MM2_d
+ N_XI0/XI15/XI15/NET33_XI0/XI15/XI15/MM2_g N_VSS_XI0/XI15/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM3 N_XI0/XI15/XI15/NET33_XI0/XI15/XI15/MM3_d
+ N_WL<26>_XI0/XI15/XI15/MM3_g N_BLN<0>_XI0/XI15/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM0 N_XI0/XI15/XI15/NET34_XI0/XI15/XI15/MM0_d
+ N_WL<26>_XI0/XI15/XI15/MM0_g N_BL<0>_XI0/XI15/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM1 N_XI0/XI15/XI15/NET33_XI0/XI15/XI15/MM1_d
+ N_XI0/XI15/XI15/NET34_XI0/XI15/XI15/MM1_g N_VSS_XI0/XI15/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM9 N_XI0/XI15/XI15/NET36_XI0/XI15/XI15/MM9_d
+ N_WL<27>_XI0/XI15/XI15/MM9_g N_BL<0>_XI0/XI15/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM6 N_XI0/XI15/XI15/NET35_XI0/XI15/XI15/MM6_d
+ N_XI0/XI15/XI15/NET36_XI0/XI15/XI15/MM6_g N_VSS_XI0/XI15/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM7 N_XI0/XI15/XI15/NET36_XI0/XI15/XI15/MM7_d
+ N_XI0/XI15/XI15/NET35_XI0/XI15/XI15/MM7_g N_VSS_XI0/XI15/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM8 N_XI0/XI15/XI15/NET35_XI0/XI15/XI15/MM8_d
+ N_WL<27>_XI0/XI15/XI15/MM8_g N_BLN<0>_XI0/XI15/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/XI15/MM5 N_XI0/XI15/XI15/NET34_XI0/XI15/XI15/MM5_d
+ N_XI0/XI15/XI15/NET33_XI0/XI15/XI15/MM5_g N_VDD_XI0/XI15/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI15/MM4 N_XI0/XI15/XI15/NET33_XI0/XI15/XI15/MM4_d
+ N_XI0/XI15/XI15/NET34_XI0/XI15/XI15/MM4_g N_VDD_XI0/XI15/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI15/MM10 N_XI0/XI15/XI15/NET35_XI0/XI15/XI15/MM10_d
+ N_XI0/XI15/XI15/NET36_XI0/XI15/XI15/MM10_g N_VDD_XI0/XI15/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/XI15/MM11 N_XI0/XI15/XI15/NET36_XI0/XI15/XI15/MM11_d
+ N_XI0/XI15/XI15/NET35_XI0/XI15/XI15/MM11_g N_VDD_XI0/XI15/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI0/MM2 N_XI0/XI16/XI0/NET34_XI0/XI16/XI0/MM2_d
+ N_XI0/XI16/XI0/NET33_XI0/XI16/XI0/MM2_g N_VSS_XI0/XI16/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM3 N_XI0/XI16/XI0/NET33_XI0/XI16/XI0/MM3_d
+ N_WL<28>_XI0/XI16/XI0/MM3_g N_BLN<15>_XI0/XI16/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM0 N_XI0/XI16/XI0/NET34_XI0/XI16/XI0/MM0_d
+ N_WL<28>_XI0/XI16/XI0/MM0_g N_BL<15>_XI0/XI16/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM1 N_XI0/XI16/XI0/NET33_XI0/XI16/XI0/MM1_d
+ N_XI0/XI16/XI0/NET34_XI0/XI16/XI0/MM1_g N_VSS_XI0/XI16/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM9 N_XI0/XI16/XI0/NET36_XI0/XI16/XI0/MM9_d
+ N_WL<29>_XI0/XI16/XI0/MM9_g N_BL<15>_XI0/XI16/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM6 N_XI0/XI16/XI0/NET35_XI0/XI16/XI0/MM6_d
+ N_XI0/XI16/XI0/NET36_XI0/XI16/XI0/MM6_g N_VSS_XI0/XI16/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM7 N_XI0/XI16/XI0/NET36_XI0/XI16/XI0/MM7_d
+ N_XI0/XI16/XI0/NET35_XI0/XI16/XI0/MM7_g N_VSS_XI0/XI16/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM8 N_XI0/XI16/XI0/NET35_XI0/XI16/XI0/MM8_d
+ N_WL<29>_XI0/XI16/XI0/MM8_g N_BLN<15>_XI0/XI16/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI0/MM5 N_XI0/XI16/XI0/NET34_XI0/XI16/XI0/MM5_d
+ N_XI0/XI16/XI0/NET33_XI0/XI16/XI0/MM5_g N_VDD_XI0/XI16/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI0/MM4 N_XI0/XI16/XI0/NET33_XI0/XI16/XI0/MM4_d
+ N_XI0/XI16/XI0/NET34_XI0/XI16/XI0/MM4_g N_VDD_XI0/XI16/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI0/MM10 N_XI0/XI16/XI0/NET35_XI0/XI16/XI0/MM10_d
+ N_XI0/XI16/XI0/NET36_XI0/XI16/XI0/MM10_g N_VDD_XI0/XI16/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI0/MM11 N_XI0/XI16/XI0/NET36_XI0/XI16/XI0/MM11_d
+ N_XI0/XI16/XI0/NET35_XI0/XI16/XI0/MM11_g N_VDD_XI0/XI16/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI1/MM2 N_XI0/XI16/XI1/NET34_XI0/XI16/XI1/MM2_d
+ N_XI0/XI16/XI1/NET33_XI0/XI16/XI1/MM2_g N_VSS_XI0/XI16/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM3 N_XI0/XI16/XI1/NET33_XI0/XI16/XI1/MM3_d
+ N_WL<28>_XI0/XI16/XI1/MM3_g N_BLN<14>_XI0/XI16/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM0 N_XI0/XI16/XI1/NET34_XI0/XI16/XI1/MM0_d
+ N_WL<28>_XI0/XI16/XI1/MM0_g N_BL<14>_XI0/XI16/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM1 N_XI0/XI16/XI1/NET33_XI0/XI16/XI1/MM1_d
+ N_XI0/XI16/XI1/NET34_XI0/XI16/XI1/MM1_g N_VSS_XI0/XI16/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM9 N_XI0/XI16/XI1/NET36_XI0/XI16/XI1/MM9_d
+ N_WL<29>_XI0/XI16/XI1/MM9_g N_BL<14>_XI0/XI16/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM6 N_XI0/XI16/XI1/NET35_XI0/XI16/XI1/MM6_d
+ N_XI0/XI16/XI1/NET36_XI0/XI16/XI1/MM6_g N_VSS_XI0/XI16/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM7 N_XI0/XI16/XI1/NET36_XI0/XI16/XI1/MM7_d
+ N_XI0/XI16/XI1/NET35_XI0/XI16/XI1/MM7_g N_VSS_XI0/XI16/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM8 N_XI0/XI16/XI1/NET35_XI0/XI16/XI1/MM8_d
+ N_WL<29>_XI0/XI16/XI1/MM8_g N_BLN<14>_XI0/XI16/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI1/MM5 N_XI0/XI16/XI1/NET34_XI0/XI16/XI1/MM5_d
+ N_XI0/XI16/XI1/NET33_XI0/XI16/XI1/MM5_g N_VDD_XI0/XI16/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI1/MM4 N_XI0/XI16/XI1/NET33_XI0/XI16/XI1/MM4_d
+ N_XI0/XI16/XI1/NET34_XI0/XI16/XI1/MM4_g N_VDD_XI0/XI16/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI1/MM10 N_XI0/XI16/XI1/NET35_XI0/XI16/XI1/MM10_d
+ N_XI0/XI16/XI1/NET36_XI0/XI16/XI1/MM10_g N_VDD_XI0/XI16/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI1/MM11 N_XI0/XI16/XI1/NET36_XI0/XI16/XI1/MM11_d
+ N_XI0/XI16/XI1/NET35_XI0/XI16/XI1/MM11_g N_VDD_XI0/XI16/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI2/MM2 N_XI0/XI16/XI2/NET34_XI0/XI16/XI2/MM2_d
+ N_XI0/XI16/XI2/NET33_XI0/XI16/XI2/MM2_g N_VSS_XI0/XI16/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM3 N_XI0/XI16/XI2/NET33_XI0/XI16/XI2/MM3_d
+ N_WL<28>_XI0/XI16/XI2/MM3_g N_BLN<13>_XI0/XI16/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM0 N_XI0/XI16/XI2/NET34_XI0/XI16/XI2/MM0_d
+ N_WL<28>_XI0/XI16/XI2/MM0_g N_BL<13>_XI0/XI16/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM1 N_XI0/XI16/XI2/NET33_XI0/XI16/XI2/MM1_d
+ N_XI0/XI16/XI2/NET34_XI0/XI16/XI2/MM1_g N_VSS_XI0/XI16/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM9 N_XI0/XI16/XI2/NET36_XI0/XI16/XI2/MM9_d
+ N_WL<29>_XI0/XI16/XI2/MM9_g N_BL<13>_XI0/XI16/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM6 N_XI0/XI16/XI2/NET35_XI0/XI16/XI2/MM6_d
+ N_XI0/XI16/XI2/NET36_XI0/XI16/XI2/MM6_g N_VSS_XI0/XI16/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM7 N_XI0/XI16/XI2/NET36_XI0/XI16/XI2/MM7_d
+ N_XI0/XI16/XI2/NET35_XI0/XI16/XI2/MM7_g N_VSS_XI0/XI16/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM8 N_XI0/XI16/XI2/NET35_XI0/XI16/XI2/MM8_d
+ N_WL<29>_XI0/XI16/XI2/MM8_g N_BLN<13>_XI0/XI16/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI2/MM5 N_XI0/XI16/XI2/NET34_XI0/XI16/XI2/MM5_d
+ N_XI0/XI16/XI2/NET33_XI0/XI16/XI2/MM5_g N_VDD_XI0/XI16/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI2/MM4 N_XI0/XI16/XI2/NET33_XI0/XI16/XI2/MM4_d
+ N_XI0/XI16/XI2/NET34_XI0/XI16/XI2/MM4_g N_VDD_XI0/XI16/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI2/MM10 N_XI0/XI16/XI2/NET35_XI0/XI16/XI2/MM10_d
+ N_XI0/XI16/XI2/NET36_XI0/XI16/XI2/MM10_g N_VDD_XI0/XI16/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI2/MM11 N_XI0/XI16/XI2/NET36_XI0/XI16/XI2/MM11_d
+ N_XI0/XI16/XI2/NET35_XI0/XI16/XI2/MM11_g N_VDD_XI0/XI16/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI3/MM2 N_XI0/XI16/XI3/NET34_XI0/XI16/XI3/MM2_d
+ N_XI0/XI16/XI3/NET33_XI0/XI16/XI3/MM2_g N_VSS_XI0/XI16/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM3 N_XI0/XI16/XI3/NET33_XI0/XI16/XI3/MM3_d
+ N_WL<28>_XI0/XI16/XI3/MM3_g N_BLN<12>_XI0/XI16/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM0 N_XI0/XI16/XI3/NET34_XI0/XI16/XI3/MM0_d
+ N_WL<28>_XI0/XI16/XI3/MM0_g N_BL<12>_XI0/XI16/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM1 N_XI0/XI16/XI3/NET33_XI0/XI16/XI3/MM1_d
+ N_XI0/XI16/XI3/NET34_XI0/XI16/XI3/MM1_g N_VSS_XI0/XI16/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM9 N_XI0/XI16/XI3/NET36_XI0/XI16/XI3/MM9_d
+ N_WL<29>_XI0/XI16/XI3/MM9_g N_BL<12>_XI0/XI16/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM6 N_XI0/XI16/XI3/NET35_XI0/XI16/XI3/MM6_d
+ N_XI0/XI16/XI3/NET36_XI0/XI16/XI3/MM6_g N_VSS_XI0/XI16/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM7 N_XI0/XI16/XI3/NET36_XI0/XI16/XI3/MM7_d
+ N_XI0/XI16/XI3/NET35_XI0/XI16/XI3/MM7_g N_VSS_XI0/XI16/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM8 N_XI0/XI16/XI3/NET35_XI0/XI16/XI3/MM8_d
+ N_WL<29>_XI0/XI16/XI3/MM8_g N_BLN<12>_XI0/XI16/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI3/MM5 N_XI0/XI16/XI3/NET34_XI0/XI16/XI3/MM5_d
+ N_XI0/XI16/XI3/NET33_XI0/XI16/XI3/MM5_g N_VDD_XI0/XI16/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI3/MM4 N_XI0/XI16/XI3/NET33_XI0/XI16/XI3/MM4_d
+ N_XI0/XI16/XI3/NET34_XI0/XI16/XI3/MM4_g N_VDD_XI0/XI16/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI3/MM10 N_XI0/XI16/XI3/NET35_XI0/XI16/XI3/MM10_d
+ N_XI0/XI16/XI3/NET36_XI0/XI16/XI3/MM10_g N_VDD_XI0/XI16/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI3/MM11 N_XI0/XI16/XI3/NET36_XI0/XI16/XI3/MM11_d
+ N_XI0/XI16/XI3/NET35_XI0/XI16/XI3/MM11_g N_VDD_XI0/XI16/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI4/MM2 N_XI0/XI16/XI4/NET34_XI0/XI16/XI4/MM2_d
+ N_XI0/XI16/XI4/NET33_XI0/XI16/XI4/MM2_g N_VSS_XI0/XI16/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM3 N_XI0/XI16/XI4/NET33_XI0/XI16/XI4/MM3_d
+ N_WL<28>_XI0/XI16/XI4/MM3_g N_BLN<11>_XI0/XI16/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM0 N_XI0/XI16/XI4/NET34_XI0/XI16/XI4/MM0_d
+ N_WL<28>_XI0/XI16/XI4/MM0_g N_BL<11>_XI0/XI16/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM1 N_XI0/XI16/XI4/NET33_XI0/XI16/XI4/MM1_d
+ N_XI0/XI16/XI4/NET34_XI0/XI16/XI4/MM1_g N_VSS_XI0/XI16/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM9 N_XI0/XI16/XI4/NET36_XI0/XI16/XI4/MM9_d
+ N_WL<29>_XI0/XI16/XI4/MM9_g N_BL<11>_XI0/XI16/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM6 N_XI0/XI16/XI4/NET35_XI0/XI16/XI4/MM6_d
+ N_XI0/XI16/XI4/NET36_XI0/XI16/XI4/MM6_g N_VSS_XI0/XI16/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM7 N_XI0/XI16/XI4/NET36_XI0/XI16/XI4/MM7_d
+ N_XI0/XI16/XI4/NET35_XI0/XI16/XI4/MM7_g N_VSS_XI0/XI16/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM8 N_XI0/XI16/XI4/NET35_XI0/XI16/XI4/MM8_d
+ N_WL<29>_XI0/XI16/XI4/MM8_g N_BLN<11>_XI0/XI16/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI4/MM5 N_XI0/XI16/XI4/NET34_XI0/XI16/XI4/MM5_d
+ N_XI0/XI16/XI4/NET33_XI0/XI16/XI4/MM5_g N_VDD_XI0/XI16/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI4/MM4 N_XI0/XI16/XI4/NET33_XI0/XI16/XI4/MM4_d
+ N_XI0/XI16/XI4/NET34_XI0/XI16/XI4/MM4_g N_VDD_XI0/XI16/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI4/MM10 N_XI0/XI16/XI4/NET35_XI0/XI16/XI4/MM10_d
+ N_XI0/XI16/XI4/NET36_XI0/XI16/XI4/MM10_g N_VDD_XI0/XI16/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI4/MM11 N_XI0/XI16/XI4/NET36_XI0/XI16/XI4/MM11_d
+ N_XI0/XI16/XI4/NET35_XI0/XI16/XI4/MM11_g N_VDD_XI0/XI16/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI5/MM2 N_XI0/XI16/XI5/NET34_XI0/XI16/XI5/MM2_d
+ N_XI0/XI16/XI5/NET33_XI0/XI16/XI5/MM2_g N_VSS_XI0/XI16/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM3 N_XI0/XI16/XI5/NET33_XI0/XI16/XI5/MM3_d
+ N_WL<28>_XI0/XI16/XI5/MM3_g N_BLN<10>_XI0/XI16/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM0 N_XI0/XI16/XI5/NET34_XI0/XI16/XI5/MM0_d
+ N_WL<28>_XI0/XI16/XI5/MM0_g N_BL<10>_XI0/XI16/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM1 N_XI0/XI16/XI5/NET33_XI0/XI16/XI5/MM1_d
+ N_XI0/XI16/XI5/NET34_XI0/XI16/XI5/MM1_g N_VSS_XI0/XI16/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM9 N_XI0/XI16/XI5/NET36_XI0/XI16/XI5/MM9_d
+ N_WL<29>_XI0/XI16/XI5/MM9_g N_BL<10>_XI0/XI16/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM6 N_XI0/XI16/XI5/NET35_XI0/XI16/XI5/MM6_d
+ N_XI0/XI16/XI5/NET36_XI0/XI16/XI5/MM6_g N_VSS_XI0/XI16/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM7 N_XI0/XI16/XI5/NET36_XI0/XI16/XI5/MM7_d
+ N_XI0/XI16/XI5/NET35_XI0/XI16/XI5/MM7_g N_VSS_XI0/XI16/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM8 N_XI0/XI16/XI5/NET35_XI0/XI16/XI5/MM8_d
+ N_WL<29>_XI0/XI16/XI5/MM8_g N_BLN<10>_XI0/XI16/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI5/MM5 N_XI0/XI16/XI5/NET34_XI0/XI16/XI5/MM5_d
+ N_XI0/XI16/XI5/NET33_XI0/XI16/XI5/MM5_g N_VDD_XI0/XI16/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI5/MM4 N_XI0/XI16/XI5/NET33_XI0/XI16/XI5/MM4_d
+ N_XI0/XI16/XI5/NET34_XI0/XI16/XI5/MM4_g N_VDD_XI0/XI16/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI5/MM10 N_XI0/XI16/XI5/NET35_XI0/XI16/XI5/MM10_d
+ N_XI0/XI16/XI5/NET36_XI0/XI16/XI5/MM10_g N_VDD_XI0/XI16/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI5/MM11 N_XI0/XI16/XI5/NET36_XI0/XI16/XI5/MM11_d
+ N_XI0/XI16/XI5/NET35_XI0/XI16/XI5/MM11_g N_VDD_XI0/XI16/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI6/MM2 N_XI0/XI16/XI6/NET34_XI0/XI16/XI6/MM2_d
+ N_XI0/XI16/XI6/NET33_XI0/XI16/XI6/MM2_g N_VSS_XI0/XI16/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM3 N_XI0/XI16/XI6/NET33_XI0/XI16/XI6/MM3_d
+ N_WL<28>_XI0/XI16/XI6/MM3_g N_BLN<9>_XI0/XI16/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM0 N_XI0/XI16/XI6/NET34_XI0/XI16/XI6/MM0_d
+ N_WL<28>_XI0/XI16/XI6/MM0_g N_BL<9>_XI0/XI16/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM1 N_XI0/XI16/XI6/NET33_XI0/XI16/XI6/MM1_d
+ N_XI0/XI16/XI6/NET34_XI0/XI16/XI6/MM1_g N_VSS_XI0/XI16/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM9 N_XI0/XI16/XI6/NET36_XI0/XI16/XI6/MM9_d
+ N_WL<29>_XI0/XI16/XI6/MM9_g N_BL<9>_XI0/XI16/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM6 N_XI0/XI16/XI6/NET35_XI0/XI16/XI6/MM6_d
+ N_XI0/XI16/XI6/NET36_XI0/XI16/XI6/MM6_g N_VSS_XI0/XI16/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM7 N_XI0/XI16/XI6/NET36_XI0/XI16/XI6/MM7_d
+ N_XI0/XI16/XI6/NET35_XI0/XI16/XI6/MM7_g N_VSS_XI0/XI16/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM8 N_XI0/XI16/XI6/NET35_XI0/XI16/XI6/MM8_d
+ N_WL<29>_XI0/XI16/XI6/MM8_g N_BLN<9>_XI0/XI16/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI6/MM5 N_XI0/XI16/XI6/NET34_XI0/XI16/XI6/MM5_d
+ N_XI0/XI16/XI6/NET33_XI0/XI16/XI6/MM5_g N_VDD_XI0/XI16/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI6/MM4 N_XI0/XI16/XI6/NET33_XI0/XI16/XI6/MM4_d
+ N_XI0/XI16/XI6/NET34_XI0/XI16/XI6/MM4_g N_VDD_XI0/XI16/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI6/MM10 N_XI0/XI16/XI6/NET35_XI0/XI16/XI6/MM10_d
+ N_XI0/XI16/XI6/NET36_XI0/XI16/XI6/MM10_g N_VDD_XI0/XI16/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI6/MM11 N_XI0/XI16/XI6/NET36_XI0/XI16/XI6/MM11_d
+ N_XI0/XI16/XI6/NET35_XI0/XI16/XI6/MM11_g N_VDD_XI0/XI16/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI7/MM2 N_XI0/XI16/XI7/NET34_XI0/XI16/XI7/MM2_d
+ N_XI0/XI16/XI7/NET33_XI0/XI16/XI7/MM2_g N_VSS_XI0/XI16/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM3 N_XI0/XI16/XI7/NET33_XI0/XI16/XI7/MM3_d
+ N_WL<28>_XI0/XI16/XI7/MM3_g N_BLN<8>_XI0/XI16/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM0 N_XI0/XI16/XI7/NET34_XI0/XI16/XI7/MM0_d
+ N_WL<28>_XI0/XI16/XI7/MM0_g N_BL<8>_XI0/XI16/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM1 N_XI0/XI16/XI7/NET33_XI0/XI16/XI7/MM1_d
+ N_XI0/XI16/XI7/NET34_XI0/XI16/XI7/MM1_g N_VSS_XI0/XI16/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM9 N_XI0/XI16/XI7/NET36_XI0/XI16/XI7/MM9_d
+ N_WL<29>_XI0/XI16/XI7/MM9_g N_BL<8>_XI0/XI16/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM6 N_XI0/XI16/XI7/NET35_XI0/XI16/XI7/MM6_d
+ N_XI0/XI16/XI7/NET36_XI0/XI16/XI7/MM6_g N_VSS_XI0/XI16/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM7 N_XI0/XI16/XI7/NET36_XI0/XI16/XI7/MM7_d
+ N_XI0/XI16/XI7/NET35_XI0/XI16/XI7/MM7_g N_VSS_XI0/XI16/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM8 N_XI0/XI16/XI7/NET35_XI0/XI16/XI7/MM8_d
+ N_WL<29>_XI0/XI16/XI7/MM8_g N_BLN<8>_XI0/XI16/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI7/MM5 N_XI0/XI16/XI7/NET34_XI0/XI16/XI7/MM5_d
+ N_XI0/XI16/XI7/NET33_XI0/XI16/XI7/MM5_g N_VDD_XI0/XI16/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI7/MM4 N_XI0/XI16/XI7/NET33_XI0/XI16/XI7/MM4_d
+ N_XI0/XI16/XI7/NET34_XI0/XI16/XI7/MM4_g N_VDD_XI0/XI16/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI7/MM10 N_XI0/XI16/XI7/NET35_XI0/XI16/XI7/MM10_d
+ N_XI0/XI16/XI7/NET36_XI0/XI16/XI7/MM10_g N_VDD_XI0/XI16/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI7/MM11 N_XI0/XI16/XI7/NET36_XI0/XI16/XI7/MM11_d
+ N_XI0/XI16/XI7/NET35_XI0/XI16/XI7/MM11_g N_VDD_XI0/XI16/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI8/MM2 N_XI0/XI16/XI8/NET34_XI0/XI16/XI8/MM2_d
+ N_XI0/XI16/XI8/NET33_XI0/XI16/XI8/MM2_g N_VSS_XI0/XI16/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM3 N_XI0/XI16/XI8/NET33_XI0/XI16/XI8/MM3_d
+ N_WL<28>_XI0/XI16/XI8/MM3_g N_BLN<7>_XI0/XI16/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM0 N_XI0/XI16/XI8/NET34_XI0/XI16/XI8/MM0_d
+ N_WL<28>_XI0/XI16/XI8/MM0_g N_BL<7>_XI0/XI16/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM1 N_XI0/XI16/XI8/NET33_XI0/XI16/XI8/MM1_d
+ N_XI0/XI16/XI8/NET34_XI0/XI16/XI8/MM1_g N_VSS_XI0/XI16/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM9 N_XI0/XI16/XI8/NET36_XI0/XI16/XI8/MM9_d
+ N_WL<29>_XI0/XI16/XI8/MM9_g N_BL<7>_XI0/XI16/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM6 N_XI0/XI16/XI8/NET35_XI0/XI16/XI8/MM6_d
+ N_XI0/XI16/XI8/NET36_XI0/XI16/XI8/MM6_g N_VSS_XI0/XI16/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM7 N_XI0/XI16/XI8/NET36_XI0/XI16/XI8/MM7_d
+ N_XI0/XI16/XI8/NET35_XI0/XI16/XI8/MM7_g N_VSS_XI0/XI16/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM8 N_XI0/XI16/XI8/NET35_XI0/XI16/XI8/MM8_d
+ N_WL<29>_XI0/XI16/XI8/MM8_g N_BLN<7>_XI0/XI16/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI8/MM5 N_XI0/XI16/XI8/NET34_XI0/XI16/XI8/MM5_d
+ N_XI0/XI16/XI8/NET33_XI0/XI16/XI8/MM5_g N_VDD_XI0/XI16/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI8/MM4 N_XI0/XI16/XI8/NET33_XI0/XI16/XI8/MM4_d
+ N_XI0/XI16/XI8/NET34_XI0/XI16/XI8/MM4_g N_VDD_XI0/XI16/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI8/MM10 N_XI0/XI16/XI8/NET35_XI0/XI16/XI8/MM10_d
+ N_XI0/XI16/XI8/NET36_XI0/XI16/XI8/MM10_g N_VDD_XI0/XI16/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI8/MM11 N_XI0/XI16/XI8/NET36_XI0/XI16/XI8/MM11_d
+ N_XI0/XI16/XI8/NET35_XI0/XI16/XI8/MM11_g N_VDD_XI0/XI16/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI9/MM2 N_XI0/XI16/XI9/NET34_XI0/XI16/XI9/MM2_d
+ N_XI0/XI16/XI9/NET33_XI0/XI16/XI9/MM2_g N_VSS_XI0/XI16/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM3 N_XI0/XI16/XI9/NET33_XI0/XI16/XI9/MM3_d
+ N_WL<28>_XI0/XI16/XI9/MM3_g N_BLN<6>_XI0/XI16/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM0 N_XI0/XI16/XI9/NET34_XI0/XI16/XI9/MM0_d
+ N_WL<28>_XI0/XI16/XI9/MM0_g N_BL<6>_XI0/XI16/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM1 N_XI0/XI16/XI9/NET33_XI0/XI16/XI9/MM1_d
+ N_XI0/XI16/XI9/NET34_XI0/XI16/XI9/MM1_g N_VSS_XI0/XI16/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM9 N_XI0/XI16/XI9/NET36_XI0/XI16/XI9/MM9_d
+ N_WL<29>_XI0/XI16/XI9/MM9_g N_BL<6>_XI0/XI16/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM6 N_XI0/XI16/XI9/NET35_XI0/XI16/XI9/MM6_d
+ N_XI0/XI16/XI9/NET36_XI0/XI16/XI9/MM6_g N_VSS_XI0/XI16/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM7 N_XI0/XI16/XI9/NET36_XI0/XI16/XI9/MM7_d
+ N_XI0/XI16/XI9/NET35_XI0/XI16/XI9/MM7_g N_VSS_XI0/XI16/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM8 N_XI0/XI16/XI9/NET35_XI0/XI16/XI9/MM8_d
+ N_WL<29>_XI0/XI16/XI9/MM8_g N_BLN<6>_XI0/XI16/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI9/MM5 N_XI0/XI16/XI9/NET34_XI0/XI16/XI9/MM5_d
+ N_XI0/XI16/XI9/NET33_XI0/XI16/XI9/MM5_g N_VDD_XI0/XI16/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI9/MM4 N_XI0/XI16/XI9/NET33_XI0/XI16/XI9/MM4_d
+ N_XI0/XI16/XI9/NET34_XI0/XI16/XI9/MM4_g N_VDD_XI0/XI16/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI9/MM10 N_XI0/XI16/XI9/NET35_XI0/XI16/XI9/MM10_d
+ N_XI0/XI16/XI9/NET36_XI0/XI16/XI9/MM10_g N_VDD_XI0/XI16/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI9/MM11 N_XI0/XI16/XI9/NET36_XI0/XI16/XI9/MM11_d
+ N_XI0/XI16/XI9/NET35_XI0/XI16/XI9/MM11_g N_VDD_XI0/XI16/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI10/MM2 N_XI0/XI16/XI10/NET34_XI0/XI16/XI10/MM2_d
+ N_XI0/XI16/XI10/NET33_XI0/XI16/XI10/MM2_g N_VSS_XI0/XI16/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM3 N_XI0/XI16/XI10/NET33_XI0/XI16/XI10/MM3_d
+ N_WL<28>_XI0/XI16/XI10/MM3_g N_BLN<5>_XI0/XI16/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM0 N_XI0/XI16/XI10/NET34_XI0/XI16/XI10/MM0_d
+ N_WL<28>_XI0/XI16/XI10/MM0_g N_BL<5>_XI0/XI16/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM1 N_XI0/XI16/XI10/NET33_XI0/XI16/XI10/MM1_d
+ N_XI0/XI16/XI10/NET34_XI0/XI16/XI10/MM1_g N_VSS_XI0/XI16/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM9 N_XI0/XI16/XI10/NET36_XI0/XI16/XI10/MM9_d
+ N_WL<29>_XI0/XI16/XI10/MM9_g N_BL<5>_XI0/XI16/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM6 N_XI0/XI16/XI10/NET35_XI0/XI16/XI10/MM6_d
+ N_XI0/XI16/XI10/NET36_XI0/XI16/XI10/MM6_g N_VSS_XI0/XI16/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM7 N_XI0/XI16/XI10/NET36_XI0/XI16/XI10/MM7_d
+ N_XI0/XI16/XI10/NET35_XI0/XI16/XI10/MM7_g N_VSS_XI0/XI16/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM8 N_XI0/XI16/XI10/NET35_XI0/XI16/XI10/MM8_d
+ N_WL<29>_XI0/XI16/XI10/MM8_g N_BLN<5>_XI0/XI16/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI10/MM5 N_XI0/XI16/XI10/NET34_XI0/XI16/XI10/MM5_d
+ N_XI0/XI16/XI10/NET33_XI0/XI16/XI10/MM5_g N_VDD_XI0/XI16/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI10/MM4 N_XI0/XI16/XI10/NET33_XI0/XI16/XI10/MM4_d
+ N_XI0/XI16/XI10/NET34_XI0/XI16/XI10/MM4_g N_VDD_XI0/XI16/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI10/MM10 N_XI0/XI16/XI10/NET35_XI0/XI16/XI10/MM10_d
+ N_XI0/XI16/XI10/NET36_XI0/XI16/XI10/MM10_g N_VDD_XI0/XI16/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI10/MM11 N_XI0/XI16/XI10/NET36_XI0/XI16/XI10/MM11_d
+ N_XI0/XI16/XI10/NET35_XI0/XI16/XI10/MM11_g N_VDD_XI0/XI16/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI11/MM2 N_XI0/XI16/XI11/NET34_XI0/XI16/XI11/MM2_d
+ N_XI0/XI16/XI11/NET33_XI0/XI16/XI11/MM2_g N_VSS_XI0/XI16/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM3 N_XI0/XI16/XI11/NET33_XI0/XI16/XI11/MM3_d
+ N_WL<28>_XI0/XI16/XI11/MM3_g N_BLN<4>_XI0/XI16/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM0 N_XI0/XI16/XI11/NET34_XI0/XI16/XI11/MM0_d
+ N_WL<28>_XI0/XI16/XI11/MM0_g N_BL<4>_XI0/XI16/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM1 N_XI0/XI16/XI11/NET33_XI0/XI16/XI11/MM1_d
+ N_XI0/XI16/XI11/NET34_XI0/XI16/XI11/MM1_g N_VSS_XI0/XI16/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM9 N_XI0/XI16/XI11/NET36_XI0/XI16/XI11/MM9_d
+ N_WL<29>_XI0/XI16/XI11/MM9_g N_BL<4>_XI0/XI16/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM6 N_XI0/XI16/XI11/NET35_XI0/XI16/XI11/MM6_d
+ N_XI0/XI16/XI11/NET36_XI0/XI16/XI11/MM6_g N_VSS_XI0/XI16/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM7 N_XI0/XI16/XI11/NET36_XI0/XI16/XI11/MM7_d
+ N_XI0/XI16/XI11/NET35_XI0/XI16/XI11/MM7_g N_VSS_XI0/XI16/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM8 N_XI0/XI16/XI11/NET35_XI0/XI16/XI11/MM8_d
+ N_WL<29>_XI0/XI16/XI11/MM8_g N_BLN<4>_XI0/XI16/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI11/MM5 N_XI0/XI16/XI11/NET34_XI0/XI16/XI11/MM5_d
+ N_XI0/XI16/XI11/NET33_XI0/XI16/XI11/MM5_g N_VDD_XI0/XI16/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI11/MM4 N_XI0/XI16/XI11/NET33_XI0/XI16/XI11/MM4_d
+ N_XI0/XI16/XI11/NET34_XI0/XI16/XI11/MM4_g N_VDD_XI0/XI16/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI11/MM10 N_XI0/XI16/XI11/NET35_XI0/XI16/XI11/MM10_d
+ N_XI0/XI16/XI11/NET36_XI0/XI16/XI11/MM10_g N_VDD_XI0/XI16/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI11/MM11 N_XI0/XI16/XI11/NET36_XI0/XI16/XI11/MM11_d
+ N_XI0/XI16/XI11/NET35_XI0/XI16/XI11/MM11_g N_VDD_XI0/XI16/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI12/MM2 N_XI0/XI16/XI12/NET34_XI0/XI16/XI12/MM2_d
+ N_XI0/XI16/XI12/NET33_XI0/XI16/XI12/MM2_g N_VSS_XI0/XI16/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM3 N_XI0/XI16/XI12/NET33_XI0/XI16/XI12/MM3_d
+ N_WL<28>_XI0/XI16/XI12/MM3_g N_BLN<3>_XI0/XI16/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM0 N_XI0/XI16/XI12/NET34_XI0/XI16/XI12/MM0_d
+ N_WL<28>_XI0/XI16/XI12/MM0_g N_BL<3>_XI0/XI16/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM1 N_XI0/XI16/XI12/NET33_XI0/XI16/XI12/MM1_d
+ N_XI0/XI16/XI12/NET34_XI0/XI16/XI12/MM1_g N_VSS_XI0/XI16/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM9 N_XI0/XI16/XI12/NET36_XI0/XI16/XI12/MM9_d
+ N_WL<29>_XI0/XI16/XI12/MM9_g N_BL<3>_XI0/XI16/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM6 N_XI0/XI16/XI12/NET35_XI0/XI16/XI12/MM6_d
+ N_XI0/XI16/XI12/NET36_XI0/XI16/XI12/MM6_g N_VSS_XI0/XI16/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM7 N_XI0/XI16/XI12/NET36_XI0/XI16/XI12/MM7_d
+ N_XI0/XI16/XI12/NET35_XI0/XI16/XI12/MM7_g N_VSS_XI0/XI16/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM8 N_XI0/XI16/XI12/NET35_XI0/XI16/XI12/MM8_d
+ N_WL<29>_XI0/XI16/XI12/MM8_g N_BLN<3>_XI0/XI16/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI12/MM5 N_XI0/XI16/XI12/NET34_XI0/XI16/XI12/MM5_d
+ N_XI0/XI16/XI12/NET33_XI0/XI16/XI12/MM5_g N_VDD_XI0/XI16/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI12/MM4 N_XI0/XI16/XI12/NET33_XI0/XI16/XI12/MM4_d
+ N_XI0/XI16/XI12/NET34_XI0/XI16/XI12/MM4_g N_VDD_XI0/XI16/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI12/MM10 N_XI0/XI16/XI12/NET35_XI0/XI16/XI12/MM10_d
+ N_XI0/XI16/XI12/NET36_XI0/XI16/XI12/MM10_g N_VDD_XI0/XI16/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI12/MM11 N_XI0/XI16/XI12/NET36_XI0/XI16/XI12/MM11_d
+ N_XI0/XI16/XI12/NET35_XI0/XI16/XI12/MM11_g N_VDD_XI0/XI16/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI13/MM2 N_XI0/XI16/XI13/NET34_XI0/XI16/XI13/MM2_d
+ N_XI0/XI16/XI13/NET33_XI0/XI16/XI13/MM2_g N_VSS_XI0/XI16/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM3 N_XI0/XI16/XI13/NET33_XI0/XI16/XI13/MM3_d
+ N_WL<28>_XI0/XI16/XI13/MM3_g N_BLN<2>_XI0/XI16/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM0 N_XI0/XI16/XI13/NET34_XI0/XI16/XI13/MM0_d
+ N_WL<28>_XI0/XI16/XI13/MM0_g N_BL<2>_XI0/XI16/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM1 N_XI0/XI16/XI13/NET33_XI0/XI16/XI13/MM1_d
+ N_XI0/XI16/XI13/NET34_XI0/XI16/XI13/MM1_g N_VSS_XI0/XI16/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM9 N_XI0/XI16/XI13/NET36_XI0/XI16/XI13/MM9_d
+ N_WL<29>_XI0/XI16/XI13/MM9_g N_BL<2>_XI0/XI16/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM6 N_XI0/XI16/XI13/NET35_XI0/XI16/XI13/MM6_d
+ N_XI0/XI16/XI13/NET36_XI0/XI16/XI13/MM6_g N_VSS_XI0/XI16/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM7 N_XI0/XI16/XI13/NET36_XI0/XI16/XI13/MM7_d
+ N_XI0/XI16/XI13/NET35_XI0/XI16/XI13/MM7_g N_VSS_XI0/XI16/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM8 N_XI0/XI16/XI13/NET35_XI0/XI16/XI13/MM8_d
+ N_WL<29>_XI0/XI16/XI13/MM8_g N_BLN<2>_XI0/XI16/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI13/MM5 N_XI0/XI16/XI13/NET34_XI0/XI16/XI13/MM5_d
+ N_XI0/XI16/XI13/NET33_XI0/XI16/XI13/MM5_g N_VDD_XI0/XI16/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI13/MM4 N_XI0/XI16/XI13/NET33_XI0/XI16/XI13/MM4_d
+ N_XI0/XI16/XI13/NET34_XI0/XI16/XI13/MM4_g N_VDD_XI0/XI16/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI13/MM10 N_XI0/XI16/XI13/NET35_XI0/XI16/XI13/MM10_d
+ N_XI0/XI16/XI13/NET36_XI0/XI16/XI13/MM10_g N_VDD_XI0/XI16/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI13/MM11 N_XI0/XI16/XI13/NET36_XI0/XI16/XI13/MM11_d
+ N_XI0/XI16/XI13/NET35_XI0/XI16/XI13/MM11_g N_VDD_XI0/XI16/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI14/MM2 N_XI0/XI16/XI14/NET34_XI0/XI16/XI14/MM2_d
+ N_XI0/XI16/XI14/NET33_XI0/XI16/XI14/MM2_g N_VSS_XI0/XI16/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM3 N_XI0/XI16/XI14/NET33_XI0/XI16/XI14/MM3_d
+ N_WL<28>_XI0/XI16/XI14/MM3_g N_BLN<1>_XI0/XI16/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM0 N_XI0/XI16/XI14/NET34_XI0/XI16/XI14/MM0_d
+ N_WL<28>_XI0/XI16/XI14/MM0_g N_BL<1>_XI0/XI16/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM1 N_XI0/XI16/XI14/NET33_XI0/XI16/XI14/MM1_d
+ N_XI0/XI16/XI14/NET34_XI0/XI16/XI14/MM1_g N_VSS_XI0/XI16/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM9 N_XI0/XI16/XI14/NET36_XI0/XI16/XI14/MM9_d
+ N_WL<29>_XI0/XI16/XI14/MM9_g N_BL<1>_XI0/XI16/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM6 N_XI0/XI16/XI14/NET35_XI0/XI16/XI14/MM6_d
+ N_XI0/XI16/XI14/NET36_XI0/XI16/XI14/MM6_g N_VSS_XI0/XI16/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM7 N_XI0/XI16/XI14/NET36_XI0/XI16/XI14/MM7_d
+ N_XI0/XI16/XI14/NET35_XI0/XI16/XI14/MM7_g N_VSS_XI0/XI16/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM8 N_XI0/XI16/XI14/NET35_XI0/XI16/XI14/MM8_d
+ N_WL<29>_XI0/XI16/XI14/MM8_g N_BLN<1>_XI0/XI16/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI14/MM5 N_XI0/XI16/XI14/NET34_XI0/XI16/XI14/MM5_d
+ N_XI0/XI16/XI14/NET33_XI0/XI16/XI14/MM5_g N_VDD_XI0/XI16/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI14/MM4 N_XI0/XI16/XI14/NET33_XI0/XI16/XI14/MM4_d
+ N_XI0/XI16/XI14/NET34_XI0/XI16/XI14/MM4_g N_VDD_XI0/XI16/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI14/MM10 N_XI0/XI16/XI14/NET35_XI0/XI16/XI14/MM10_d
+ N_XI0/XI16/XI14/NET36_XI0/XI16/XI14/MM10_g N_VDD_XI0/XI16/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI14/MM11 N_XI0/XI16/XI14/NET36_XI0/XI16/XI14/MM11_d
+ N_XI0/XI16/XI14/NET35_XI0/XI16/XI14/MM11_g N_VDD_XI0/XI16/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI15/MM2 N_XI0/XI16/XI15/NET34_XI0/XI16/XI15/MM2_d
+ N_XI0/XI16/XI15/NET33_XI0/XI16/XI15/MM2_g N_VSS_XI0/XI16/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM3 N_XI0/XI16/XI15/NET33_XI0/XI16/XI15/MM3_d
+ N_WL<28>_XI0/XI16/XI15/MM3_g N_BLN<0>_XI0/XI16/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM0 N_XI0/XI16/XI15/NET34_XI0/XI16/XI15/MM0_d
+ N_WL<28>_XI0/XI16/XI15/MM0_g N_BL<0>_XI0/XI16/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM1 N_XI0/XI16/XI15/NET33_XI0/XI16/XI15/MM1_d
+ N_XI0/XI16/XI15/NET34_XI0/XI16/XI15/MM1_g N_VSS_XI0/XI16/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM9 N_XI0/XI16/XI15/NET36_XI0/XI16/XI15/MM9_d
+ N_WL<29>_XI0/XI16/XI15/MM9_g N_BL<0>_XI0/XI16/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM6 N_XI0/XI16/XI15/NET35_XI0/XI16/XI15/MM6_d
+ N_XI0/XI16/XI15/NET36_XI0/XI16/XI15/MM6_g N_VSS_XI0/XI16/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM7 N_XI0/XI16/XI15/NET36_XI0/XI16/XI15/MM7_d
+ N_XI0/XI16/XI15/NET35_XI0/XI16/XI15/MM7_g N_VSS_XI0/XI16/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM8 N_XI0/XI16/XI15/NET35_XI0/XI16/XI15/MM8_d
+ N_WL<29>_XI0/XI16/XI15/MM8_g N_BLN<0>_XI0/XI16/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI16/XI15/MM5 N_XI0/XI16/XI15/NET34_XI0/XI16/XI15/MM5_d
+ N_XI0/XI16/XI15/NET33_XI0/XI16/XI15/MM5_g N_VDD_XI0/XI16/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI15/MM4 N_XI0/XI16/XI15/NET33_XI0/XI16/XI15/MM4_d
+ N_XI0/XI16/XI15/NET34_XI0/XI16/XI15/MM4_g N_VDD_XI0/XI16/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI15/MM10 N_XI0/XI16/XI15/NET35_XI0/XI16/XI15/MM10_d
+ N_XI0/XI16/XI15/NET36_XI0/XI16/XI15/MM10_g N_VDD_XI0/XI16/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI16/XI15/MM11 N_XI0/XI16/XI15/NET36_XI0/XI16/XI15/MM11_d
+ N_XI0/XI16/XI15/NET35_XI0/XI16/XI15/MM11_g N_VDD_XI0/XI16/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI0/MM2 N_XI0/XI17/XI0/NET34_XI0/XI17/XI0/MM2_d
+ N_XI0/XI17/XI0/NET33_XI0/XI17/XI0/MM2_g N_VSS_XI0/XI17/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM3 N_XI0/XI17/XI0/NET33_XI0/XI17/XI0/MM3_d
+ N_WL<30>_XI0/XI17/XI0/MM3_g N_BLN<15>_XI0/XI17/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM0 N_XI0/XI17/XI0/NET34_XI0/XI17/XI0/MM0_d
+ N_WL<30>_XI0/XI17/XI0/MM0_g N_BL<15>_XI0/XI17/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM1 N_XI0/XI17/XI0/NET33_XI0/XI17/XI0/MM1_d
+ N_XI0/XI17/XI0/NET34_XI0/XI17/XI0/MM1_g N_VSS_XI0/XI17/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM9 N_XI0/XI17/XI0/NET36_XI0/XI17/XI0/MM9_d
+ N_WL<31>_XI0/XI17/XI0/MM9_g N_BL<15>_XI0/XI17/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM6 N_XI0/XI17/XI0/NET35_XI0/XI17/XI0/MM6_d
+ N_XI0/XI17/XI0/NET36_XI0/XI17/XI0/MM6_g N_VSS_XI0/XI17/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM7 N_XI0/XI17/XI0/NET36_XI0/XI17/XI0/MM7_d
+ N_XI0/XI17/XI0/NET35_XI0/XI17/XI0/MM7_g N_VSS_XI0/XI17/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM8 N_XI0/XI17/XI0/NET35_XI0/XI17/XI0/MM8_d
+ N_WL<31>_XI0/XI17/XI0/MM8_g N_BLN<15>_XI0/XI17/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI0/MM5 N_XI0/XI17/XI0/NET34_XI0/XI17/XI0/MM5_d
+ N_XI0/XI17/XI0/NET33_XI0/XI17/XI0/MM5_g N_VDD_XI0/XI17/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI0/MM4 N_XI0/XI17/XI0/NET33_XI0/XI17/XI0/MM4_d
+ N_XI0/XI17/XI0/NET34_XI0/XI17/XI0/MM4_g N_VDD_XI0/XI17/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI0/MM10 N_XI0/XI17/XI0/NET35_XI0/XI17/XI0/MM10_d
+ N_XI0/XI17/XI0/NET36_XI0/XI17/XI0/MM10_g N_VDD_XI0/XI17/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI0/MM11 N_XI0/XI17/XI0/NET36_XI0/XI17/XI0/MM11_d
+ N_XI0/XI17/XI0/NET35_XI0/XI17/XI0/MM11_g N_VDD_XI0/XI17/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI1/MM2 N_XI0/XI17/XI1/NET34_XI0/XI17/XI1/MM2_d
+ N_XI0/XI17/XI1/NET33_XI0/XI17/XI1/MM2_g N_VSS_XI0/XI17/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM3 N_XI0/XI17/XI1/NET33_XI0/XI17/XI1/MM3_d
+ N_WL<30>_XI0/XI17/XI1/MM3_g N_BLN<14>_XI0/XI17/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM0 N_XI0/XI17/XI1/NET34_XI0/XI17/XI1/MM0_d
+ N_WL<30>_XI0/XI17/XI1/MM0_g N_BL<14>_XI0/XI17/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM1 N_XI0/XI17/XI1/NET33_XI0/XI17/XI1/MM1_d
+ N_XI0/XI17/XI1/NET34_XI0/XI17/XI1/MM1_g N_VSS_XI0/XI17/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM9 N_XI0/XI17/XI1/NET36_XI0/XI17/XI1/MM9_d
+ N_WL<31>_XI0/XI17/XI1/MM9_g N_BL<14>_XI0/XI17/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM6 N_XI0/XI17/XI1/NET35_XI0/XI17/XI1/MM6_d
+ N_XI0/XI17/XI1/NET36_XI0/XI17/XI1/MM6_g N_VSS_XI0/XI17/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM7 N_XI0/XI17/XI1/NET36_XI0/XI17/XI1/MM7_d
+ N_XI0/XI17/XI1/NET35_XI0/XI17/XI1/MM7_g N_VSS_XI0/XI17/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM8 N_XI0/XI17/XI1/NET35_XI0/XI17/XI1/MM8_d
+ N_WL<31>_XI0/XI17/XI1/MM8_g N_BLN<14>_XI0/XI17/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI1/MM5 N_XI0/XI17/XI1/NET34_XI0/XI17/XI1/MM5_d
+ N_XI0/XI17/XI1/NET33_XI0/XI17/XI1/MM5_g N_VDD_XI0/XI17/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI1/MM4 N_XI0/XI17/XI1/NET33_XI0/XI17/XI1/MM4_d
+ N_XI0/XI17/XI1/NET34_XI0/XI17/XI1/MM4_g N_VDD_XI0/XI17/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI1/MM10 N_XI0/XI17/XI1/NET35_XI0/XI17/XI1/MM10_d
+ N_XI0/XI17/XI1/NET36_XI0/XI17/XI1/MM10_g N_VDD_XI0/XI17/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI1/MM11 N_XI0/XI17/XI1/NET36_XI0/XI17/XI1/MM11_d
+ N_XI0/XI17/XI1/NET35_XI0/XI17/XI1/MM11_g N_VDD_XI0/XI17/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI2/MM2 N_XI0/XI17/XI2/NET34_XI0/XI17/XI2/MM2_d
+ N_XI0/XI17/XI2/NET33_XI0/XI17/XI2/MM2_g N_VSS_XI0/XI17/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM3 N_XI0/XI17/XI2/NET33_XI0/XI17/XI2/MM3_d
+ N_WL<30>_XI0/XI17/XI2/MM3_g N_BLN<13>_XI0/XI17/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM0 N_XI0/XI17/XI2/NET34_XI0/XI17/XI2/MM0_d
+ N_WL<30>_XI0/XI17/XI2/MM0_g N_BL<13>_XI0/XI17/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM1 N_XI0/XI17/XI2/NET33_XI0/XI17/XI2/MM1_d
+ N_XI0/XI17/XI2/NET34_XI0/XI17/XI2/MM1_g N_VSS_XI0/XI17/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM9 N_XI0/XI17/XI2/NET36_XI0/XI17/XI2/MM9_d
+ N_WL<31>_XI0/XI17/XI2/MM9_g N_BL<13>_XI0/XI17/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM6 N_XI0/XI17/XI2/NET35_XI0/XI17/XI2/MM6_d
+ N_XI0/XI17/XI2/NET36_XI0/XI17/XI2/MM6_g N_VSS_XI0/XI17/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM7 N_XI0/XI17/XI2/NET36_XI0/XI17/XI2/MM7_d
+ N_XI0/XI17/XI2/NET35_XI0/XI17/XI2/MM7_g N_VSS_XI0/XI17/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM8 N_XI0/XI17/XI2/NET35_XI0/XI17/XI2/MM8_d
+ N_WL<31>_XI0/XI17/XI2/MM8_g N_BLN<13>_XI0/XI17/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI2/MM5 N_XI0/XI17/XI2/NET34_XI0/XI17/XI2/MM5_d
+ N_XI0/XI17/XI2/NET33_XI0/XI17/XI2/MM5_g N_VDD_XI0/XI17/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI2/MM4 N_XI0/XI17/XI2/NET33_XI0/XI17/XI2/MM4_d
+ N_XI0/XI17/XI2/NET34_XI0/XI17/XI2/MM4_g N_VDD_XI0/XI17/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI2/MM10 N_XI0/XI17/XI2/NET35_XI0/XI17/XI2/MM10_d
+ N_XI0/XI17/XI2/NET36_XI0/XI17/XI2/MM10_g N_VDD_XI0/XI17/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI2/MM11 N_XI0/XI17/XI2/NET36_XI0/XI17/XI2/MM11_d
+ N_XI0/XI17/XI2/NET35_XI0/XI17/XI2/MM11_g N_VDD_XI0/XI17/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI3/MM2 N_XI0/XI17/XI3/NET34_XI0/XI17/XI3/MM2_d
+ N_XI0/XI17/XI3/NET33_XI0/XI17/XI3/MM2_g N_VSS_XI0/XI17/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM3 N_XI0/XI17/XI3/NET33_XI0/XI17/XI3/MM3_d
+ N_WL<30>_XI0/XI17/XI3/MM3_g N_BLN<12>_XI0/XI17/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM0 N_XI0/XI17/XI3/NET34_XI0/XI17/XI3/MM0_d
+ N_WL<30>_XI0/XI17/XI3/MM0_g N_BL<12>_XI0/XI17/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM1 N_XI0/XI17/XI3/NET33_XI0/XI17/XI3/MM1_d
+ N_XI0/XI17/XI3/NET34_XI0/XI17/XI3/MM1_g N_VSS_XI0/XI17/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM9 N_XI0/XI17/XI3/NET36_XI0/XI17/XI3/MM9_d
+ N_WL<31>_XI0/XI17/XI3/MM9_g N_BL<12>_XI0/XI17/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM6 N_XI0/XI17/XI3/NET35_XI0/XI17/XI3/MM6_d
+ N_XI0/XI17/XI3/NET36_XI0/XI17/XI3/MM6_g N_VSS_XI0/XI17/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM7 N_XI0/XI17/XI3/NET36_XI0/XI17/XI3/MM7_d
+ N_XI0/XI17/XI3/NET35_XI0/XI17/XI3/MM7_g N_VSS_XI0/XI17/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM8 N_XI0/XI17/XI3/NET35_XI0/XI17/XI3/MM8_d
+ N_WL<31>_XI0/XI17/XI3/MM8_g N_BLN<12>_XI0/XI17/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI3/MM5 N_XI0/XI17/XI3/NET34_XI0/XI17/XI3/MM5_d
+ N_XI0/XI17/XI3/NET33_XI0/XI17/XI3/MM5_g N_VDD_XI0/XI17/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI3/MM4 N_XI0/XI17/XI3/NET33_XI0/XI17/XI3/MM4_d
+ N_XI0/XI17/XI3/NET34_XI0/XI17/XI3/MM4_g N_VDD_XI0/XI17/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI3/MM10 N_XI0/XI17/XI3/NET35_XI0/XI17/XI3/MM10_d
+ N_XI0/XI17/XI3/NET36_XI0/XI17/XI3/MM10_g N_VDD_XI0/XI17/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI3/MM11 N_XI0/XI17/XI3/NET36_XI0/XI17/XI3/MM11_d
+ N_XI0/XI17/XI3/NET35_XI0/XI17/XI3/MM11_g N_VDD_XI0/XI17/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI4/MM2 N_XI0/XI17/XI4/NET34_XI0/XI17/XI4/MM2_d
+ N_XI0/XI17/XI4/NET33_XI0/XI17/XI4/MM2_g N_VSS_XI0/XI17/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM3 N_XI0/XI17/XI4/NET33_XI0/XI17/XI4/MM3_d
+ N_WL<30>_XI0/XI17/XI4/MM3_g N_BLN<11>_XI0/XI17/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM0 N_XI0/XI17/XI4/NET34_XI0/XI17/XI4/MM0_d
+ N_WL<30>_XI0/XI17/XI4/MM0_g N_BL<11>_XI0/XI17/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM1 N_XI0/XI17/XI4/NET33_XI0/XI17/XI4/MM1_d
+ N_XI0/XI17/XI4/NET34_XI0/XI17/XI4/MM1_g N_VSS_XI0/XI17/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM9 N_XI0/XI17/XI4/NET36_XI0/XI17/XI4/MM9_d
+ N_WL<31>_XI0/XI17/XI4/MM9_g N_BL<11>_XI0/XI17/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM6 N_XI0/XI17/XI4/NET35_XI0/XI17/XI4/MM6_d
+ N_XI0/XI17/XI4/NET36_XI0/XI17/XI4/MM6_g N_VSS_XI0/XI17/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM7 N_XI0/XI17/XI4/NET36_XI0/XI17/XI4/MM7_d
+ N_XI0/XI17/XI4/NET35_XI0/XI17/XI4/MM7_g N_VSS_XI0/XI17/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM8 N_XI0/XI17/XI4/NET35_XI0/XI17/XI4/MM8_d
+ N_WL<31>_XI0/XI17/XI4/MM8_g N_BLN<11>_XI0/XI17/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI4/MM5 N_XI0/XI17/XI4/NET34_XI0/XI17/XI4/MM5_d
+ N_XI0/XI17/XI4/NET33_XI0/XI17/XI4/MM5_g N_VDD_XI0/XI17/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI4/MM4 N_XI0/XI17/XI4/NET33_XI0/XI17/XI4/MM4_d
+ N_XI0/XI17/XI4/NET34_XI0/XI17/XI4/MM4_g N_VDD_XI0/XI17/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI4/MM10 N_XI0/XI17/XI4/NET35_XI0/XI17/XI4/MM10_d
+ N_XI0/XI17/XI4/NET36_XI0/XI17/XI4/MM10_g N_VDD_XI0/XI17/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI4/MM11 N_XI0/XI17/XI4/NET36_XI0/XI17/XI4/MM11_d
+ N_XI0/XI17/XI4/NET35_XI0/XI17/XI4/MM11_g N_VDD_XI0/XI17/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI5/MM2 N_XI0/XI17/XI5/NET34_XI0/XI17/XI5/MM2_d
+ N_XI0/XI17/XI5/NET33_XI0/XI17/XI5/MM2_g N_VSS_XI0/XI17/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM3 N_XI0/XI17/XI5/NET33_XI0/XI17/XI5/MM3_d
+ N_WL<30>_XI0/XI17/XI5/MM3_g N_BLN<10>_XI0/XI17/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM0 N_XI0/XI17/XI5/NET34_XI0/XI17/XI5/MM0_d
+ N_WL<30>_XI0/XI17/XI5/MM0_g N_BL<10>_XI0/XI17/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM1 N_XI0/XI17/XI5/NET33_XI0/XI17/XI5/MM1_d
+ N_XI0/XI17/XI5/NET34_XI0/XI17/XI5/MM1_g N_VSS_XI0/XI17/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM9 N_XI0/XI17/XI5/NET36_XI0/XI17/XI5/MM9_d
+ N_WL<31>_XI0/XI17/XI5/MM9_g N_BL<10>_XI0/XI17/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM6 N_XI0/XI17/XI5/NET35_XI0/XI17/XI5/MM6_d
+ N_XI0/XI17/XI5/NET36_XI0/XI17/XI5/MM6_g N_VSS_XI0/XI17/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM7 N_XI0/XI17/XI5/NET36_XI0/XI17/XI5/MM7_d
+ N_XI0/XI17/XI5/NET35_XI0/XI17/XI5/MM7_g N_VSS_XI0/XI17/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM8 N_XI0/XI17/XI5/NET35_XI0/XI17/XI5/MM8_d
+ N_WL<31>_XI0/XI17/XI5/MM8_g N_BLN<10>_XI0/XI17/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI5/MM5 N_XI0/XI17/XI5/NET34_XI0/XI17/XI5/MM5_d
+ N_XI0/XI17/XI5/NET33_XI0/XI17/XI5/MM5_g N_VDD_XI0/XI17/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI5/MM4 N_XI0/XI17/XI5/NET33_XI0/XI17/XI5/MM4_d
+ N_XI0/XI17/XI5/NET34_XI0/XI17/XI5/MM4_g N_VDD_XI0/XI17/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI5/MM10 N_XI0/XI17/XI5/NET35_XI0/XI17/XI5/MM10_d
+ N_XI0/XI17/XI5/NET36_XI0/XI17/XI5/MM10_g N_VDD_XI0/XI17/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI5/MM11 N_XI0/XI17/XI5/NET36_XI0/XI17/XI5/MM11_d
+ N_XI0/XI17/XI5/NET35_XI0/XI17/XI5/MM11_g N_VDD_XI0/XI17/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI6/MM2 N_XI0/XI17/XI6/NET34_XI0/XI17/XI6/MM2_d
+ N_XI0/XI17/XI6/NET33_XI0/XI17/XI6/MM2_g N_VSS_XI0/XI17/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM3 N_XI0/XI17/XI6/NET33_XI0/XI17/XI6/MM3_d
+ N_WL<30>_XI0/XI17/XI6/MM3_g N_BLN<9>_XI0/XI17/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM0 N_XI0/XI17/XI6/NET34_XI0/XI17/XI6/MM0_d
+ N_WL<30>_XI0/XI17/XI6/MM0_g N_BL<9>_XI0/XI17/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM1 N_XI0/XI17/XI6/NET33_XI0/XI17/XI6/MM1_d
+ N_XI0/XI17/XI6/NET34_XI0/XI17/XI6/MM1_g N_VSS_XI0/XI17/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM9 N_XI0/XI17/XI6/NET36_XI0/XI17/XI6/MM9_d
+ N_WL<31>_XI0/XI17/XI6/MM9_g N_BL<9>_XI0/XI17/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM6 N_XI0/XI17/XI6/NET35_XI0/XI17/XI6/MM6_d
+ N_XI0/XI17/XI6/NET36_XI0/XI17/XI6/MM6_g N_VSS_XI0/XI17/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM7 N_XI0/XI17/XI6/NET36_XI0/XI17/XI6/MM7_d
+ N_XI0/XI17/XI6/NET35_XI0/XI17/XI6/MM7_g N_VSS_XI0/XI17/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM8 N_XI0/XI17/XI6/NET35_XI0/XI17/XI6/MM8_d
+ N_WL<31>_XI0/XI17/XI6/MM8_g N_BLN<9>_XI0/XI17/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI6/MM5 N_XI0/XI17/XI6/NET34_XI0/XI17/XI6/MM5_d
+ N_XI0/XI17/XI6/NET33_XI0/XI17/XI6/MM5_g N_VDD_XI0/XI17/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI6/MM4 N_XI0/XI17/XI6/NET33_XI0/XI17/XI6/MM4_d
+ N_XI0/XI17/XI6/NET34_XI0/XI17/XI6/MM4_g N_VDD_XI0/XI17/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI6/MM10 N_XI0/XI17/XI6/NET35_XI0/XI17/XI6/MM10_d
+ N_XI0/XI17/XI6/NET36_XI0/XI17/XI6/MM10_g N_VDD_XI0/XI17/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI6/MM11 N_XI0/XI17/XI6/NET36_XI0/XI17/XI6/MM11_d
+ N_XI0/XI17/XI6/NET35_XI0/XI17/XI6/MM11_g N_VDD_XI0/XI17/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI7/MM2 N_XI0/XI17/XI7/NET34_XI0/XI17/XI7/MM2_d
+ N_XI0/XI17/XI7/NET33_XI0/XI17/XI7/MM2_g N_VSS_XI0/XI17/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM3 N_XI0/XI17/XI7/NET33_XI0/XI17/XI7/MM3_d
+ N_WL<30>_XI0/XI17/XI7/MM3_g N_BLN<8>_XI0/XI17/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM0 N_XI0/XI17/XI7/NET34_XI0/XI17/XI7/MM0_d
+ N_WL<30>_XI0/XI17/XI7/MM0_g N_BL<8>_XI0/XI17/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM1 N_XI0/XI17/XI7/NET33_XI0/XI17/XI7/MM1_d
+ N_XI0/XI17/XI7/NET34_XI0/XI17/XI7/MM1_g N_VSS_XI0/XI17/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM9 N_XI0/XI17/XI7/NET36_XI0/XI17/XI7/MM9_d
+ N_WL<31>_XI0/XI17/XI7/MM9_g N_BL<8>_XI0/XI17/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM6 N_XI0/XI17/XI7/NET35_XI0/XI17/XI7/MM6_d
+ N_XI0/XI17/XI7/NET36_XI0/XI17/XI7/MM6_g N_VSS_XI0/XI17/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM7 N_XI0/XI17/XI7/NET36_XI0/XI17/XI7/MM7_d
+ N_XI0/XI17/XI7/NET35_XI0/XI17/XI7/MM7_g N_VSS_XI0/XI17/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM8 N_XI0/XI17/XI7/NET35_XI0/XI17/XI7/MM8_d
+ N_WL<31>_XI0/XI17/XI7/MM8_g N_BLN<8>_XI0/XI17/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI7/MM5 N_XI0/XI17/XI7/NET34_XI0/XI17/XI7/MM5_d
+ N_XI0/XI17/XI7/NET33_XI0/XI17/XI7/MM5_g N_VDD_XI0/XI17/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI7/MM4 N_XI0/XI17/XI7/NET33_XI0/XI17/XI7/MM4_d
+ N_XI0/XI17/XI7/NET34_XI0/XI17/XI7/MM4_g N_VDD_XI0/XI17/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI7/MM10 N_XI0/XI17/XI7/NET35_XI0/XI17/XI7/MM10_d
+ N_XI0/XI17/XI7/NET36_XI0/XI17/XI7/MM10_g N_VDD_XI0/XI17/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI7/MM11 N_XI0/XI17/XI7/NET36_XI0/XI17/XI7/MM11_d
+ N_XI0/XI17/XI7/NET35_XI0/XI17/XI7/MM11_g N_VDD_XI0/XI17/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI8/MM2 N_XI0/XI17/XI8/NET34_XI0/XI17/XI8/MM2_d
+ N_XI0/XI17/XI8/NET33_XI0/XI17/XI8/MM2_g N_VSS_XI0/XI17/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM3 N_XI0/XI17/XI8/NET33_XI0/XI17/XI8/MM3_d
+ N_WL<30>_XI0/XI17/XI8/MM3_g N_BLN<7>_XI0/XI17/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM0 N_XI0/XI17/XI8/NET34_XI0/XI17/XI8/MM0_d
+ N_WL<30>_XI0/XI17/XI8/MM0_g N_BL<7>_XI0/XI17/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM1 N_XI0/XI17/XI8/NET33_XI0/XI17/XI8/MM1_d
+ N_XI0/XI17/XI8/NET34_XI0/XI17/XI8/MM1_g N_VSS_XI0/XI17/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM9 N_XI0/XI17/XI8/NET36_XI0/XI17/XI8/MM9_d
+ N_WL<31>_XI0/XI17/XI8/MM9_g N_BL<7>_XI0/XI17/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM6 N_XI0/XI17/XI8/NET35_XI0/XI17/XI8/MM6_d
+ N_XI0/XI17/XI8/NET36_XI0/XI17/XI8/MM6_g N_VSS_XI0/XI17/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM7 N_XI0/XI17/XI8/NET36_XI0/XI17/XI8/MM7_d
+ N_XI0/XI17/XI8/NET35_XI0/XI17/XI8/MM7_g N_VSS_XI0/XI17/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM8 N_XI0/XI17/XI8/NET35_XI0/XI17/XI8/MM8_d
+ N_WL<31>_XI0/XI17/XI8/MM8_g N_BLN<7>_XI0/XI17/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI8/MM5 N_XI0/XI17/XI8/NET34_XI0/XI17/XI8/MM5_d
+ N_XI0/XI17/XI8/NET33_XI0/XI17/XI8/MM5_g N_VDD_XI0/XI17/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI8/MM4 N_XI0/XI17/XI8/NET33_XI0/XI17/XI8/MM4_d
+ N_XI0/XI17/XI8/NET34_XI0/XI17/XI8/MM4_g N_VDD_XI0/XI17/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI8/MM10 N_XI0/XI17/XI8/NET35_XI0/XI17/XI8/MM10_d
+ N_XI0/XI17/XI8/NET36_XI0/XI17/XI8/MM10_g N_VDD_XI0/XI17/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI8/MM11 N_XI0/XI17/XI8/NET36_XI0/XI17/XI8/MM11_d
+ N_XI0/XI17/XI8/NET35_XI0/XI17/XI8/MM11_g N_VDD_XI0/XI17/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI9/MM2 N_XI0/XI17/XI9/NET34_XI0/XI17/XI9/MM2_d
+ N_XI0/XI17/XI9/NET33_XI0/XI17/XI9/MM2_g N_VSS_XI0/XI17/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM3 N_XI0/XI17/XI9/NET33_XI0/XI17/XI9/MM3_d
+ N_WL<30>_XI0/XI17/XI9/MM3_g N_BLN<6>_XI0/XI17/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM0 N_XI0/XI17/XI9/NET34_XI0/XI17/XI9/MM0_d
+ N_WL<30>_XI0/XI17/XI9/MM0_g N_BL<6>_XI0/XI17/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM1 N_XI0/XI17/XI9/NET33_XI0/XI17/XI9/MM1_d
+ N_XI0/XI17/XI9/NET34_XI0/XI17/XI9/MM1_g N_VSS_XI0/XI17/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM9 N_XI0/XI17/XI9/NET36_XI0/XI17/XI9/MM9_d
+ N_WL<31>_XI0/XI17/XI9/MM9_g N_BL<6>_XI0/XI17/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM6 N_XI0/XI17/XI9/NET35_XI0/XI17/XI9/MM6_d
+ N_XI0/XI17/XI9/NET36_XI0/XI17/XI9/MM6_g N_VSS_XI0/XI17/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM7 N_XI0/XI17/XI9/NET36_XI0/XI17/XI9/MM7_d
+ N_XI0/XI17/XI9/NET35_XI0/XI17/XI9/MM7_g N_VSS_XI0/XI17/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM8 N_XI0/XI17/XI9/NET35_XI0/XI17/XI9/MM8_d
+ N_WL<31>_XI0/XI17/XI9/MM8_g N_BLN<6>_XI0/XI17/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI9/MM5 N_XI0/XI17/XI9/NET34_XI0/XI17/XI9/MM5_d
+ N_XI0/XI17/XI9/NET33_XI0/XI17/XI9/MM5_g N_VDD_XI0/XI17/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI9/MM4 N_XI0/XI17/XI9/NET33_XI0/XI17/XI9/MM4_d
+ N_XI0/XI17/XI9/NET34_XI0/XI17/XI9/MM4_g N_VDD_XI0/XI17/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI9/MM10 N_XI0/XI17/XI9/NET35_XI0/XI17/XI9/MM10_d
+ N_XI0/XI17/XI9/NET36_XI0/XI17/XI9/MM10_g N_VDD_XI0/XI17/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI9/MM11 N_XI0/XI17/XI9/NET36_XI0/XI17/XI9/MM11_d
+ N_XI0/XI17/XI9/NET35_XI0/XI17/XI9/MM11_g N_VDD_XI0/XI17/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI10/MM2 N_XI0/XI17/XI10/NET34_XI0/XI17/XI10/MM2_d
+ N_XI0/XI17/XI10/NET33_XI0/XI17/XI10/MM2_g N_VSS_XI0/XI17/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM3 N_XI0/XI17/XI10/NET33_XI0/XI17/XI10/MM3_d
+ N_WL<30>_XI0/XI17/XI10/MM3_g N_BLN<5>_XI0/XI17/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM0 N_XI0/XI17/XI10/NET34_XI0/XI17/XI10/MM0_d
+ N_WL<30>_XI0/XI17/XI10/MM0_g N_BL<5>_XI0/XI17/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM1 N_XI0/XI17/XI10/NET33_XI0/XI17/XI10/MM1_d
+ N_XI0/XI17/XI10/NET34_XI0/XI17/XI10/MM1_g N_VSS_XI0/XI17/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM9 N_XI0/XI17/XI10/NET36_XI0/XI17/XI10/MM9_d
+ N_WL<31>_XI0/XI17/XI10/MM9_g N_BL<5>_XI0/XI17/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM6 N_XI0/XI17/XI10/NET35_XI0/XI17/XI10/MM6_d
+ N_XI0/XI17/XI10/NET36_XI0/XI17/XI10/MM6_g N_VSS_XI0/XI17/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM7 N_XI0/XI17/XI10/NET36_XI0/XI17/XI10/MM7_d
+ N_XI0/XI17/XI10/NET35_XI0/XI17/XI10/MM7_g N_VSS_XI0/XI17/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM8 N_XI0/XI17/XI10/NET35_XI0/XI17/XI10/MM8_d
+ N_WL<31>_XI0/XI17/XI10/MM8_g N_BLN<5>_XI0/XI17/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI10/MM5 N_XI0/XI17/XI10/NET34_XI0/XI17/XI10/MM5_d
+ N_XI0/XI17/XI10/NET33_XI0/XI17/XI10/MM5_g N_VDD_XI0/XI17/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI10/MM4 N_XI0/XI17/XI10/NET33_XI0/XI17/XI10/MM4_d
+ N_XI0/XI17/XI10/NET34_XI0/XI17/XI10/MM4_g N_VDD_XI0/XI17/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI10/MM10 N_XI0/XI17/XI10/NET35_XI0/XI17/XI10/MM10_d
+ N_XI0/XI17/XI10/NET36_XI0/XI17/XI10/MM10_g N_VDD_XI0/XI17/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI10/MM11 N_XI0/XI17/XI10/NET36_XI0/XI17/XI10/MM11_d
+ N_XI0/XI17/XI10/NET35_XI0/XI17/XI10/MM11_g N_VDD_XI0/XI17/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI11/MM2 N_XI0/XI17/XI11/NET34_XI0/XI17/XI11/MM2_d
+ N_XI0/XI17/XI11/NET33_XI0/XI17/XI11/MM2_g N_VSS_XI0/XI17/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM3 N_XI0/XI17/XI11/NET33_XI0/XI17/XI11/MM3_d
+ N_WL<30>_XI0/XI17/XI11/MM3_g N_BLN<4>_XI0/XI17/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM0 N_XI0/XI17/XI11/NET34_XI0/XI17/XI11/MM0_d
+ N_WL<30>_XI0/XI17/XI11/MM0_g N_BL<4>_XI0/XI17/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM1 N_XI0/XI17/XI11/NET33_XI0/XI17/XI11/MM1_d
+ N_XI0/XI17/XI11/NET34_XI0/XI17/XI11/MM1_g N_VSS_XI0/XI17/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM9 N_XI0/XI17/XI11/NET36_XI0/XI17/XI11/MM9_d
+ N_WL<31>_XI0/XI17/XI11/MM9_g N_BL<4>_XI0/XI17/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM6 N_XI0/XI17/XI11/NET35_XI0/XI17/XI11/MM6_d
+ N_XI0/XI17/XI11/NET36_XI0/XI17/XI11/MM6_g N_VSS_XI0/XI17/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM7 N_XI0/XI17/XI11/NET36_XI0/XI17/XI11/MM7_d
+ N_XI0/XI17/XI11/NET35_XI0/XI17/XI11/MM7_g N_VSS_XI0/XI17/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM8 N_XI0/XI17/XI11/NET35_XI0/XI17/XI11/MM8_d
+ N_WL<31>_XI0/XI17/XI11/MM8_g N_BLN<4>_XI0/XI17/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI11/MM5 N_XI0/XI17/XI11/NET34_XI0/XI17/XI11/MM5_d
+ N_XI0/XI17/XI11/NET33_XI0/XI17/XI11/MM5_g N_VDD_XI0/XI17/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI11/MM4 N_XI0/XI17/XI11/NET33_XI0/XI17/XI11/MM4_d
+ N_XI0/XI17/XI11/NET34_XI0/XI17/XI11/MM4_g N_VDD_XI0/XI17/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI11/MM10 N_XI0/XI17/XI11/NET35_XI0/XI17/XI11/MM10_d
+ N_XI0/XI17/XI11/NET36_XI0/XI17/XI11/MM10_g N_VDD_XI0/XI17/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI11/MM11 N_XI0/XI17/XI11/NET36_XI0/XI17/XI11/MM11_d
+ N_XI0/XI17/XI11/NET35_XI0/XI17/XI11/MM11_g N_VDD_XI0/XI17/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI12/MM2 N_XI0/XI17/XI12/NET34_XI0/XI17/XI12/MM2_d
+ N_XI0/XI17/XI12/NET33_XI0/XI17/XI12/MM2_g N_VSS_XI0/XI17/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM3 N_XI0/XI17/XI12/NET33_XI0/XI17/XI12/MM3_d
+ N_WL<30>_XI0/XI17/XI12/MM3_g N_BLN<3>_XI0/XI17/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM0 N_XI0/XI17/XI12/NET34_XI0/XI17/XI12/MM0_d
+ N_WL<30>_XI0/XI17/XI12/MM0_g N_BL<3>_XI0/XI17/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM1 N_XI0/XI17/XI12/NET33_XI0/XI17/XI12/MM1_d
+ N_XI0/XI17/XI12/NET34_XI0/XI17/XI12/MM1_g N_VSS_XI0/XI17/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM9 N_XI0/XI17/XI12/NET36_XI0/XI17/XI12/MM9_d
+ N_WL<31>_XI0/XI17/XI12/MM9_g N_BL<3>_XI0/XI17/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM6 N_XI0/XI17/XI12/NET35_XI0/XI17/XI12/MM6_d
+ N_XI0/XI17/XI12/NET36_XI0/XI17/XI12/MM6_g N_VSS_XI0/XI17/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM7 N_XI0/XI17/XI12/NET36_XI0/XI17/XI12/MM7_d
+ N_XI0/XI17/XI12/NET35_XI0/XI17/XI12/MM7_g N_VSS_XI0/XI17/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM8 N_XI0/XI17/XI12/NET35_XI0/XI17/XI12/MM8_d
+ N_WL<31>_XI0/XI17/XI12/MM8_g N_BLN<3>_XI0/XI17/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI12/MM5 N_XI0/XI17/XI12/NET34_XI0/XI17/XI12/MM5_d
+ N_XI0/XI17/XI12/NET33_XI0/XI17/XI12/MM5_g N_VDD_XI0/XI17/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI12/MM4 N_XI0/XI17/XI12/NET33_XI0/XI17/XI12/MM4_d
+ N_XI0/XI17/XI12/NET34_XI0/XI17/XI12/MM4_g N_VDD_XI0/XI17/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI12/MM10 N_XI0/XI17/XI12/NET35_XI0/XI17/XI12/MM10_d
+ N_XI0/XI17/XI12/NET36_XI0/XI17/XI12/MM10_g N_VDD_XI0/XI17/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI12/MM11 N_XI0/XI17/XI12/NET36_XI0/XI17/XI12/MM11_d
+ N_XI0/XI17/XI12/NET35_XI0/XI17/XI12/MM11_g N_VDD_XI0/XI17/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI13/MM2 N_XI0/XI17/XI13/NET34_XI0/XI17/XI13/MM2_d
+ N_XI0/XI17/XI13/NET33_XI0/XI17/XI13/MM2_g N_VSS_XI0/XI17/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM3 N_XI0/XI17/XI13/NET33_XI0/XI17/XI13/MM3_d
+ N_WL<30>_XI0/XI17/XI13/MM3_g N_BLN<2>_XI0/XI17/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM0 N_XI0/XI17/XI13/NET34_XI0/XI17/XI13/MM0_d
+ N_WL<30>_XI0/XI17/XI13/MM0_g N_BL<2>_XI0/XI17/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM1 N_XI0/XI17/XI13/NET33_XI0/XI17/XI13/MM1_d
+ N_XI0/XI17/XI13/NET34_XI0/XI17/XI13/MM1_g N_VSS_XI0/XI17/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM9 N_XI0/XI17/XI13/NET36_XI0/XI17/XI13/MM9_d
+ N_WL<31>_XI0/XI17/XI13/MM9_g N_BL<2>_XI0/XI17/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM6 N_XI0/XI17/XI13/NET35_XI0/XI17/XI13/MM6_d
+ N_XI0/XI17/XI13/NET36_XI0/XI17/XI13/MM6_g N_VSS_XI0/XI17/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM7 N_XI0/XI17/XI13/NET36_XI0/XI17/XI13/MM7_d
+ N_XI0/XI17/XI13/NET35_XI0/XI17/XI13/MM7_g N_VSS_XI0/XI17/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM8 N_XI0/XI17/XI13/NET35_XI0/XI17/XI13/MM8_d
+ N_WL<31>_XI0/XI17/XI13/MM8_g N_BLN<2>_XI0/XI17/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI13/MM5 N_XI0/XI17/XI13/NET34_XI0/XI17/XI13/MM5_d
+ N_XI0/XI17/XI13/NET33_XI0/XI17/XI13/MM5_g N_VDD_XI0/XI17/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI13/MM4 N_XI0/XI17/XI13/NET33_XI0/XI17/XI13/MM4_d
+ N_XI0/XI17/XI13/NET34_XI0/XI17/XI13/MM4_g N_VDD_XI0/XI17/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI13/MM10 N_XI0/XI17/XI13/NET35_XI0/XI17/XI13/MM10_d
+ N_XI0/XI17/XI13/NET36_XI0/XI17/XI13/MM10_g N_VDD_XI0/XI17/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI13/MM11 N_XI0/XI17/XI13/NET36_XI0/XI17/XI13/MM11_d
+ N_XI0/XI17/XI13/NET35_XI0/XI17/XI13/MM11_g N_VDD_XI0/XI17/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI14/MM2 N_XI0/XI17/XI14/NET34_XI0/XI17/XI14/MM2_d
+ N_XI0/XI17/XI14/NET33_XI0/XI17/XI14/MM2_g N_VSS_XI0/XI17/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM3 N_XI0/XI17/XI14/NET33_XI0/XI17/XI14/MM3_d
+ N_WL<30>_XI0/XI17/XI14/MM3_g N_BLN<1>_XI0/XI17/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM0 N_XI0/XI17/XI14/NET34_XI0/XI17/XI14/MM0_d
+ N_WL<30>_XI0/XI17/XI14/MM0_g N_BL<1>_XI0/XI17/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM1 N_XI0/XI17/XI14/NET33_XI0/XI17/XI14/MM1_d
+ N_XI0/XI17/XI14/NET34_XI0/XI17/XI14/MM1_g N_VSS_XI0/XI17/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM9 N_XI0/XI17/XI14/NET36_XI0/XI17/XI14/MM9_d
+ N_WL<31>_XI0/XI17/XI14/MM9_g N_BL<1>_XI0/XI17/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM6 N_XI0/XI17/XI14/NET35_XI0/XI17/XI14/MM6_d
+ N_XI0/XI17/XI14/NET36_XI0/XI17/XI14/MM6_g N_VSS_XI0/XI17/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM7 N_XI0/XI17/XI14/NET36_XI0/XI17/XI14/MM7_d
+ N_XI0/XI17/XI14/NET35_XI0/XI17/XI14/MM7_g N_VSS_XI0/XI17/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM8 N_XI0/XI17/XI14/NET35_XI0/XI17/XI14/MM8_d
+ N_WL<31>_XI0/XI17/XI14/MM8_g N_BLN<1>_XI0/XI17/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI14/MM5 N_XI0/XI17/XI14/NET34_XI0/XI17/XI14/MM5_d
+ N_XI0/XI17/XI14/NET33_XI0/XI17/XI14/MM5_g N_VDD_XI0/XI17/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI14/MM4 N_XI0/XI17/XI14/NET33_XI0/XI17/XI14/MM4_d
+ N_XI0/XI17/XI14/NET34_XI0/XI17/XI14/MM4_g N_VDD_XI0/XI17/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI14/MM10 N_XI0/XI17/XI14/NET35_XI0/XI17/XI14/MM10_d
+ N_XI0/XI17/XI14/NET36_XI0/XI17/XI14/MM10_g N_VDD_XI0/XI17/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI14/MM11 N_XI0/XI17/XI14/NET36_XI0/XI17/XI14/MM11_d
+ N_XI0/XI17/XI14/NET35_XI0/XI17/XI14/MM11_g N_VDD_XI0/XI17/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI15/MM2 N_XI0/XI17/XI15/NET34_XI0/XI17/XI15/MM2_d
+ N_XI0/XI17/XI15/NET33_XI0/XI17/XI15/MM2_g N_VSS_XI0/XI17/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM3 N_XI0/XI17/XI15/NET33_XI0/XI17/XI15/MM3_d
+ N_WL<30>_XI0/XI17/XI15/MM3_g N_BLN<0>_XI0/XI17/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM0 N_XI0/XI17/XI15/NET34_XI0/XI17/XI15/MM0_d
+ N_WL<30>_XI0/XI17/XI15/MM0_g N_BL<0>_XI0/XI17/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM1 N_XI0/XI17/XI15/NET33_XI0/XI17/XI15/MM1_d
+ N_XI0/XI17/XI15/NET34_XI0/XI17/XI15/MM1_g N_VSS_XI0/XI17/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM9 N_XI0/XI17/XI15/NET36_XI0/XI17/XI15/MM9_d
+ N_WL<31>_XI0/XI17/XI15/MM9_g N_BL<0>_XI0/XI17/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM6 N_XI0/XI17/XI15/NET35_XI0/XI17/XI15/MM6_d
+ N_XI0/XI17/XI15/NET36_XI0/XI17/XI15/MM6_g N_VSS_XI0/XI17/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM7 N_XI0/XI17/XI15/NET36_XI0/XI17/XI15/MM7_d
+ N_XI0/XI17/XI15/NET35_XI0/XI17/XI15/MM7_g N_VSS_XI0/XI17/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM8 N_XI0/XI17/XI15/NET35_XI0/XI17/XI15/MM8_d
+ N_WL<31>_XI0/XI17/XI15/MM8_g N_BLN<0>_XI0/XI17/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI17/XI15/MM5 N_XI0/XI17/XI15/NET34_XI0/XI17/XI15/MM5_d
+ N_XI0/XI17/XI15/NET33_XI0/XI17/XI15/MM5_g N_VDD_XI0/XI17/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI15/MM4 N_XI0/XI17/XI15/NET33_XI0/XI17/XI15/MM4_d
+ N_XI0/XI17/XI15/NET34_XI0/XI17/XI15/MM4_g N_VDD_XI0/XI17/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI15/MM10 N_XI0/XI17/XI15/NET35_XI0/XI17/XI15/MM10_d
+ N_XI0/XI17/XI15/NET36_XI0/XI17/XI15/MM10_g N_VDD_XI0/XI17/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI17/XI15/MM11 N_XI0/XI17/XI15/NET36_XI0/XI17/XI15/MM11_d
+ N_XI0/XI17/XI15/NET35_XI0/XI17/XI15/MM11_g N_VDD_XI0/XI17/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI0/MM2 N_XI0/XI18/XI0/NET34_XI0/XI18/XI0/MM2_d
+ N_XI0/XI18/XI0/NET33_XI0/XI18/XI0/MM2_g N_VSS_XI0/XI18/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM3 N_XI0/XI18/XI0/NET33_XI0/XI18/XI0/MM3_d
+ N_WL<32>_XI0/XI18/XI0/MM3_g N_BLN<15>_XI0/XI18/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM0 N_XI0/XI18/XI0/NET34_XI0/XI18/XI0/MM0_d
+ N_WL<32>_XI0/XI18/XI0/MM0_g N_BL<15>_XI0/XI18/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM1 N_XI0/XI18/XI0/NET33_XI0/XI18/XI0/MM1_d
+ N_XI0/XI18/XI0/NET34_XI0/XI18/XI0/MM1_g N_VSS_XI0/XI18/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM9 N_XI0/XI18/XI0/NET36_XI0/XI18/XI0/MM9_d
+ N_WL<33>_XI0/XI18/XI0/MM9_g N_BL<15>_XI0/XI18/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM6 N_XI0/XI18/XI0/NET35_XI0/XI18/XI0/MM6_d
+ N_XI0/XI18/XI0/NET36_XI0/XI18/XI0/MM6_g N_VSS_XI0/XI18/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM7 N_XI0/XI18/XI0/NET36_XI0/XI18/XI0/MM7_d
+ N_XI0/XI18/XI0/NET35_XI0/XI18/XI0/MM7_g N_VSS_XI0/XI18/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM8 N_XI0/XI18/XI0/NET35_XI0/XI18/XI0/MM8_d
+ N_WL<33>_XI0/XI18/XI0/MM8_g N_BLN<15>_XI0/XI18/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI0/MM5 N_XI0/XI18/XI0/NET34_XI0/XI18/XI0/MM5_d
+ N_XI0/XI18/XI0/NET33_XI0/XI18/XI0/MM5_g N_VDD_XI0/XI18/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI0/MM4 N_XI0/XI18/XI0/NET33_XI0/XI18/XI0/MM4_d
+ N_XI0/XI18/XI0/NET34_XI0/XI18/XI0/MM4_g N_VDD_XI0/XI18/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI0/MM10 N_XI0/XI18/XI0/NET35_XI0/XI18/XI0/MM10_d
+ N_XI0/XI18/XI0/NET36_XI0/XI18/XI0/MM10_g N_VDD_XI0/XI18/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI0/MM11 N_XI0/XI18/XI0/NET36_XI0/XI18/XI0/MM11_d
+ N_XI0/XI18/XI0/NET35_XI0/XI18/XI0/MM11_g N_VDD_XI0/XI18/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI1/MM2 N_XI0/XI18/XI1/NET34_XI0/XI18/XI1/MM2_d
+ N_XI0/XI18/XI1/NET33_XI0/XI18/XI1/MM2_g N_VSS_XI0/XI18/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM3 N_XI0/XI18/XI1/NET33_XI0/XI18/XI1/MM3_d
+ N_WL<32>_XI0/XI18/XI1/MM3_g N_BLN<14>_XI0/XI18/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM0 N_XI0/XI18/XI1/NET34_XI0/XI18/XI1/MM0_d
+ N_WL<32>_XI0/XI18/XI1/MM0_g N_BL<14>_XI0/XI18/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM1 N_XI0/XI18/XI1/NET33_XI0/XI18/XI1/MM1_d
+ N_XI0/XI18/XI1/NET34_XI0/XI18/XI1/MM1_g N_VSS_XI0/XI18/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM9 N_XI0/XI18/XI1/NET36_XI0/XI18/XI1/MM9_d
+ N_WL<33>_XI0/XI18/XI1/MM9_g N_BL<14>_XI0/XI18/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM6 N_XI0/XI18/XI1/NET35_XI0/XI18/XI1/MM6_d
+ N_XI0/XI18/XI1/NET36_XI0/XI18/XI1/MM6_g N_VSS_XI0/XI18/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM7 N_XI0/XI18/XI1/NET36_XI0/XI18/XI1/MM7_d
+ N_XI0/XI18/XI1/NET35_XI0/XI18/XI1/MM7_g N_VSS_XI0/XI18/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM8 N_XI0/XI18/XI1/NET35_XI0/XI18/XI1/MM8_d
+ N_WL<33>_XI0/XI18/XI1/MM8_g N_BLN<14>_XI0/XI18/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI1/MM5 N_XI0/XI18/XI1/NET34_XI0/XI18/XI1/MM5_d
+ N_XI0/XI18/XI1/NET33_XI0/XI18/XI1/MM5_g N_VDD_XI0/XI18/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI1/MM4 N_XI0/XI18/XI1/NET33_XI0/XI18/XI1/MM4_d
+ N_XI0/XI18/XI1/NET34_XI0/XI18/XI1/MM4_g N_VDD_XI0/XI18/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI1/MM10 N_XI0/XI18/XI1/NET35_XI0/XI18/XI1/MM10_d
+ N_XI0/XI18/XI1/NET36_XI0/XI18/XI1/MM10_g N_VDD_XI0/XI18/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI1/MM11 N_XI0/XI18/XI1/NET36_XI0/XI18/XI1/MM11_d
+ N_XI0/XI18/XI1/NET35_XI0/XI18/XI1/MM11_g N_VDD_XI0/XI18/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI2/MM2 N_XI0/XI18/XI2/NET34_XI0/XI18/XI2/MM2_d
+ N_XI0/XI18/XI2/NET33_XI0/XI18/XI2/MM2_g N_VSS_XI0/XI18/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM3 N_XI0/XI18/XI2/NET33_XI0/XI18/XI2/MM3_d
+ N_WL<32>_XI0/XI18/XI2/MM3_g N_BLN<13>_XI0/XI18/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM0 N_XI0/XI18/XI2/NET34_XI0/XI18/XI2/MM0_d
+ N_WL<32>_XI0/XI18/XI2/MM0_g N_BL<13>_XI0/XI18/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM1 N_XI0/XI18/XI2/NET33_XI0/XI18/XI2/MM1_d
+ N_XI0/XI18/XI2/NET34_XI0/XI18/XI2/MM1_g N_VSS_XI0/XI18/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM9 N_XI0/XI18/XI2/NET36_XI0/XI18/XI2/MM9_d
+ N_WL<33>_XI0/XI18/XI2/MM9_g N_BL<13>_XI0/XI18/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM6 N_XI0/XI18/XI2/NET35_XI0/XI18/XI2/MM6_d
+ N_XI0/XI18/XI2/NET36_XI0/XI18/XI2/MM6_g N_VSS_XI0/XI18/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM7 N_XI0/XI18/XI2/NET36_XI0/XI18/XI2/MM7_d
+ N_XI0/XI18/XI2/NET35_XI0/XI18/XI2/MM7_g N_VSS_XI0/XI18/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM8 N_XI0/XI18/XI2/NET35_XI0/XI18/XI2/MM8_d
+ N_WL<33>_XI0/XI18/XI2/MM8_g N_BLN<13>_XI0/XI18/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI2/MM5 N_XI0/XI18/XI2/NET34_XI0/XI18/XI2/MM5_d
+ N_XI0/XI18/XI2/NET33_XI0/XI18/XI2/MM5_g N_VDD_XI0/XI18/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI2/MM4 N_XI0/XI18/XI2/NET33_XI0/XI18/XI2/MM4_d
+ N_XI0/XI18/XI2/NET34_XI0/XI18/XI2/MM4_g N_VDD_XI0/XI18/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI2/MM10 N_XI0/XI18/XI2/NET35_XI0/XI18/XI2/MM10_d
+ N_XI0/XI18/XI2/NET36_XI0/XI18/XI2/MM10_g N_VDD_XI0/XI18/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI2/MM11 N_XI0/XI18/XI2/NET36_XI0/XI18/XI2/MM11_d
+ N_XI0/XI18/XI2/NET35_XI0/XI18/XI2/MM11_g N_VDD_XI0/XI18/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI3/MM2 N_XI0/XI18/XI3/NET34_XI0/XI18/XI3/MM2_d
+ N_XI0/XI18/XI3/NET33_XI0/XI18/XI3/MM2_g N_VSS_XI0/XI18/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM3 N_XI0/XI18/XI3/NET33_XI0/XI18/XI3/MM3_d
+ N_WL<32>_XI0/XI18/XI3/MM3_g N_BLN<12>_XI0/XI18/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM0 N_XI0/XI18/XI3/NET34_XI0/XI18/XI3/MM0_d
+ N_WL<32>_XI0/XI18/XI3/MM0_g N_BL<12>_XI0/XI18/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM1 N_XI0/XI18/XI3/NET33_XI0/XI18/XI3/MM1_d
+ N_XI0/XI18/XI3/NET34_XI0/XI18/XI3/MM1_g N_VSS_XI0/XI18/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM9 N_XI0/XI18/XI3/NET36_XI0/XI18/XI3/MM9_d
+ N_WL<33>_XI0/XI18/XI3/MM9_g N_BL<12>_XI0/XI18/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM6 N_XI0/XI18/XI3/NET35_XI0/XI18/XI3/MM6_d
+ N_XI0/XI18/XI3/NET36_XI0/XI18/XI3/MM6_g N_VSS_XI0/XI18/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM7 N_XI0/XI18/XI3/NET36_XI0/XI18/XI3/MM7_d
+ N_XI0/XI18/XI3/NET35_XI0/XI18/XI3/MM7_g N_VSS_XI0/XI18/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM8 N_XI0/XI18/XI3/NET35_XI0/XI18/XI3/MM8_d
+ N_WL<33>_XI0/XI18/XI3/MM8_g N_BLN<12>_XI0/XI18/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI3/MM5 N_XI0/XI18/XI3/NET34_XI0/XI18/XI3/MM5_d
+ N_XI0/XI18/XI3/NET33_XI0/XI18/XI3/MM5_g N_VDD_XI0/XI18/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI3/MM4 N_XI0/XI18/XI3/NET33_XI0/XI18/XI3/MM4_d
+ N_XI0/XI18/XI3/NET34_XI0/XI18/XI3/MM4_g N_VDD_XI0/XI18/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI3/MM10 N_XI0/XI18/XI3/NET35_XI0/XI18/XI3/MM10_d
+ N_XI0/XI18/XI3/NET36_XI0/XI18/XI3/MM10_g N_VDD_XI0/XI18/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI3/MM11 N_XI0/XI18/XI3/NET36_XI0/XI18/XI3/MM11_d
+ N_XI0/XI18/XI3/NET35_XI0/XI18/XI3/MM11_g N_VDD_XI0/XI18/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI4/MM2 N_XI0/XI18/XI4/NET34_XI0/XI18/XI4/MM2_d
+ N_XI0/XI18/XI4/NET33_XI0/XI18/XI4/MM2_g N_VSS_XI0/XI18/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM3 N_XI0/XI18/XI4/NET33_XI0/XI18/XI4/MM3_d
+ N_WL<32>_XI0/XI18/XI4/MM3_g N_BLN<11>_XI0/XI18/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM0 N_XI0/XI18/XI4/NET34_XI0/XI18/XI4/MM0_d
+ N_WL<32>_XI0/XI18/XI4/MM0_g N_BL<11>_XI0/XI18/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM1 N_XI0/XI18/XI4/NET33_XI0/XI18/XI4/MM1_d
+ N_XI0/XI18/XI4/NET34_XI0/XI18/XI4/MM1_g N_VSS_XI0/XI18/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM9 N_XI0/XI18/XI4/NET36_XI0/XI18/XI4/MM9_d
+ N_WL<33>_XI0/XI18/XI4/MM9_g N_BL<11>_XI0/XI18/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM6 N_XI0/XI18/XI4/NET35_XI0/XI18/XI4/MM6_d
+ N_XI0/XI18/XI4/NET36_XI0/XI18/XI4/MM6_g N_VSS_XI0/XI18/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM7 N_XI0/XI18/XI4/NET36_XI0/XI18/XI4/MM7_d
+ N_XI0/XI18/XI4/NET35_XI0/XI18/XI4/MM7_g N_VSS_XI0/XI18/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM8 N_XI0/XI18/XI4/NET35_XI0/XI18/XI4/MM8_d
+ N_WL<33>_XI0/XI18/XI4/MM8_g N_BLN<11>_XI0/XI18/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI4/MM5 N_XI0/XI18/XI4/NET34_XI0/XI18/XI4/MM5_d
+ N_XI0/XI18/XI4/NET33_XI0/XI18/XI4/MM5_g N_VDD_XI0/XI18/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI4/MM4 N_XI0/XI18/XI4/NET33_XI0/XI18/XI4/MM4_d
+ N_XI0/XI18/XI4/NET34_XI0/XI18/XI4/MM4_g N_VDD_XI0/XI18/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI4/MM10 N_XI0/XI18/XI4/NET35_XI0/XI18/XI4/MM10_d
+ N_XI0/XI18/XI4/NET36_XI0/XI18/XI4/MM10_g N_VDD_XI0/XI18/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI4/MM11 N_XI0/XI18/XI4/NET36_XI0/XI18/XI4/MM11_d
+ N_XI0/XI18/XI4/NET35_XI0/XI18/XI4/MM11_g N_VDD_XI0/XI18/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI5/MM2 N_XI0/XI18/XI5/NET34_XI0/XI18/XI5/MM2_d
+ N_XI0/XI18/XI5/NET33_XI0/XI18/XI5/MM2_g N_VSS_XI0/XI18/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM3 N_XI0/XI18/XI5/NET33_XI0/XI18/XI5/MM3_d
+ N_WL<32>_XI0/XI18/XI5/MM3_g N_BLN<10>_XI0/XI18/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM0 N_XI0/XI18/XI5/NET34_XI0/XI18/XI5/MM0_d
+ N_WL<32>_XI0/XI18/XI5/MM0_g N_BL<10>_XI0/XI18/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM1 N_XI0/XI18/XI5/NET33_XI0/XI18/XI5/MM1_d
+ N_XI0/XI18/XI5/NET34_XI0/XI18/XI5/MM1_g N_VSS_XI0/XI18/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM9 N_XI0/XI18/XI5/NET36_XI0/XI18/XI5/MM9_d
+ N_WL<33>_XI0/XI18/XI5/MM9_g N_BL<10>_XI0/XI18/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM6 N_XI0/XI18/XI5/NET35_XI0/XI18/XI5/MM6_d
+ N_XI0/XI18/XI5/NET36_XI0/XI18/XI5/MM6_g N_VSS_XI0/XI18/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM7 N_XI0/XI18/XI5/NET36_XI0/XI18/XI5/MM7_d
+ N_XI0/XI18/XI5/NET35_XI0/XI18/XI5/MM7_g N_VSS_XI0/XI18/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM8 N_XI0/XI18/XI5/NET35_XI0/XI18/XI5/MM8_d
+ N_WL<33>_XI0/XI18/XI5/MM8_g N_BLN<10>_XI0/XI18/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI5/MM5 N_XI0/XI18/XI5/NET34_XI0/XI18/XI5/MM5_d
+ N_XI0/XI18/XI5/NET33_XI0/XI18/XI5/MM5_g N_VDD_XI0/XI18/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI5/MM4 N_XI0/XI18/XI5/NET33_XI0/XI18/XI5/MM4_d
+ N_XI0/XI18/XI5/NET34_XI0/XI18/XI5/MM4_g N_VDD_XI0/XI18/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI5/MM10 N_XI0/XI18/XI5/NET35_XI0/XI18/XI5/MM10_d
+ N_XI0/XI18/XI5/NET36_XI0/XI18/XI5/MM10_g N_VDD_XI0/XI18/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI5/MM11 N_XI0/XI18/XI5/NET36_XI0/XI18/XI5/MM11_d
+ N_XI0/XI18/XI5/NET35_XI0/XI18/XI5/MM11_g N_VDD_XI0/XI18/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI6/MM2 N_XI0/XI18/XI6/NET34_XI0/XI18/XI6/MM2_d
+ N_XI0/XI18/XI6/NET33_XI0/XI18/XI6/MM2_g N_VSS_XI0/XI18/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM3 N_XI0/XI18/XI6/NET33_XI0/XI18/XI6/MM3_d
+ N_WL<32>_XI0/XI18/XI6/MM3_g N_BLN<9>_XI0/XI18/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM0 N_XI0/XI18/XI6/NET34_XI0/XI18/XI6/MM0_d
+ N_WL<32>_XI0/XI18/XI6/MM0_g N_BL<9>_XI0/XI18/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM1 N_XI0/XI18/XI6/NET33_XI0/XI18/XI6/MM1_d
+ N_XI0/XI18/XI6/NET34_XI0/XI18/XI6/MM1_g N_VSS_XI0/XI18/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM9 N_XI0/XI18/XI6/NET36_XI0/XI18/XI6/MM9_d
+ N_WL<33>_XI0/XI18/XI6/MM9_g N_BL<9>_XI0/XI18/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM6 N_XI0/XI18/XI6/NET35_XI0/XI18/XI6/MM6_d
+ N_XI0/XI18/XI6/NET36_XI0/XI18/XI6/MM6_g N_VSS_XI0/XI18/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM7 N_XI0/XI18/XI6/NET36_XI0/XI18/XI6/MM7_d
+ N_XI0/XI18/XI6/NET35_XI0/XI18/XI6/MM7_g N_VSS_XI0/XI18/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM8 N_XI0/XI18/XI6/NET35_XI0/XI18/XI6/MM8_d
+ N_WL<33>_XI0/XI18/XI6/MM8_g N_BLN<9>_XI0/XI18/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI6/MM5 N_XI0/XI18/XI6/NET34_XI0/XI18/XI6/MM5_d
+ N_XI0/XI18/XI6/NET33_XI0/XI18/XI6/MM5_g N_VDD_XI0/XI18/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI6/MM4 N_XI0/XI18/XI6/NET33_XI0/XI18/XI6/MM4_d
+ N_XI0/XI18/XI6/NET34_XI0/XI18/XI6/MM4_g N_VDD_XI0/XI18/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI6/MM10 N_XI0/XI18/XI6/NET35_XI0/XI18/XI6/MM10_d
+ N_XI0/XI18/XI6/NET36_XI0/XI18/XI6/MM10_g N_VDD_XI0/XI18/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI6/MM11 N_XI0/XI18/XI6/NET36_XI0/XI18/XI6/MM11_d
+ N_XI0/XI18/XI6/NET35_XI0/XI18/XI6/MM11_g N_VDD_XI0/XI18/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI7/MM2 N_XI0/XI18/XI7/NET34_XI0/XI18/XI7/MM2_d
+ N_XI0/XI18/XI7/NET33_XI0/XI18/XI7/MM2_g N_VSS_XI0/XI18/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM3 N_XI0/XI18/XI7/NET33_XI0/XI18/XI7/MM3_d
+ N_WL<32>_XI0/XI18/XI7/MM3_g N_BLN<8>_XI0/XI18/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM0 N_XI0/XI18/XI7/NET34_XI0/XI18/XI7/MM0_d
+ N_WL<32>_XI0/XI18/XI7/MM0_g N_BL<8>_XI0/XI18/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM1 N_XI0/XI18/XI7/NET33_XI0/XI18/XI7/MM1_d
+ N_XI0/XI18/XI7/NET34_XI0/XI18/XI7/MM1_g N_VSS_XI0/XI18/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM9 N_XI0/XI18/XI7/NET36_XI0/XI18/XI7/MM9_d
+ N_WL<33>_XI0/XI18/XI7/MM9_g N_BL<8>_XI0/XI18/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM6 N_XI0/XI18/XI7/NET35_XI0/XI18/XI7/MM6_d
+ N_XI0/XI18/XI7/NET36_XI0/XI18/XI7/MM6_g N_VSS_XI0/XI18/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM7 N_XI0/XI18/XI7/NET36_XI0/XI18/XI7/MM7_d
+ N_XI0/XI18/XI7/NET35_XI0/XI18/XI7/MM7_g N_VSS_XI0/XI18/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM8 N_XI0/XI18/XI7/NET35_XI0/XI18/XI7/MM8_d
+ N_WL<33>_XI0/XI18/XI7/MM8_g N_BLN<8>_XI0/XI18/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI7/MM5 N_XI0/XI18/XI7/NET34_XI0/XI18/XI7/MM5_d
+ N_XI0/XI18/XI7/NET33_XI0/XI18/XI7/MM5_g N_VDD_XI0/XI18/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI7/MM4 N_XI0/XI18/XI7/NET33_XI0/XI18/XI7/MM4_d
+ N_XI0/XI18/XI7/NET34_XI0/XI18/XI7/MM4_g N_VDD_XI0/XI18/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI7/MM10 N_XI0/XI18/XI7/NET35_XI0/XI18/XI7/MM10_d
+ N_XI0/XI18/XI7/NET36_XI0/XI18/XI7/MM10_g N_VDD_XI0/XI18/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI7/MM11 N_XI0/XI18/XI7/NET36_XI0/XI18/XI7/MM11_d
+ N_XI0/XI18/XI7/NET35_XI0/XI18/XI7/MM11_g N_VDD_XI0/XI18/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI8/MM2 N_XI0/XI18/XI8/NET34_XI0/XI18/XI8/MM2_d
+ N_XI0/XI18/XI8/NET33_XI0/XI18/XI8/MM2_g N_VSS_XI0/XI18/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM3 N_XI0/XI18/XI8/NET33_XI0/XI18/XI8/MM3_d
+ N_WL<32>_XI0/XI18/XI8/MM3_g N_BLN<7>_XI0/XI18/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM0 N_XI0/XI18/XI8/NET34_XI0/XI18/XI8/MM0_d
+ N_WL<32>_XI0/XI18/XI8/MM0_g N_BL<7>_XI0/XI18/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM1 N_XI0/XI18/XI8/NET33_XI0/XI18/XI8/MM1_d
+ N_XI0/XI18/XI8/NET34_XI0/XI18/XI8/MM1_g N_VSS_XI0/XI18/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM9 N_XI0/XI18/XI8/NET36_XI0/XI18/XI8/MM9_d
+ N_WL<33>_XI0/XI18/XI8/MM9_g N_BL<7>_XI0/XI18/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM6 N_XI0/XI18/XI8/NET35_XI0/XI18/XI8/MM6_d
+ N_XI0/XI18/XI8/NET36_XI0/XI18/XI8/MM6_g N_VSS_XI0/XI18/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM7 N_XI0/XI18/XI8/NET36_XI0/XI18/XI8/MM7_d
+ N_XI0/XI18/XI8/NET35_XI0/XI18/XI8/MM7_g N_VSS_XI0/XI18/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM8 N_XI0/XI18/XI8/NET35_XI0/XI18/XI8/MM8_d
+ N_WL<33>_XI0/XI18/XI8/MM8_g N_BLN<7>_XI0/XI18/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI8/MM5 N_XI0/XI18/XI8/NET34_XI0/XI18/XI8/MM5_d
+ N_XI0/XI18/XI8/NET33_XI0/XI18/XI8/MM5_g N_VDD_XI0/XI18/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI8/MM4 N_XI0/XI18/XI8/NET33_XI0/XI18/XI8/MM4_d
+ N_XI0/XI18/XI8/NET34_XI0/XI18/XI8/MM4_g N_VDD_XI0/XI18/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI8/MM10 N_XI0/XI18/XI8/NET35_XI0/XI18/XI8/MM10_d
+ N_XI0/XI18/XI8/NET36_XI0/XI18/XI8/MM10_g N_VDD_XI0/XI18/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI8/MM11 N_XI0/XI18/XI8/NET36_XI0/XI18/XI8/MM11_d
+ N_XI0/XI18/XI8/NET35_XI0/XI18/XI8/MM11_g N_VDD_XI0/XI18/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI9/MM2 N_XI0/XI18/XI9/NET34_XI0/XI18/XI9/MM2_d
+ N_XI0/XI18/XI9/NET33_XI0/XI18/XI9/MM2_g N_VSS_XI0/XI18/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM3 N_XI0/XI18/XI9/NET33_XI0/XI18/XI9/MM3_d
+ N_WL<32>_XI0/XI18/XI9/MM3_g N_BLN<6>_XI0/XI18/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM0 N_XI0/XI18/XI9/NET34_XI0/XI18/XI9/MM0_d
+ N_WL<32>_XI0/XI18/XI9/MM0_g N_BL<6>_XI0/XI18/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM1 N_XI0/XI18/XI9/NET33_XI0/XI18/XI9/MM1_d
+ N_XI0/XI18/XI9/NET34_XI0/XI18/XI9/MM1_g N_VSS_XI0/XI18/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM9 N_XI0/XI18/XI9/NET36_XI0/XI18/XI9/MM9_d
+ N_WL<33>_XI0/XI18/XI9/MM9_g N_BL<6>_XI0/XI18/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM6 N_XI0/XI18/XI9/NET35_XI0/XI18/XI9/MM6_d
+ N_XI0/XI18/XI9/NET36_XI0/XI18/XI9/MM6_g N_VSS_XI0/XI18/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM7 N_XI0/XI18/XI9/NET36_XI0/XI18/XI9/MM7_d
+ N_XI0/XI18/XI9/NET35_XI0/XI18/XI9/MM7_g N_VSS_XI0/XI18/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM8 N_XI0/XI18/XI9/NET35_XI0/XI18/XI9/MM8_d
+ N_WL<33>_XI0/XI18/XI9/MM8_g N_BLN<6>_XI0/XI18/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI9/MM5 N_XI0/XI18/XI9/NET34_XI0/XI18/XI9/MM5_d
+ N_XI0/XI18/XI9/NET33_XI0/XI18/XI9/MM5_g N_VDD_XI0/XI18/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI9/MM4 N_XI0/XI18/XI9/NET33_XI0/XI18/XI9/MM4_d
+ N_XI0/XI18/XI9/NET34_XI0/XI18/XI9/MM4_g N_VDD_XI0/XI18/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI9/MM10 N_XI0/XI18/XI9/NET35_XI0/XI18/XI9/MM10_d
+ N_XI0/XI18/XI9/NET36_XI0/XI18/XI9/MM10_g N_VDD_XI0/XI18/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI9/MM11 N_XI0/XI18/XI9/NET36_XI0/XI18/XI9/MM11_d
+ N_XI0/XI18/XI9/NET35_XI0/XI18/XI9/MM11_g N_VDD_XI0/XI18/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI10/MM2 N_XI0/XI18/XI10/NET34_XI0/XI18/XI10/MM2_d
+ N_XI0/XI18/XI10/NET33_XI0/XI18/XI10/MM2_g N_VSS_XI0/XI18/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM3 N_XI0/XI18/XI10/NET33_XI0/XI18/XI10/MM3_d
+ N_WL<32>_XI0/XI18/XI10/MM3_g N_BLN<5>_XI0/XI18/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM0 N_XI0/XI18/XI10/NET34_XI0/XI18/XI10/MM0_d
+ N_WL<32>_XI0/XI18/XI10/MM0_g N_BL<5>_XI0/XI18/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM1 N_XI0/XI18/XI10/NET33_XI0/XI18/XI10/MM1_d
+ N_XI0/XI18/XI10/NET34_XI0/XI18/XI10/MM1_g N_VSS_XI0/XI18/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM9 N_XI0/XI18/XI10/NET36_XI0/XI18/XI10/MM9_d
+ N_WL<33>_XI0/XI18/XI10/MM9_g N_BL<5>_XI0/XI18/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM6 N_XI0/XI18/XI10/NET35_XI0/XI18/XI10/MM6_d
+ N_XI0/XI18/XI10/NET36_XI0/XI18/XI10/MM6_g N_VSS_XI0/XI18/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM7 N_XI0/XI18/XI10/NET36_XI0/XI18/XI10/MM7_d
+ N_XI0/XI18/XI10/NET35_XI0/XI18/XI10/MM7_g N_VSS_XI0/XI18/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM8 N_XI0/XI18/XI10/NET35_XI0/XI18/XI10/MM8_d
+ N_WL<33>_XI0/XI18/XI10/MM8_g N_BLN<5>_XI0/XI18/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI10/MM5 N_XI0/XI18/XI10/NET34_XI0/XI18/XI10/MM5_d
+ N_XI0/XI18/XI10/NET33_XI0/XI18/XI10/MM5_g N_VDD_XI0/XI18/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI10/MM4 N_XI0/XI18/XI10/NET33_XI0/XI18/XI10/MM4_d
+ N_XI0/XI18/XI10/NET34_XI0/XI18/XI10/MM4_g N_VDD_XI0/XI18/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI10/MM10 N_XI0/XI18/XI10/NET35_XI0/XI18/XI10/MM10_d
+ N_XI0/XI18/XI10/NET36_XI0/XI18/XI10/MM10_g N_VDD_XI0/XI18/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI10/MM11 N_XI0/XI18/XI10/NET36_XI0/XI18/XI10/MM11_d
+ N_XI0/XI18/XI10/NET35_XI0/XI18/XI10/MM11_g N_VDD_XI0/XI18/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI11/MM2 N_XI0/XI18/XI11/NET34_XI0/XI18/XI11/MM2_d
+ N_XI0/XI18/XI11/NET33_XI0/XI18/XI11/MM2_g N_VSS_XI0/XI18/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM3 N_XI0/XI18/XI11/NET33_XI0/XI18/XI11/MM3_d
+ N_WL<32>_XI0/XI18/XI11/MM3_g N_BLN<4>_XI0/XI18/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM0 N_XI0/XI18/XI11/NET34_XI0/XI18/XI11/MM0_d
+ N_WL<32>_XI0/XI18/XI11/MM0_g N_BL<4>_XI0/XI18/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM1 N_XI0/XI18/XI11/NET33_XI0/XI18/XI11/MM1_d
+ N_XI0/XI18/XI11/NET34_XI0/XI18/XI11/MM1_g N_VSS_XI0/XI18/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM9 N_XI0/XI18/XI11/NET36_XI0/XI18/XI11/MM9_d
+ N_WL<33>_XI0/XI18/XI11/MM9_g N_BL<4>_XI0/XI18/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM6 N_XI0/XI18/XI11/NET35_XI0/XI18/XI11/MM6_d
+ N_XI0/XI18/XI11/NET36_XI0/XI18/XI11/MM6_g N_VSS_XI0/XI18/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM7 N_XI0/XI18/XI11/NET36_XI0/XI18/XI11/MM7_d
+ N_XI0/XI18/XI11/NET35_XI0/XI18/XI11/MM7_g N_VSS_XI0/XI18/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM8 N_XI0/XI18/XI11/NET35_XI0/XI18/XI11/MM8_d
+ N_WL<33>_XI0/XI18/XI11/MM8_g N_BLN<4>_XI0/XI18/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI11/MM5 N_XI0/XI18/XI11/NET34_XI0/XI18/XI11/MM5_d
+ N_XI0/XI18/XI11/NET33_XI0/XI18/XI11/MM5_g N_VDD_XI0/XI18/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI11/MM4 N_XI0/XI18/XI11/NET33_XI0/XI18/XI11/MM4_d
+ N_XI0/XI18/XI11/NET34_XI0/XI18/XI11/MM4_g N_VDD_XI0/XI18/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI11/MM10 N_XI0/XI18/XI11/NET35_XI0/XI18/XI11/MM10_d
+ N_XI0/XI18/XI11/NET36_XI0/XI18/XI11/MM10_g N_VDD_XI0/XI18/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI11/MM11 N_XI0/XI18/XI11/NET36_XI0/XI18/XI11/MM11_d
+ N_XI0/XI18/XI11/NET35_XI0/XI18/XI11/MM11_g N_VDD_XI0/XI18/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI12/MM2 N_XI0/XI18/XI12/NET34_XI0/XI18/XI12/MM2_d
+ N_XI0/XI18/XI12/NET33_XI0/XI18/XI12/MM2_g N_VSS_XI0/XI18/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM3 N_XI0/XI18/XI12/NET33_XI0/XI18/XI12/MM3_d
+ N_WL<32>_XI0/XI18/XI12/MM3_g N_BLN<3>_XI0/XI18/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM0 N_XI0/XI18/XI12/NET34_XI0/XI18/XI12/MM0_d
+ N_WL<32>_XI0/XI18/XI12/MM0_g N_BL<3>_XI0/XI18/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM1 N_XI0/XI18/XI12/NET33_XI0/XI18/XI12/MM1_d
+ N_XI0/XI18/XI12/NET34_XI0/XI18/XI12/MM1_g N_VSS_XI0/XI18/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM9 N_XI0/XI18/XI12/NET36_XI0/XI18/XI12/MM9_d
+ N_WL<33>_XI0/XI18/XI12/MM9_g N_BL<3>_XI0/XI18/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM6 N_XI0/XI18/XI12/NET35_XI0/XI18/XI12/MM6_d
+ N_XI0/XI18/XI12/NET36_XI0/XI18/XI12/MM6_g N_VSS_XI0/XI18/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM7 N_XI0/XI18/XI12/NET36_XI0/XI18/XI12/MM7_d
+ N_XI0/XI18/XI12/NET35_XI0/XI18/XI12/MM7_g N_VSS_XI0/XI18/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM8 N_XI0/XI18/XI12/NET35_XI0/XI18/XI12/MM8_d
+ N_WL<33>_XI0/XI18/XI12/MM8_g N_BLN<3>_XI0/XI18/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI12/MM5 N_XI0/XI18/XI12/NET34_XI0/XI18/XI12/MM5_d
+ N_XI0/XI18/XI12/NET33_XI0/XI18/XI12/MM5_g N_VDD_XI0/XI18/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI12/MM4 N_XI0/XI18/XI12/NET33_XI0/XI18/XI12/MM4_d
+ N_XI0/XI18/XI12/NET34_XI0/XI18/XI12/MM4_g N_VDD_XI0/XI18/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI12/MM10 N_XI0/XI18/XI12/NET35_XI0/XI18/XI12/MM10_d
+ N_XI0/XI18/XI12/NET36_XI0/XI18/XI12/MM10_g N_VDD_XI0/XI18/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI12/MM11 N_XI0/XI18/XI12/NET36_XI0/XI18/XI12/MM11_d
+ N_XI0/XI18/XI12/NET35_XI0/XI18/XI12/MM11_g N_VDD_XI0/XI18/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI13/MM2 N_XI0/XI18/XI13/NET34_XI0/XI18/XI13/MM2_d
+ N_XI0/XI18/XI13/NET33_XI0/XI18/XI13/MM2_g N_VSS_XI0/XI18/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM3 N_XI0/XI18/XI13/NET33_XI0/XI18/XI13/MM3_d
+ N_WL<32>_XI0/XI18/XI13/MM3_g N_BLN<2>_XI0/XI18/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM0 N_XI0/XI18/XI13/NET34_XI0/XI18/XI13/MM0_d
+ N_WL<32>_XI0/XI18/XI13/MM0_g N_BL<2>_XI0/XI18/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM1 N_XI0/XI18/XI13/NET33_XI0/XI18/XI13/MM1_d
+ N_XI0/XI18/XI13/NET34_XI0/XI18/XI13/MM1_g N_VSS_XI0/XI18/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM9 N_XI0/XI18/XI13/NET36_XI0/XI18/XI13/MM9_d
+ N_WL<33>_XI0/XI18/XI13/MM9_g N_BL<2>_XI0/XI18/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM6 N_XI0/XI18/XI13/NET35_XI0/XI18/XI13/MM6_d
+ N_XI0/XI18/XI13/NET36_XI0/XI18/XI13/MM6_g N_VSS_XI0/XI18/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM7 N_XI0/XI18/XI13/NET36_XI0/XI18/XI13/MM7_d
+ N_XI0/XI18/XI13/NET35_XI0/XI18/XI13/MM7_g N_VSS_XI0/XI18/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM8 N_XI0/XI18/XI13/NET35_XI0/XI18/XI13/MM8_d
+ N_WL<33>_XI0/XI18/XI13/MM8_g N_BLN<2>_XI0/XI18/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI13/MM5 N_XI0/XI18/XI13/NET34_XI0/XI18/XI13/MM5_d
+ N_XI0/XI18/XI13/NET33_XI0/XI18/XI13/MM5_g N_VDD_XI0/XI18/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI13/MM4 N_XI0/XI18/XI13/NET33_XI0/XI18/XI13/MM4_d
+ N_XI0/XI18/XI13/NET34_XI0/XI18/XI13/MM4_g N_VDD_XI0/XI18/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI13/MM10 N_XI0/XI18/XI13/NET35_XI0/XI18/XI13/MM10_d
+ N_XI0/XI18/XI13/NET36_XI0/XI18/XI13/MM10_g N_VDD_XI0/XI18/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI13/MM11 N_XI0/XI18/XI13/NET36_XI0/XI18/XI13/MM11_d
+ N_XI0/XI18/XI13/NET35_XI0/XI18/XI13/MM11_g N_VDD_XI0/XI18/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI14/MM2 N_XI0/XI18/XI14/NET34_XI0/XI18/XI14/MM2_d
+ N_XI0/XI18/XI14/NET33_XI0/XI18/XI14/MM2_g N_VSS_XI0/XI18/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM3 N_XI0/XI18/XI14/NET33_XI0/XI18/XI14/MM3_d
+ N_WL<32>_XI0/XI18/XI14/MM3_g N_BLN<1>_XI0/XI18/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM0 N_XI0/XI18/XI14/NET34_XI0/XI18/XI14/MM0_d
+ N_WL<32>_XI0/XI18/XI14/MM0_g N_BL<1>_XI0/XI18/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM1 N_XI0/XI18/XI14/NET33_XI0/XI18/XI14/MM1_d
+ N_XI0/XI18/XI14/NET34_XI0/XI18/XI14/MM1_g N_VSS_XI0/XI18/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM9 N_XI0/XI18/XI14/NET36_XI0/XI18/XI14/MM9_d
+ N_WL<33>_XI0/XI18/XI14/MM9_g N_BL<1>_XI0/XI18/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM6 N_XI0/XI18/XI14/NET35_XI0/XI18/XI14/MM6_d
+ N_XI0/XI18/XI14/NET36_XI0/XI18/XI14/MM6_g N_VSS_XI0/XI18/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM7 N_XI0/XI18/XI14/NET36_XI0/XI18/XI14/MM7_d
+ N_XI0/XI18/XI14/NET35_XI0/XI18/XI14/MM7_g N_VSS_XI0/XI18/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM8 N_XI0/XI18/XI14/NET35_XI0/XI18/XI14/MM8_d
+ N_WL<33>_XI0/XI18/XI14/MM8_g N_BLN<1>_XI0/XI18/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI14/MM5 N_XI0/XI18/XI14/NET34_XI0/XI18/XI14/MM5_d
+ N_XI0/XI18/XI14/NET33_XI0/XI18/XI14/MM5_g N_VDD_XI0/XI18/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI14/MM4 N_XI0/XI18/XI14/NET33_XI0/XI18/XI14/MM4_d
+ N_XI0/XI18/XI14/NET34_XI0/XI18/XI14/MM4_g N_VDD_XI0/XI18/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI14/MM10 N_XI0/XI18/XI14/NET35_XI0/XI18/XI14/MM10_d
+ N_XI0/XI18/XI14/NET36_XI0/XI18/XI14/MM10_g N_VDD_XI0/XI18/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI14/MM11 N_XI0/XI18/XI14/NET36_XI0/XI18/XI14/MM11_d
+ N_XI0/XI18/XI14/NET35_XI0/XI18/XI14/MM11_g N_VDD_XI0/XI18/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI15/MM2 N_XI0/XI18/XI15/NET34_XI0/XI18/XI15/MM2_d
+ N_XI0/XI18/XI15/NET33_XI0/XI18/XI15/MM2_g N_VSS_XI0/XI18/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM3 N_XI0/XI18/XI15/NET33_XI0/XI18/XI15/MM3_d
+ N_WL<32>_XI0/XI18/XI15/MM3_g N_BLN<0>_XI0/XI18/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM0 N_XI0/XI18/XI15/NET34_XI0/XI18/XI15/MM0_d
+ N_WL<32>_XI0/XI18/XI15/MM0_g N_BL<0>_XI0/XI18/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM1 N_XI0/XI18/XI15/NET33_XI0/XI18/XI15/MM1_d
+ N_XI0/XI18/XI15/NET34_XI0/XI18/XI15/MM1_g N_VSS_XI0/XI18/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM9 N_XI0/XI18/XI15/NET36_XI0/XI18/XI15/MM9_d
+ N_WL<33>_XI0/XI18/XI15/MM9_g N_BL<0>_XI0/XI18/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM6 N_XI0/XI18/XI15/NET35_XI0/XI18/XI15/MM6_d
+ N_XI0/XI18/XI15/NET36_XI0/XI18/XI15/MM6_g N_VSS_XI0/XI18/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM7 N_XI0/XI18/XI15/NET36_XI0/XI18/XI15/MM7_d
+ N_XI0/XI18/XI15/NET35_XI0/XI18/XI15/MM7_g N_VSS_XI0/XI18/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM8 N_XI0/XI18/XI15/NET35_XI0/XI18/XI15/MM8_d
+ N_WL<33>_XI0/XI18/XI15/MM8_g N_BLN<0>_XI0/XI18/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI18/XI15/MM5 N_XI0/XI18/XI15/NET34_XI0/XI18/XI15/MM5_d
+ N_XI0/XI18/XI15/NET33_XI0/XI18/XI15/MM5_g N_VDD_XI0/XI18/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI15/MM4 N_XI0/XI18/XI15/NET33_XI0/XI18/XI15/MM4_d
+ N_XI0/XI18/XI15/NET34_XI0/XI18/XI15/MM4_g N_VDD_XI0/XI18/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI15/MM10 N_XI0/XI18/XI15/NET35_XI0/XI18/XI15/MM10_d
+ N_XI0/XI18/XI15/NET36_XI0/XI18/XI15/MM10_g N_VDD_XI0/XI18/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI18/XI15/MM11 N_XI0/XI18/XI15/NET36_XI0/XI18/XI15/MM11_d
+ N_XI0/XI18/XI15/NET35_XI0/XI18/XI15/MM11_g N_VDD_XI0/XI18/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI0/MM2 N_XI0/XI19/XI0/NET34_XI0/XI19/XI0/MM2_d
+ N_XI0/XI19/XI0/NET33_XI0/XI19/XI0/MM2_g N_VSS_XI0/XI19/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM3 N_XI0/XI19/XI0/NET33_XI0/XI19/XI0/MM3_d
+ N_WL<34>_XI0/XI19/XI0/MM3_g N_BLN<15>_XI0/XI19/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM0 N_XI0/XI19/XI0/NET34_XI0/XI19/XI0/MM0_d
+ N_WL<34>_XI0/XI19/XI0/MM0_g N_BL<15>_XI0/XI19/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM1 N_XI0/XI19/XI0/NET33_XI0/XI19/XI0/MM1_d
+ N_XI0/XI19/XI0/NET34_XI0/XI19/XI0/MM1_g N_VSS_XI0/XI19/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM9 N_XI0/XI19/XI0/NET36_XI0/XI19/XI0/MM9_d
+ N_WL<35>_XI0/XI19/XI0/MM9_g N_BL<15>_XI0/XI19/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM6 N_XI0/XI19/XI0/NET35_XI0/XI19/XI0/MM6_d
+ N_XI0/XI19/XI0/NET36_XI0/XI19/XI0/MM6_g N_VSS_XI0/XI19/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM7 N_XI0/XI19/XI0/NET36_XI0/XI19/XI0/MM7_d
+ N_XI0/XI19/XI0/NET35_XI0/XI19/XI0/MM7_g N_VSS_XI0/XI19/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM8 N_XI0/XI19/XI0/NET35_XI0/XI19/XI0/MM8_d
+ N_WL<35>_XI0/XI19/XI0/MM8_g N_BLN<15>_XI0/XI19/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI0/MM5 N_XI0/XI19/XI0/NET34_XI0/XI19/XI0/MM5_d
+ N_XI0/XI19/XI0/NET33_XI0/XI19/XI0/MM5_g N_VDD_XI0/XI19/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI0/MM4 N_XI0/XI19/XI0/NET33_XI0/XI19/XI0/MM4_d
+ N_XI0/XI19/XI0/NET34_XI0/XI19/XI0/MM4_g N_VDD_XI0/XI19/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI0/MM10 N_XI0/XI19/XI0/NET35_XI0/XI19/XI0/MM10_d
+ N_XI0/XI19/XI0/NET36_XI0/XI19/XI0/MM10_g N_VDD_XI0/XI19/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI0/MM11 N_XI0/XI19/XI0/NET36_XI0/XI19/XI0/MM11_d
+ N_XI0/XI19/XI0/NET35_XI0/XI19/XI0/MM11_g N_VDD_XI0/XI19/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI1/MM2 N_XI0/XI19/XI1/NET34_XI0/XI19/XI1/MM2_d
+ N_XI0/XI19/XI1/NET33_XI0/XI19/XI1/MM2_g N_VSS_XI0/XI19/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM3 N_XI0/XI19/XI1/NET33_XI0/XI19/XI1/MM3_d
+ N_WL<34>_XI0/XI19/XI1/MM3_g N_BLN<14>_XI0/XI19/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM0 N_XI0/XI19/XI1/NET34_XI0/XI19/XI1/MM0_d
+ N_WL<34>_XI0/XI19/XI1/MM0_g N_BL<14>_XI0/XI19/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM1 N_XI0/XI19/XI1/NET33_XI0/XI19/XI1/MM1_d
+ N_XI0/XI19/XI1/NET34_XI0/XI19/XI1/MM1_g N_VSS_XI0/XI19/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM9 N_XI0/XI19/XI1/NET36_XI0/XI19/XI1/MM9_d
+ N_WL<35>_XI0/XI19/XI1/MM9_g N_BL<14>_XI0/XI19/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM6 N_XI0/XI19/XI1/NET35_XI0/XI19/XI1/MM6_d
+ N_XI0/XI19/XI1/NET36_XI0/XI19/XI1/MM6_g N_VSS_XI0/XI19/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM7 N_XI0/XI19/XI1/NET36_XI0/XI19/XI1/MM7_d
+ N_XI0/XI19/XI1/NET35_XI0/XI19/XI1/MM7_g N_VSS_XI0/XI19/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM8 N_XI0/XI19/XI1/NET35_XI0/XI19/XI1/MM8_d
+ N_WL<35>_XI0/XI19/XI1/MM8_g N_BLN<14>_XI0/XI19/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI1/MM5 N_XI0/XI19/XI1/NET34_XI0/XI19/XI1/MM5_d
+ N_XI0/XI19/XI1/NET33_XI0/XI19/XI1/MM5_g N_VDD_XI0/XI19/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI1/MM4 N_XI0/XI19/XI1/NET33_XI0/XI19/XI1/MM4_d
+ N_XI0/XI19/XI1/NET34_XI0/XI19/XI1/MM4_g N_VDD_XI0/XI19/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI1/MM10 N_XI0/XI19/XI1/NET35_XI0/XI19/XI1/MM10_d
+ N_XI0/XI19/XI1/NET36_XI0/XI19/XI1/MM10_g N_VDD_XI0/XI19/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI1/MM11 N_XI0/XI19/XI1/NET36_XI0/XI19/XI1/MM11_d
+ N_XI0/XI19/XI1/NET35_XI0/XI19/XI1/MM11_g N_VDD_XI0/XI19/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI2/MM2 N_XI0/XI19/XI2/NET34_XI0/XI19/XI2/MM2_d
+ N_XI0/XI19/XI2/NET33_XI0/XI19/XI2/MM2_g N_VSS_XI0/XI19/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM3 N_XI0/XI19/XI2/NET33_XI0/XI19/XI2/MM3_d
+ N_WL<34>_XI0/XI19/XI2/MM3_g N_BLN<13>_XI0/XI19/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM0 N_XI0/XI19/XI2/NET34_XI0/XI19/XI2/MM0_d
+ N_WL<34>_XI0/XI19/XI2/MM0_g N_BL<13>_XI0/XI19/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM1 N_XI0/XI19/XI2/NET33_XI0/XI19/XI2/MM1_d
+ N_XI0/XI19/XI2/NET34_XI0/XI19/XI2/MM1_g N_VSS_XI0/XI19/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM9 N_XI0/XI19/XI2/NET36_XI0/XI19/XI2/MM9_d
+ N_WL<35>_XI0/XI19/XI2/MM9_g N_BL<13>_XI0/XI19/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM6 N_XI0/XI19/XI2/NET35_XI0/XI19/XI2/MM6_d
+ N_XI0/XI19/XI2/NET36_XI0/XI19/XI2/MM6_g N_VSS_XI0/XI19/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM7 N_XI0/XI19/XI2/NET36_XI0/XI19/XI2/MM7_d
+ N_XI0/XI19/XI2/NET35_XI0/XI19/XI2/MM7_g N_VSS_XI0/XI19/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM8 N_XI0/XI19/XI2/NET35_XI0/XI19/XI2/MM8_d
+ N_WL<35>_XI0/XI19/XI2/MM8_g N_BLN<13>_XI0/XI19/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI2/MM5 N_XI0/XI19/XI2/NET34_XI0/XI19/XI2/MM5_d
+ N_XI0/XI19/XI2/NET33_XI0/XI19/XI2/MM5_g N_VDD_XI0/XI19/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI2/MM4 N_XI0/XI19/XI2/NET33_XI0/XI19/XI2/MM4_d
+ N_XI0/XI19/XI2/NET34_XI0/XI19/XI2/MM4_g N_VDD_XI0/XI19/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI2/MM10 N_XI0/XI19/XI2/NET35_XI0/XI19/XI2/MM10_d
+ N_XI0/XI19/XI2/NET36_XI0/XI19/XI2/MM10_g N_VDD_XI0/XI19/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI2/MM11 N_XI0/XI19/XI2/NET36_XI0/XI19/XI2/MM11_d
+ N_XI0/XI19/XI2/NET35_XI0/XI19/XI2/MM11_g N_VDD_XI0/XI19/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI3/MM2 N_XI0/XI19/XI3/NET34_XI0/XI19/XI3/MM2_d
+ N_XI0/XI19/XI3/NET33_XI0/XI19/XI3/MM2_g N_VSS_XI0/XI19/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM3 N_XI0/XI19/XI3/NET33_XI0/XI19/XI3/MM3_d
+ N_WL<34>_XI0/XI19/XI3/MM3_g N_BLN<12>_XI0/XI19/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM0 N_XI0/XI19/XI3/NET34_XI0/XI19/XI3/MM0_d
+ N_WL<34>_XI0/XI19/XI3/MM0_g N_BL<12>_XI0/XI19/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM1 N_XI0/XI19/XI3/NET33_XI0/XI19/XI3/MM1_d
+ N_XI0/XI19/XI3/NET34_XI0/XI19/XI3/MM1_g N_VSS_XI0/XI19/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM9 N_XI0/XI19/XI3/NET36_XI0/XI19/XI3/MM9_d
+ N_WL<35>_XI0/XI19/XI3/MM9_g N_BL<12>_XI0/XI19/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM6 N_XI0/XI19/XI3/NET35_XI0/XI19/XI3/MM6_d
+ N_XI0/XI19/XI3/NET36_XI0/XI19/XI3/MM6_g N_VSS_XI0/XI19/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM7 N_XI0/XI19/XI3/NET36_XI0/XI19/XI3/MM7_d
+ N_XI0/XI19/XI3/NET35_XI0/XI19/XI3/MM7_g N_VSS_XI0/XI19/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM8 N_XI0/XI19/XI3/NET35_XI0/XI19/XI3/MM8_d
+ N_WL<35>_XI0/XI19/XI3/MM8_g N_BLN<12>_XI0/XI19/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI3/MM5 N_XI0/XI19/XI3/NET34_XI0/XI19/XI3/MM5_d
+ N_XI0/XI19/XI3/NET33_XI0/XI19/XI3/MM5_g N_VDD_XI0/XI19/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI3/MM4 N_XI0/XI19/XI3/NET33_XI0/XI19/XI3/MM4_d
+ N_XI0/XI19/XI3/NET34_XI0/XI19/XI3/MM4_g N_VDD_XI0/XI19/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI3/MM10 N_XI0/XI19/XI3/NET35_XI0/XI19/XI3/MM10_d
+ N_XI0/XI19/XI3/NET36_XI0/XI19/XI3/MM10_g N_VDD_XI0/XI19/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI3/MM11 N_XI0/XI19/XI3/NET36_XI0/XI19/XI3/MM11_d
+ N_XI0/XI19/XI3/NET35_XI0/XI19/XI3/MM11_g N_VDD_XI0/XI19/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI4/MM2 N_XI0/XI19/XI4/NET34_XI0/XI19/XI4/MM2_d
+ N_XI0/XI19/XI4/NET33_XI0/XI19/XI4/MM2_g N_VSS_XI0/XI19/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM3 N_XI0/XI19/XI4/NET33_XI0/XI19/XI4/MM3_d
+ N_WL<34>_XI0/XI19/XI4/MM3_g N_BLN<11>_XI0/XI19/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM0 N_XI0/XI19/XI4/NET34_XI0/XI19/XI4/MM0_d
+ N_WL<34>_XI0/XI19/XI4/MM0_g N_BL<11>_XI0/XI19/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM1 N_XI0/XI19/XI4/NET33_XI0/XI19/XI4/MM1_d
+ N_XI0/XI19/XI4/NET34_XI0/XI19/XI4/MM1_g N_VSS_XI0/XI19/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM9 N_XI0/XI19/XI4/NET36_XI0/XI19/XI4/MM9_d
+ N_WL<35>_XI0/XI19/XI4/MM9_g N_BL<11>_XI0/XI19/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM6 N_XI0/XI19/XI4/NET35_XI0/XI19/XI4/MM6_d
+ N_XI0/XI19/XI4/NET36_XI0/XI19/XI4/MM6_g N_VSS_XI0/XI19/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM7 N_XI0/XI19/XI4/NET36_XI0/XI19/XI4/MM7_d
+ N_XI0/XI19/XI4/NET35_XI0/XI19/XI4/MM7_g N_VSS_XI0/XI19/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM8 N_XI0/XI19/XI4/NET35_XI0/XI19/XI4/MM8_d
+ N_WL<35>_XI0/XI19/XI4/MM8_g N_BLN<11>_XI0/XI19/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI4/MM5 N_XI0/XI19/XI4/NET34_XI0/XI19/XI4/MM5_d
+ N_XI0/XI19/XI4/NET33_XI0/XI19/XI4/MM5_g N_VDD_XI0/XI19/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI4/MM4 N_XI0/XI19/XI4/NET33_XI0/XI19/XI4/MM4_d
+ N_XI0/XI19/XI4/NET34_XI0/XI19/XI4/MM4_g N_VDD_XI0/XI19/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI4/MM10 N_XI0/XI19/XI4/NET35_XI0/XI19/XI4/MM10_d
+ N_XI0/XI19/XI4/NET36_XI0/XI19/XI4/MM10_g N_VDD_XI0/XI19/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI4/MM11 N_XI0/XI19/XI4/NET36_XI0/XI19/XI4/MM11_d
+ N_XI0/XI19/XI4/NET35_XI0/XI19/XI4/MM11_g N_VDD_XI0/XI19/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI5/MM2 N_XI0/XI19/XI5/NET34_XI0/XI19/XI5/MM2_d
+ N_XI0/XI19/XI5/NET33_XI0/XI19/XI5/MM2_g N_VSS_XI0/XI19/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM3 N_XI0/XI19/XI5/NET33_XI0/XI19/XI5/MM3_d
+ N_WL<34>_XI0/XI19/XI5/MM3_g N_BLN<10>_XI0/XI19/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM0 N_XI0/XI19/XI5/NET34_XI0/XI19/XI5/MM0_d
+ N_WL<34>_XI0/XI19/XI5/MM0_g N_BL<10>_XI0/XI19/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM1 N_XI0/XI19/XI5/NET33_XI0/XI19/XI5/MM1_d
+ N_XI0/XI19/XI5/NET34_XI0/XI19/XI5/MM1_g N_VSS_XI0/XI19/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM9 N_XI0/XI19/XI5/NET36_XI0/XI19/XI5/MM9_d
+ N_WL<35>_XI0/XI19/XI5/MM9_g N_BL<10>_XI0/XI19/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM6 N_XI0/XI19/XI5/NET35_XI0/XI19/XI5/MM6_d
+ N_XI0/XI19/XI5/NET36_XI0/XI19/XI5/MM6_g N_VSS_XI0/XI19/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM7 N_XI0/XI19/XI5/NET36_XI0/XI19/XI5/MM7_d
+ N_XI0/XI19/XI5/NET35_XI0/XI19/XI5/MM7_g N_VSS_XI0/XI19/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM8 N_XI0/XI19/XI5/NET35_XI0/XI19/XI5/MM8_d
+ N_WL<35>_XI0/XI19/XI5/MM8_g N_BLN<10>_XI0/XI19/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI5/MM5 N_XI0/XI19/XI5/NET34_XI0/XI19/XI5/MM5_d
+ N_XI0/XI19/XI5/NET33_XI0/XI19/XI5/MM5_g N_VDD_XI0/XI19/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI5/MM4 N_XI0/XI19/XI5/NET33_XI0/XI19/XI5/MM4_d
+ N_XI0/XI19/XI5/NET34_XI0/XI19/XI5/MM4_g N_VDD_XI0/XI19/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI5/MM10 N_XI0/XI19/XI5/NET35_XI0/XI19/XI5/MM10_d
+ N_XI0/XI19/XI5/NET36_XI0/XI19/XI5/MM10_g N_VDD_XI0/XI19/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI5/MM11 N_XI0/XI19/XI5/NET36_XI0/XI19/XI5/MM11_d
+ N_XI0/XI19/XI5/NET35_XI0/XI19/XI5/MM11_g N_VDD_XI0/XI19/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI6/MM2 N_XI0/XI19/XI6/NET34_XI0/XI19/XI6/MM2_d
+ N_XI0/XI19/XI6/NET33_XI0/XI19/XI6/MM2_g N_VSS_XI0/XI19/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM3 N_XI0/XI19/XI6/NET33_XI0/XI19/XI6/MM3_d
+ N_WL<34>_XI0/XI19/XI6/MM3_g N_BLN<9>_XI0/XI19/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM0 N_XI0/XI19/XI6/NET34_XI0/XI19/XI6/MM0_d
+ N_WL<34>_XI0/XI19/XI6/MM0_g N_BL<9>_XI0/XI19/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM1 N_XI0/XI19/XI6/NET33_XI0/XI19/XI6/MM1_d
+ N_XI0/XI19/XI6/NET34_XI0/XI19/XI6/MM1_g N_VSS_XI0/XI19/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM9 N_XI0/XI19/XI6/NET36_XI0/XI19/XI6/MM9_d
+ N_WL<35>_XI0/XI19/XI6/MM9_g N_BL<9>_XI0/XI19/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM6 N_XI0/XI19/XI6/NET35_XI0/XI19/XI6/MM6_d
+ N_XI0/XI19/XI6/NET36_XI0/XI19/XI6/MM6_g N_VSS_XI0/XI19/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM7 N_XI0/XI19/XI6/NET36_XI0/XI19/XI6/MM7_d
+ N_XI0/XI19/XI6/NET35_XI0/XI19/XI6/MM7_g N_VSS_XI0/XI19/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM8 N_XI0/XI19/XI6/NET35_XI0/XI19/XI6/MM8_d
+ N_WL<35>_XI0/XI19/XI6/MM8_g N_BLN<9>_XI0/XI19/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI6/MM5 N_XI0/XI19/XI6/NET34_XI0/XI19/XI6/MM5_d
+ N_XI0/XI19/XI6/NET33_XI0/XI19/XI6/MM5_g N_VDD_XI0/XI19/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI6/MM4 N_XI0/XI19/XI6/NET33_XI0/XI19/XI6/MM4_d
+ N_XI0/XI19/XI6/NET34_XI0/XI19/XI6/MM4_g N_VDD_XI0/XI19/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI6/MM10 N_XI0/XI19/XI6/NET35_XI0/XI19/XI6/MM10_d
+ N_XI0/XI19/XI6/NET36_XI0/XI19/XI6/MM10_g N_VDD_XI0/XI19/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI6/MM11 N_XI0/XI19/XI6/NET36_XI0/XI19/XI6/MM11_d
+ N_XI0/XI19/XI6/NET35_XI0/XI19/XI6/MM11_g N_VDD_XI0/XI19/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI7/MM2 N_XI0/XI19/XI7/NET34_XI0/XI19/XI7/MM2_d
+ N_XI0/XI19/XI7/NET33_XI0/XI19/XI7/MM2_g N_VSS_XI0/XI19/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM3 N_XI0/XI19/XI7/NET33_XI0/XI19/XI7/MM3_d
+ N_WL<34>_XI0/XI19/XI7/MM3_g N_BLN<8>_XI0/XI19/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM0 N_XI0/XI19/XI7/NET34_XI0/XI19/XI7/MM0_d
+ N_WL<34>_XI0/XI19/XI7/MM0_g N_BL<8>_XI0/XI19/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM1 N_XI0/XI19/XI7/NET33_XI0/XI19/XI7/MM1_d
+ N_XI0/XI19/XI7/NET34_XI0/XI19/XI7/MM1_g N_VSS_XI0/XI19/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM9 N_XI0/XI19/XI7/NET36_XI0/XI19/XI7/MM9_d
+ N_WL<35>_XI0/XI19/XI7/MM9_g N_BL<8>_XI0/XI19/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM6 N_XI0/XI19/XI7/NET35_XI0/XI19/XI7/MM6_d
+ N_XI0/XI19/XI7/NET36_XI0/XI19/XI7/MM6_g N_VSS_XI0/XI19/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM7 N_XI0/XI19/XI7/NET36_XI0/XI19/XI7/MM7_d
+ N_XI0/XI19/XI7/NET35_XI0/XI19/XI7/MM7_g N_VSS_XI0/XI19/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM8 N_XI0/XI19/XI7/NET35_XI0/XI19/XI7/MM8_d
+ N_WL<35>_XI0/XI19/XI7/MM8_g N_BLN<8>_XI0/XI19/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI7/MM5 N_XI0/XI19/XI7/NET34_XI0/XI19/XI7/MM5_d
+ N_XI0/XI19/XI7/NET33_XI0/XI19/XI7/MM5_g N_VDD_XI0/XI19/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI7/MM4 N_XI0/XI19/XI7/NET33_XI0/XI19/XI7/MM4_d
+ N_XI0/XI19/XI7/NET34_XI0/XI19/XI7/MM4_g N_VDD_XI0/XI19/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI7/MM10 N_XI0/XI19/XI7/NET35_XI0/XI19/XI7/MM10_d
+ N_XI0/XI19/XI7/NET36_XI0/XI19/XI7/MM10_g N_VDD_XI0/XI19/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI7/MM11 N_XI0/XI19/XI7/NET36_XI0/XI19/XI7/MM11_d
+ N_XI0/XI19/XI7/NET35_XI0/XI19/XI7/MM11_g N_VDD_XI0/XI19/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI8/MM2 N_XI0/XI19/XI8/NET34_XI0/XI19/XI8/MM2_d
+ N_XI0/XI19/XI8/NET33_XI0/XI19/XI8/MM2_g N_VSS_XI0/XI19/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM3 N_XI0/XI19/XI8/NET33_XI0/XI19/XI8/MM3_d
+ N_WL<34>_XI0/XI19/XI8/MM3_g N_BLN<7>_XI0/XI19/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM0 N_XI0/XI19/XI8/NET34_XI0/XI19/XI8/MM0_d
+ N_WL<34>_XI0/XI19/XI8/MM0_g N_BL<7>_XI0/XI19/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM1 N_XI0/XI19/XI8/NET33_XI0/XI19/XI8/MM1_d
+ N_XI0/XI19/XI8/NET34_XI0/XI19/XI8/MM1_g N_VSS_XI0/XI19/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM9 N_XI0/XI19/XI8/NET36_XI0/XI19/XI8/MM9_d
+ N_WL<35>_XI0/XI19/XI8/MM9_g N_BL<7>_XI0/XI19/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM6 N_XI0/XI19/XI8/NET35_XI0/XI19/XI8/MM6_d
+ N_XI0/XI19/XI8/NET36_XI0/XI19/XI8/MM6_g N_VSS_XI0/XI19/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM7 N_XI0/XI19/XI8/NET36_XI0/XI19/XI8/MM7_d
+ N_XI0/XI19/XI8/NET35_XI0/XI19/XI8/MM7_g N_VSS_XI0/XI19/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM8 N_XI0/XI19/XI8/NET35_XI0/XI19/XI8/MM8_d
+ N_WL<35>_XI0/XI19/XI8/MM8_g N_BLN<7>_XI0/XI19/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI8/MM5 N_XI0/XI19/XI8/NET34_XI0/XI19/XI8/MM5_d
+ N_XI0/XI19/XI8/NET33_XI0/XI19/XI8/MM5_g N_VDD_XI0/XI19/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI8/MM4 N_XI0/XI19/XI8/NET33_XI0/XI19/XI8/MM4_d
+ N_XI0/XI19/XI8/NET34_XI0/XI19/XI8/MM4_g N_VDD_XI0/XI19/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI8/MM10 N_XI0/XI19/XI8/NET35_XI0/XI19/XI8/MM10_d
+ N_XI0/XI19/XI8/NET36_XI0/XI19/XI8/MM10_g N_VDD_XI0/XI19/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI8/MM11 N_XI0/XI19/XI8/NET36_XI0/XI19/XI8/MM11_d
+ N_XI0/XI19/XI8/NET35_XI0/XI19/XI8/MM11_g N_VDD_XI0/XI19/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI9/MM2 N_XI0/XI19/XI9/NET34_XI0/XI19/XI9/MM2_d
+ N_XI0/XI19/XI9/NET33_XI0/XI19/XI9/MM2_g N_VSS_XI0/XI19/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM3 N_XI0/XI19/XI9/NET33_XI0/XI19/XI9/MM3_d
+ N_WL<34>_XI0/XI19/XI9/MM3_g N_BLN<6>_XI0/XI19/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM0 N_XI0/XI19/XI9/NET34_XI0/XI19/XI9/MM0_d
+ N_WL<34>_XI0/XI19/XI9/MM0_g N_BL<6>_XI0/XI19/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM1 N_XI0/XI19/XI9/NET33_XI0/XI19/XI9/MM1_d
+ N_XI0/XI19/XI9/NET34_XI0/XI19/XI9/MM1_g N_VSS_XI0/XI19/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM9 N_XI0/XI19/XI9/NET36_XI0/XI19/XI9/MM9_d
+ N_WL<35>_XI0/XI19/XI9/MM9_g N_BL<6>_XI0/XI19/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM6 N_XI0/XI19/XI9/NET35_XI0/XI19/XI9/MM6_d
+ N_XI0/XI19/XI9/NET36_XI0/XI19/XI9/MM6_g N_VSS_XI0/XI19/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM7 N_XI0/XI19/XI9/NET36_XI0/XI19/XI9/MM7_d
+ N_XI0/XI19/XI9/NET35_XI0/XI19/XI9/MM7_g N_VSS_XI0/XI19/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM8 N_XI0/XI19/XI9/NET35_XI0/XI19/XI9/MM8_d
+ N_WL<35>_XI0/XI19/XI9/MM8_g N_BLN<6>_XI0/XI19/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI9/MM5 N_XI0/XI19/XI9/NET34_XI0/XI19/XI9/MM5_d
+ N_XI0/XI19/XI9/NET33_XI0/XI19/XI9/MM5_g N_VDD_XI0/XI19/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI9/MM4 N_XI0/XI19/XI9/NET33_XI0/XI19/XI9/MM4_d
+ N_XI0/XI19/XI9/NET34_XI0/XI19/XI9/MM4_g N_VDD_XI0/XI19/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI9/MM10 N_XI0/XI19/XI9/NET35_XI0/XI19/XI9/MM10_d
+ N_XI0/XI19/XI9/NET36_XI0/XI19/XI9/MM10_g N_VDD_XI0/XI19/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI9/MM11 N_XI0/XI19/XI9/NET36_XI0/XI19/XI9/MM11_d
+ N_XI0/XI19/XI9/NET35_XI0/XI19/XI9/MM11_g N_VDD_XI0/XI19/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI10/MM2 N_XI0/XI19/XI10/NET34_XI0/XI19/XI10/MM2_d
+ N_XI0/XI19/XI10/NET33_XI0/XI19/XI10/MM2_g N_VSS_XI0/XI19/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM3 N_XI0/XI19/XI10/NET33_XI0/XI19/XI10/MM3_d
+ N_WL<34>_XI0/XI19/XI10/MM3_g N_BLN<5>_XI0/XI19/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM0 N_XI0/XI19/XI10/NET34_XI0/XI19/XI10/MM0_d
+ N_WL<34>_XI0/XI19/XI10/MM0_g N_BL<5>_XI0/XI19/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM1 N_XI0/XI19/XI10/NET33_XI0/XI19/XI10/MM1_d
+ N_XI0/XI19/XI10/NET34_XI0/XI19/XI10/MM1_g N_VSS_XI0/XI19/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM9 N_XI0/XI19/XI10/NET36_XI0/XI19/XI10/MM9_d
+ N_WL<35>_XI0/XI19/XI10/MM9_g N_BL<5>_XI0/XI19/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM6 N_XI0/XI19/XI10/NET35_XI0/XI19/XI10/MM6_d
+ N_XI0/XI19/XI10/NET36_XI0/XI19/XI10/MM6_g N_VSS_XI0/XI19/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM7 N_XI0/XI19/XI10/NET36_XI0/XI19/XI10/MM7_d
+ N_XI0/XI19/XI10/NET35_XI0/XI19/XI10/MM7_g N_VSS_XI0/XI19/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM8 N_XI0/XI19/XI10/NET35_XI0/XI19/XI10/MM8_d
+ N_WL<35>_XI0/XI19/XI10/MM8_g N_BLN<5>_XI0/XI19/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI10/MM5 N_XI0/XI19/XI10/NET34_XI0/XI19/XI10/MM5_d
+ N_XI0/XI19/XI10/NET33_XI0/XI19/XI10/MM5_g N_VDD_XI0/XI19/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI10/MM4 N_XI0/XI19/XI10/NET33_XI0/XI19/XI10/MM4_d
+ N_XI0/XI19/XI10/NET34_XI0/XI19/XI10/MM4_g N_VDD_XI0/XI19/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI10/MM10 N_XI0/XI19/XI10/NET35_XI0/XI19/XI10/MM10_d
+ N_XI0/XI19/XI10/NET36_XI0/XI19/XI10/MM10_g N_VDD_XI0/XI19/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI10/MM11 N_XI0/XI19/XI10/NET36_XI0/XI19/XI10/MM11_d
+ N_XI0/XI19/XI10/NET35_XI0/XI19/XI10/MM11_g N_VDD_XI0/XI19/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI11/MM2 N_XI0/XI19/XI11/NET34_XI0/XI19/XI11/MM2_d
+ N_XI0/XI19/XI11/NET33_XI0/XI19/XI11/MM2_g N_VSS_XI0/XI19/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM3 N_XI0/XI19/XI11/NET33_XI0/XI19/XI11/MM3_d
+ N_WL<34>_XI0/XI19/XI11/MM3_g N_BLN<4>_XI0/XI19/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM0 N_XI0/XI19/XI11/NET34_XI0/XI19/XI11/MM0_d
+ N_WL<34>_XI0/XI19/XI11/MM0_g N_BL<4>_XI0/XI19/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM1 N_XI0/XI19/XI11/NET33_XI0/XI19/XI11/MM1_d
+ N_XI0/XI19/XI11/NET34_XI0/XI19/XI11/MM1_g N_VSS_XI0/XI19/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM9 N_XI0/XI19/XI11/NET36_XI0/XI19/XI11/MM9_d
+ N_WL<35>_XI0/XI19/XI11/MM9_g N_BL<4>_XI0/XI19/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM6 N_XI0/XI19/XI11/NET35_XI0/XI19/XI11/MM6_d
+ N_XI0/XI19/XI11/NET36_XI0/XI19/XI11/MM6_g N_VSS_XI0/XI19/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM7 N_XI0/XI19/XI11/NET36_XI0/XI19/XI11/MM7_d
+ N_XI0/XI19/XI11/NET35_XI0/XI19/XI11/MM7_g N_VSS_XI0/XI19/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM8 N_XI0/XI19/XI11/NET35_XI0/XI19/XI11/MM8_d
+ N_WL<35>_XI0/XI19/XI11/MM8_g N_BLN<4>_XI0/XI19/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI11/MM5 N_XI0/XI19/XI11/NET34_XI0/XI19/XI11/MM5_d
+ N_XI0/XI19/XI11/NET33_XI0/XI19/XI11/MM5_g N_VDD_XI0/XI19/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI11/MM4 N_XI0/XI19/XI11/NET33_XI0/XI19/XI11/MM4_d
+ N_XI0/XI19/XI11/NET34_XI0/XI19/XI11/MM4_g N_VDD_XI0/XI19/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI11/MM10 N_XI0/XI19/XI11/NET35_XI0/XI19/XI11/MM10_d
+ N_XI0/XI19/XI11/NET36_XI0/XI19/XI11/MM10_g N_VDD_XI0/XI19/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI11/MM11 N_XI0/XI19/XI11/NET36_XI0/XI19/XI11/MM11_d
+ N_XI0/XI19/XI11/NET35_XI0/XI19/XI11/MM11_g N_VDD_XI0/XI19/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI12/MM2 N_XI0/XI19/XI12/NET34_XI0/XI19/XI12/MM2_d
+ N_XI0/XI19/XI12/NET33_XI0/XI19/XI12/MM2_g N_VSS_XI0/XI19/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM3 N_XI0/XI19/XI12/NET33_XI0/XI19/XI12/MM3_d
+ N_WL<34>_XI0/XI19/XI12/MM3_g N_BLN<3>_XI0/XI19/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM0 N_XI0/XI19/XI12/NET34_XI0/XI19/XI12/MM0_d
+ N_WL<34>_XI0/XI19/XI12/MM0_g N_BL<3>_XI0/XI19/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM1 N_XI0/XI19/XI12/NET33_XI0/XI19/XI12/MM1_d
+ N_XI0/XI19/XI12/NET34_XI0/XI19/XI12/MM1_g N_VSS_XI0/XI19/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM9 N_XI0/XI19/XI12/NET36_XI0/XI19/XI12/MM9_d
+ N_WL<35>_XI0/XI19/XI12/MM9_g N_BL<3>_XI0/XI19/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM6 N_XI0/XI19/XI12/NET35_XI0/XI19/XI12/MM6_d
+ N_XI0/XI19/XI12/NET36_XI0/XI19/XI12/MM6_g N_VSS_XI0/XI19/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM7 N_XI0/XI19/XI12/NET36_XI0/XI19/XI12/MM7_d
+ N_XI0/XI19/XI12/NET35_XI0/XI19/XI12/MM7_g N_VSS_XI0/XI19/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM8 N_XI0/XI19/XI12/NET35_XI0/XI19/XI12/MM8_d
+ N_WL<35>_XI0/XI19/XI12/MM8_g N_BLN<3>_XI0/XI19/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI12/MM5 N_XI0/XI19/XI12/NET34_XI0/XI19/XI12/MM5_d
+ N_XI0/XI19/XI12/NET33_XI0/XI19/XI12/MM5_g N_VDD_XI0/XI19/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI12/MM4 N_XI0/XI19/XI12/NET33_XI0/XI19/XI12/MM4_d
+ N_XI0/XI19/XI12/NET34_XI0/XI19/XI12/MM4_g N_VDD_XI0/XI19/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI12/MM10 N_XI0/XI19/XI12/NET35_XI0/XI19/XI12/MM10_d
+ N_XI0/XI19/XI12/NET36_XI0/XI19/XI12/MM10_g N_VDD_XI0/XI19/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI12/MM11 N_XI0/XI19/XI12/NET36_XI0/XI19/XI12/MM11_d
+ N_XI0/XI19/XI12/NET35_XI0/XI19/XI12/MM11_g N_VDD_XI0/XI19/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI13/MM2 N_XI0/XI19/XI13/NET34_XI0/XI19/XI13/MM2_d
+ N_XI0/XI19/XI13/NET33_XI0/XI19/XI13/MM2_g N_VSS_XI0/XI19/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM3 N_XI0/XI19/XI13/NET33_XI0/XI19/XI13/MM3_d
+ N_WL<34>_XI0/XI19/XI13/MM3_g N_BLN<2>_XI0/XI19/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM0 N_XI0/XI19/XI13/NET34_XI0/XI19/XI13/MM0_d
+ N_WL<34>_XI0/XI19/XI13/MM0_g N_BL<2>_XI0/XI19/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM1 N_XI0/XI19/XI13/NET33_XI0/XI19/XI13/MM1_d
+ N_XI0/XI19/XI13/NET34_XI0/XI19/XI13/MM1_g N_VSS_XI0/XI19/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM9 N_XI0/XI19/XI13/NET36_XI0/XI19/XI13/MM9_d
+ N_WL<35>_XI0/XI19/XI13/MM9_g N_BL<2>_XI0/XI19/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM6 N_XI0/XI19/XI13/NET35_XI0/XI19/XI13/MM6_d
+ N_XI0/XI19/XI13/NET36_XI0/XI19/XI13/MM6_g N_VSS_XI0/XI19/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM7 N_XI0/XI19/XI13/NET36_XI0/XI19/XI13/MM7_d
+ N_XI0/XI19/XI13/NET35_XI0/XI19/XI13/MM7_g N_VSS_XI0/XI19/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM8 N_XI0/XI19/XI13/NET35_XI0/XI19/XI13/MM8_d
+ N_WL<35>_XI0/XI19/XI13/MM8_g N_BLN<2>_XI0/XI19/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI13/MM5 N_XI0/XI19/XI13/NET34_XI0/XI19/XI13/MM5_d
+ N_XI0/XI19/XI13/NET33_XI0/XI19/XI13/MM5_g N_VDD_XI0/XI19/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI13/MM4 N_XI0/XI19/XI13/NET33_XI0/XI19/XI13/MM4_d
+ N_XI0/XI19/XI13/NET34_XI0/XI19/XI13/MM4_g N_VDD_XI0/XI19/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI13/MM10 N_XI0/XI19/XI13/NET35_XI0/XI19/XI13/MM10_d
+ N_XI0/XI19/XI13/NET36_XI0/XI19/XI13/MM10_g N_VDD_XI0/XI19/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI13/MM11 N_XI0/XI19/XI13/NET36_XI0/XI19/XI13/MM11_d
+ N_XI0/XI19/XI13/NET35_XI0/XI19/XI13/MM11_g N_VDD_XI0/XI19/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI14/MM2 N_XI0/XI19/XI14/NET34_XI0/XI19/XI14/MM2_d
+ N_XI0/XI19/XI14/NET33_XI0/XI19/XI14/MM2_g N_VSS_XI0/XI19/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM3 N_XI0/XI19/XI14/NET33_XI0/XI19/XI14/MM3_d
+ N_WL<34>_XI0/XI19/XI14/MM3_g N_BLN<1>_XI0/XI19/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM0 N_XI0/XI19/XI14/NET34_XI0/XI19/XI14/MM0_d
+ N_WL<34>_XI0/XI19/XI14/MM0_g N_BL<1>_XI0/XI19/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM1 N_XI0/XI19/XI14/NET33_XI0/XI19/XI14/MM1_d
+ N_XI0/XI19/XI14/NET34_XI0/XI19/XI14/MM1_g N_VSS_XI0/XI19/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM9 N_XI0/XI19/XI14/NET36_XI0/XI19/XI14/MM9_d
+ N_WL<35>_XI0/XI19/XI14/MM9_g N_BL<1>_XI0/XI19/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM6 N_XI0/XI19/XI14/NET35_XI0/XI19/XI14/MM6_d
+ N_XI0/XI19/XI14/NET36_XI0/XI19/XI14/MM6_g N_VSS_XI0/XI19/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM7 N_XI0/XI19/XI14/NET36_XI0/XI19/XI14/MM7_d
+ N_XI0/XI19/XI14/NET35_XI0/XI19/XI14/MM7_g N_VSS_XI0/XI19/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM8 N_XI0/XI19/XI14/NET35_XI0/XI19/XI14/MM8_d
+ N_WL<35>_XI0/XI19/XI14/MM8_g N_BLN<1>_XI0/XI19/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI14/MM5 N_XI0/XI19/XI14/NET34_XI0/XI19/XI14/MM5_d
+ N_XI0/XI19/XI14/NET33_XI0/XI19/XI14/MM5_g N_VDD_XI0/XI19/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI14/MM4 N_XI0/XI19/XI14/NET33_XI0/XI19/XI14/MM4_d
+ N_XI0/XI19/XI14/NET34_XI0/XI19/XI14/MM4_g N_VDD_XI0/XI19/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI14/MM10 N_XI0/XI19/XI14/NET35_XI0/XI19/XI14/MM10_d
+ N_XI0/XI19/XI14/NET36_XI0/XI19/XI14/MM10_g N_VDD_XI0/XI19/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI14/MM11 N_XI0/XI19/XI14/NET36_XI0/XI19/XI14/MM11_d
+ N_XI0/XI19/XI14/NET35_XI0/XI19/XI14/MM11_g N_VDD_XI0/XI19/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI15/MM2 N_XI0/XI19/XI15/NET34_XI0/XI19/XI15/MM2_d
+ N_XI0/XI19/XI15/NET33_XI0/XI19/XI15/MM2_g N_VSS_XI0/XI19/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM3 N_XI0/XI19/XI15/NET33_XI0/XI19/XI15/MM3_d
+ N_WL<34>_XI0/XI19/XI15/MM3_g N_BLN<0>_XI0/XI19/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM0 N_XI0/XI19/XI15/NET34_XI0/XI19/XI15/MM0_d
+ N_WL<34>_XI0/XI19/XI15/MM0_g N_BL<0>_XI0/XI19/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM1 N_XI0/XI19/XI15/NET33_XI0/XI19/XI15/MM1_d
+ N_XI0/XI19/XI15/NET34_XI0/XI19/XI15/MM1_g N_VSS_XI0/XI19/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM9 N_XI0/XI19/XI15/NET36_XI0/XI19/XI15/MM9_d
+ N_WL<35>_XI0/XI19/XI15/MM9_g N_BL<0>_XI0/XI19/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM6 N_XI0/XI19/XI15/NET35_XI0/XI19/XI15/MM6_d
+ N_XI0/XI19/XI15/NET36_XI0/XI19/XI15/MM6_g N_VSS_XI0/XI19/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM7 N_XI0/XI19/XI15/NET36_XI0/XI19/XI15/MM7_d
+ N_XI0/XI19/XI15/NET35_XI0/XI19/XI15/MM7_g N_VSS_XI0/XI19/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM8 N_XI0/XI19/XI15/NET35_XI0/XI19/XI15/MM8_d
+ N_WL<35>_XI0/XI19/XI15/MM8_g N_BLN<0>_XI0/XI19/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI19/XI15/MM5 N_XI0/XI19/XI15/NET34_XI0/XI19/XI15/MM5_d
+ N_XI0/XI19/XI15/NET33_XI0/XI19/XI15/MM5_g N_VDD_XI0/XI19/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI15/MM4 N_XI0/XI19/XI15/NET33_XI0/XI19/XI15/MM4_d
+ N_XI0/XI19/XI15/NET34_XI0/XI19/XI15/MM4_g N_VDD_XI0/XI19/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI15/MM10 N_XI0/XI19/XI15/NET35_XI0/XI19/XI15/MM10_d
+ N_XI0/XI19/XI15/NET36_XI0/XI19/XI15/MM10_g N_VDD_XI0/XI19/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI19/XI15/MM11 N_XI0/XI19/XI15/NET36_XI0/XI19/XI15/MM11_d
+ N_XI0/XI19/XI15/NET35_XI0/XI19/XI15/MM11_g N_VDD_XI0/XI19/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI0/MM2 N_XI0/XI20/XI0/NET34_XI0/XI20/XI0/MM2_d
+ N_XI0/XI20/XI0/NET33_XI0/XI20/XI0/MM2_g N_VSS_XI0/XI20/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM3 N_XI0/XI20/XI0/NET33_XI0/XI20/XI0/MM3_d
+ N_WL<36>_XI0/XI20/XI0/MM3_g N_BLN<15>_XI0/XI20/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM0 N_XI0/XI20/XI0/NET34_XI0/XI20/XI0/MM0_d
+ N_WL<36>_XI0/XI20/XI0/MM0_g N_BL<15>_XI0/XI20/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM1 N_XI0/XI20/XI0/NET33_XI0/XI20/XI0/MM1_d
+ N_XI0/XI20/XI0/NET34_XI0/XI20/XI0/MM1_g N_VSS_XI0/XI20/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM9 N_XI0/XI20/XI0/NET36_XI0/XI20/XI0/MM9_d
+ N_WL<37>_XI0/XI20/XI0/MM9_g N_BL<15>_XI0/XI20/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM6 N_XI0/XI20/XI0/NET35_XI0/XI20/XI0/MM6_d
+ N_XI0/XI20/XI0/NET36_XI0/XI20/XI0/MM6_g N_VSS_XI0/XI20/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM7 N_XI0/XI20/XI0/NET36_XI0/XI20/XI0/MM7_d
+ N_XI0/XI20/XI0/NET35_XI0/XI20/XI0/MM7_g N_VSS_XI0/XI20/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM8 N_XI0/XI20/XI0/NET35_XI0/XI20/XI0/MM8_d
+ N_WL<37>_XI0/XI20/XI0/MM8_g N_BLN<15>_XI0/XI20/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI0/MM5 N_XI0/XI20/XI0/NET34_XI0/XI20/XI0/MM5_d
+ N_XI0/XI20/XI0/NET33_XI0/XI20/XI0/MM5_g N_VDD_XI0/XI20/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI0/MM4 N_XI0/XI20/XI0/NET33_XI0/XI20/XI0/MM4_d
+ N_XI0/XI20/XI0/NET34_XI0/XI20/XI0/MM4_g N_VDD_XI0/XI20/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI0/MM10 N_XI0/XI20/XI0/NET35_XI0/XI20/XI0/MM10_d
+ N_XI0/XI20/XI0/NET36_XI0/XI20/XI0/MM10_g N_VDD_XI0/XI20/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI0/MM11 N_XI0/XI20/XI0/NET36_XI0/XI20/XI0/MM11_d
+ N_XI0/XI20/XI0/NET35_XI0/XI20/XI0/MM11_g N_VDD_XI0/XI20/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI1/MM2 N_XI0/XI20/XI1/NET34_XI0/XI20/XI1/MM2_d
+ N_XI0/XI20/XI1/NET33_XI0/XI20/XI1/MM2_g N_VSS_XI0/XI20/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM3 N_XI0/XI20/XI1/NET33_XI0/XI20/XI1/MM3_d
+ N_WL<36>_XI0/XI20/XI1/MM3_g N_BLN<14>_XI0/XI20/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM0 N_XI0/XI20/XI1/NET34_XI0/XI20/XI1/MM0_d
+ N_WL<36>_XI0/XI20/XI1/MM0_g N_BL<14>_XI0/XI20/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM1 N_XI0/XI20/XI1/NET33_XI0/XI20/XI1/MM1_d
+ N_XI0/XI20/XI1/NET34_XI0/XI20/XI1/MM1_g N_VSS_XI0/XI20/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM9 N_XI0/XI20/XI1/NET36_XI0/XI20/XI1/MM9_d
+ N_WL<37>_XI0/XI20/XI1/MM9_g N_BL<14>_XI0/XI20/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM6 N_XI0/XI20/XI1/NET35_XI0/XI20/XI1/MM6_d
+ N_XI0/XI20/XI1/NET36_XI0/XI20/XI1/MM6_g N_VSS_XI0/XI20/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM7 N_XI0/XI20/XI1/NET36_XI0/XI20/XI1/MM7_d
+ N_XI0/XI20/XI1/NET35_XI0/XI20/XI1/MM7_g N_VSS_XI0/XI20/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM8 N_XI0/XI20/XI1/NET35_XI0/XI20/XI1/MM8_d
+ N_WL<37>_XI0/XI20/XI1/MM8_g N_BLN<14>_XI0/XI20/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI1/MM5 N_XI0/XI20/XI1/NET34_XI0/XI20/XI1/MM5_d
+ N_XI0/XI20/XI1/NET33_XI0/XI20/XI1/MM5_g N_VDD_XI0/XI20/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI1/MM4 N_XI0/XI20/XI1/NET33_XI0/XI20/XI1/MM4_d
+ N_XI0/XI20/XI1/NET34_XI0/XI20/XI1/MM4_g N_VDD_XI0/XI20/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI1/MM10 N_XI0/XI20/XI1/NET35_XI0/XI20/XI1/MM10_d
+ N_XI0/XI20/XI1/NET36_XI0/XI20/XI1/MM10_g N_VDD_XI0/XI20/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI1/MM11 N_XI0/XI20/XI1/NET36_XI0/XI20/XI1/MM11_d
+ N_XI0/XI20/XI1/NET35_XI0/XI20/XI1/MM11_g N_VDD_XI0/XI20/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI2/MM2 N_XI0/XI20/XI2/NET34_XI0/XI20/XI2/MM2_d
+ N_XI0/XI20/XI2/NET33_XI0/XI20/XI2/MM2_g N_VSS_XI0/XI20/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM3 N_XI0/XI20/XI2/NET33_XI0/XI20/XI2/MM3_d
+ N_WL<36>_XI0/XI20/XI2/MM3_g N_BLN<13>_XI0/XI20/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM0 N_XI0/XI20/XI2/NET34_XI0/XI20/XI2/MM0_d
+ N_WL<36>_XI0/XI20/XI2/MM0_g N_BL<13>_XI0/XI20/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM1 N_XI0/XI20/XI2/NET33_XI0/XI20/XI2/MM1_d
+ N_XI0/XI20/XI2/NET34_XI0/XI20/XI2/MM1_g N_VSS_XI0/XI20/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM9 N_XI0/XI20/XI2/NET36_XI0/XI20/XI2/MM9_d
+ N_WL<37>_XI0/XI20/XI2/MM9_g N_BL<13>_XI0/XI20/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM6 N_XI0/XI20/XI2/NET35_XI0/XI20/XI2/MM6_d
+ N_XI0/XI20/XI2/NET36_XI0/XI20/XI2/MM6_g N_VSS_XI0/XI20/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM7 N_XI0/XI20/XI2/NET36_XI0/XI20/XI2/MM7_d
+ N_XI0/XI20/XI2/NET35_XI0/XI20/XI2/MM7_g N_VSS_XI0/XI20/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM8 N_XI0/XI20/XI2/NET35_XI0/XI20/XI2/MM8_d
+ N_WL<37>_XI0/XI20/XI2/MM8_g N_BLN<13>_XI0/XI20/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI2/MM5 N_XI0/XI20/XI2/NET34_XI0/XI20/XI2/MM5_d
+ N_XI0/XI20/XI2/NET33_XI0/XI20/XI2/MM5_g N_VDD_XI0/XI20/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI2/MM4 N_XI0/XI20/XI2/NET33_XI0/XI20/XI2/MM4_d
+ N_XI0/XI20/XI2/NET34_XI0/XI20/XI2/MM4_g N_VDD_XI0/XI20/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI2/MM10 N_XI0/XI20/XI2/NET35_XI0/XI20/XI2/MM10_d
+ N_XI0/XI20/XI2/NET36_XI0/XI20/XI2/MM10_g N_VDD_XI0/XI20/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI2/MM11 N_XI0/XI20/XI2/NET36_XI0/XI20/XI2/MM11_d
+ N_XI0/XI20/XI2/NET35_XI0/XI20/XI2/MM11_g N_VDD_XI0/XI20/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI3/MM2 N_XI0/XI20/XI3/NET34_XI0/XI20/XI3/MM2_d
+ N_XI0/XI20/XI3/NET33_XI0/XI20/XI3/MM2_g N_VSS_XI0/XI20/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM3 N_XI0/XI20/XI3/NET33_XI0/XI20/XI3/MM3_d
+ N_WL<36>_XI0/XI20/XI3/MM3_g N_BLN<12>_XI0/XI20/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM0 N_XI0/XI20/XI3/NET34_XI0/XI20/XI3/MM0_d
+ N_WL<36>_XI0/XI20/XI3/MM0_g N_BL<12>_XI0/XI20/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM1 N_XI0/XI20/XI3/NET33_XI0/XI20/XI3/MM1_d
+ N_XI0/XI20/XI3/NET34_XI0/XI20/XI3/MM1_g N_VSS_XI0/XI20/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM9 N_XI0/XI20/XI3/NET36_XI0/XI20/XI3/MM9_d
+ N_WL<37>_XI0/XI20/XI3/MM9_g N_BL<12>_XI0/XI20/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM6 N_XI0/XI20/XI3/NET35_XI0/XI20/XI3/MM6_d
+ N_XI0/XI20/XI3/NET36_XI0/XI20/XI3/MM6_g N_VSS_XI0/XI20/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM7 N_XI0/XI20/XI3/NET36_XI0/XI20/XI3/MM7_d
+ N_XI0/XI20/XI3/NET35_XI0/XI20/XI3/MM7_g N_VSS_XI0/XI20/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM8 N_XI0/XI20/XI3/NET35_XI0/XI20/XI3/MM8_d
+ N_WL<37>_XI0/XI20/XI3/MM8_g N_BLN<12>_XI0/XI20/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI3/MM5 N_XI0/XI20/XI3/NET34_XI0/XI20/XI3/MM5_d
+ N_XI0/XI20/XI3/NET33_XI0/XI20/XI3/MM5_g N_VDD_XI0/XI20/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI3/MM4 N_XI0/XI20/XI3/NET33_XI0/XI20/XI3/MM4_d
+ N_XI0/XI20/XI3/NET34_XI0/XI20/XI3/MM4_g N_VDD_XI0/XI20/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI3/MM10 N_XI0/XI20/XI3/NET35_XI0/XI20/XI3/MM10_d
+ N_XI0/XI20/XI3/NET36_XI0/XI20/XI3/MM10_g N_VDD_XI0/XI20/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI3/MM11 N_XI0/XI20/XI3/NET36_XI0/XI20/XI3/MM11_d
+ N_XI0/XI20/XI3/NET35_XI0/XI20/XI3/MM11_g N_VDD_XI0/XI20/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI4/MM2 N_XI0/XI20/XI4/NET34_XI0/XI20/XI4/MM2_d
+ N_XI0/XI20/XI4/NET33_XI0/XI20/XI4/MM2_g N_VSS_XI0/XI20/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM3 N_XI0/XI20/XI4/NET33_XI0/XI20/XI4/MM3_d
+ N_WL<36>_XI0/XI20/XI4/MM3_g N_BLN<11>_XI0/XI20/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM0 N_XI0/XI20/XI4/NET34_XI0/XI20/XI4/MM0_d
+ N_WL<36>_XI0/XI20/XI4/MM0_g N_BL<11>_XI0/XI20/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM1 N_XI0/XI20/XI4/NET33_XI0/XI20/XI4/MM1_d
+ N_XI0/XI20/XI4/NET34_XI0/XI20/XI4/MM1_g N_VSS_XI0/XI20/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM9 N_XI0/XI20/XI4/NET36_XI0/XI20/XI4/MM9_d
+ N_WL<37>_XI0/XI20/XI4/MM9_g N_BL<11>_XI0/XI20/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM6 N_XI0/XI20/XI4/NET35_XI0/XI20/XI4/MM6_d
+ N_XI0/XI20/XI4/NET36_XI0/XI20/XI4/MM6_g N_VSS_XI0/XI20/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM7 N_XI0/XI20/XI4/NET36_XI0/XI20/XI4/MM7_d
+ N_XI0/XI20/XI4/NET35_XI0/XI20/XI4/MM7_g N_VSS_XI0/XI20/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM8 N_XI0/XI20/XI4/NET35_XI0/XI20/XI4/MM8_d
+ N_WL<37>_XI0/XI20/XI4/MM8_g N_BLN<11>_XI0/XI20/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI4/MM5 N_XI0/XI20/XI4/NET34_XI0/XI20/XI4/MM5_d
+ N_XI0/XI20/XI4/NET33_XI0/XI20/XI4/MM5_g N_VDD_XI0/XI20/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI4/MM4 N_XI0/XI20/XI4/NET33_XI0/XI20/XI4/MM4_d
+ N_XI0/XI20/XI4/NET34_XI0/XI20/XI4/MM4_g N_VDD_XI0/XI20/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI4/MM10 N_XI0/XI20/XI4/NET35_XI0/XI20/XI4/MM10_d
+ N_XI0/XI20/XI4/NET36_XI0/XI20/XI4/MM10_g N_VDD_XI0/XI20/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI4/MM11 N_XI0/XI20/XI4/NET36_XI0/XI20/XI4/MM11_d
+ N_XI0/XI20/XI4/NET35_XI0/XI20/XI4/MM11_g N_VDD_XI0/XI20/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI5/MM2 N_XI0/XI20/XI5/NET34_XI0/XI20/XI5/MM2_d
+ N_XI0/XI20/XI5/NET33_XI0/XI20/XI5/MM2_g N_VSS_XI0/XI20/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM3 N_XI0/XI20/XI5/NET33_XI0/XI20/XI5/MM3_d
+ N_WL<36>_XI0/XI20/XI5/MM3_g N_BLN<10>_XI0/XI20/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM0 N_XI0/XI20/XI5/NET34_XI0/XI20/XI5/MM0_d
+ N_WL<36>_XI0/XI20/XI5/MM0_g N_BL<10>_XI0/XI20/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM1 N_XI0/XI20/XI5/NET33_XI0/XI20/XI5/MM1_d
+ N_XI0/XI20/XI5/NET34_XI0/XI20/XI5/MM1_g N_VSS_XI0/XI20/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM9 N_XI0/XI20/XI5/NET36_XI0/XI20/XI5/MM9_d
+ N_WL<37>_XI0/XI20/XI5/MM9_g N_BL<10>_XI0/XI20/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM6 N_XI0/XI20/XI5/NET35_XI0/XI20/XI5/MM6_d
+ N_XI0/XI20/XI5/NET36_XI0/XI20/XI5/MM6_g N_VSS_XI0/XI20/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM7 N_XI0/XI20/XI5/NET36_XI0/XI20/XI5/MM7_d
+ N_XI0/XI20/XI5/NET35_XI0/XI20/XI5/MM7_g N_VSS_XI0/XI20/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM8 N_XI0/XI20/XI5/NET35_XI0/XI20/XI5/MM8_d
+ N_WL<37>_XI0/XI20/XI5/MM8_g N_BLN<10>_XI0/XI20/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI5/MM5 N_XI0/XI20/XI5/NET34_XI0/XI20/XI5/MM5_d
+ N_XI0/XI20/XI5/NET33_XI0/XI20/XI5/MM5_g N_VDD_XI0/XI20/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI5/MM4 N_XI0/XI20/XI5/NET33_XI0/XI20/XI5/MM4_d
+ N_XI0/XI20/XI5/NET34_XI0/XI20/XI5/MM4_g N_VDD_XI0/XI20/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI5/MM10 N_XI0/XI20/XI5/NET35_XI0/XI20/XI5/MM10_d
+ N_XI0/XI20/XI5/NET36_XI0/XI20/XI5/MM10_g N_VDD_XI0/XI20/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI5/MM11 N_XI0/XI20/XI5/NET36_XI0/XI20/XI5/MM11_d
+ N_XI0/XI20/XI5/NET35_XI0/XI20/XI5/MM11_g N_VDD_XI0/XI20/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI6/MM2 N_XI0/XI20/XI6/NET34_XI0/XI20/XI6/MM2_d
+ N_XI0/XI20/XI6/NET33_XI0/XI20/XI6/MM2_g N_VSS_XI0/XI20/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM3 N_XI0/XI20/XI6/NET33_XI0/XI20/XI6/MM3_d
+ N_WL<36>_XI0/XI20/XI6/MM3_g N_BLN<9>_XI0/XI20/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM0 N_XI0/XI20/XI6/NET34_XI0/XI20/XI6/MM0_d
+ N_WL<36>_XI0/XI20/XI6/MM0_g N_BL<9>_XI0/XI20/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM1 N_XI0/XI20/XI6/NET33_XI0/XI20/XI6/MM1_d
+ N_XI0/XI20/XI6/NET34_XI0/XI20/XI6/MM1_g N_VSS_XI0/XI20/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM9 N_XI0/XI20/XI6/NET36_XI0/XI20/XI6/MM9_d
+ N_WL<37>_XI0/XI20/XI6/MM9_g N_BL<9>_XI0/XI20/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM6 N_XI0/XI20/XI6/NET35_XI0/XI20/XI6/MM6_d
+ N_XI0/XI20/XI6/NET36_XI0/XI20/XI6/MM6_g N_VSS_XI0/XI20/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM7 N_XI0/XI20/XI6/NET36_XI0/XI20/XI6/MM7_d
+ N_XI0/XI20/XI6/NET35_XI0/XI20/XI6/MM7_g N_VSS_XI0/XI20/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM8 N_XI0/XI20/XI6/NET35_XI0/XI20/XI6/MM8_d
+ N_WL<37>_XI0/XI20/XI6/MM8_g N_BLN<9>_XI0/XI20/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI6/MM5 N_XI0/XI20/XI6/NET34_XI0/XI20/XI6/MM5_d
+ N_XI0/XI20/XI6/NET33_XI0/XI20/XI6/MM5_g N_VDD_XI0/XI20/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI6/MM4 N_XI0/XI20/XI6/NET33_XI0/XI20/XI6/MM4_d
+ N_XI0/XI20/XI6/NET34_XI0/XI20/XI6/MM4_g N_VDD_XI0/XI20/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI6/MM10 N_XI0/XI20/XI6/NET35_XI0/XI20/XI6/MM10_d
+ N_XI0/XI20/XI6/NET36_XI0/XI20/XI6/MM10_g N_VDD_XI0/XI20/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI6/MM11 N_XI0/XI20/XI6/NET36_XI0/XI20/XI6/MM11_d
+ N_XI0/XI20/XI6/NET35_XI0/XI20/XI6/MM11_g N_VDD_XI0/XI20/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI7/MM2 N_XI0/XI20/XI7/NET34_XI0/XI20/XI7/MM2_d
+ N_XI0/XI20/XI7/NET33_XI0/XI20/XI7/MM2_g N_VSS_XI0/XI20/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM3 N_XI0/XI20/XI7/NET33_XI0/XI20/XI7/MM3_d
+ N_WL<36>_XI0/XI20/XI7/MM3_g N_BLN<8>_XI0/XI20/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM0 N_XI0/XI20/XI7/NET34_XI0/XI20/XI7/MM0_d
+ N_WL<36>_XI0/XI20/XI7/MM0_g N_BL<8>_XI0/XI20/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM1 N_XI0/XI20/XI7/NET33_XI0/XI20/XI7/MM1_d
+ N_XI0/XI20/XI7/NET34_XI0/XI20/XI7/MM1_g N_VSS_XI0/XI20/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM9 N_XI0/XI20/XI7/NET36_XI0/XI20/XI7/MM9_d
+ N_WL<37>_XI0/XI20/XI7/MM9_g N_BL<8>_XI0/XI20/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM6 N_XI0/XI20/XI7/NET35_XI0/XI20/XI7/MM6_d
+ N_XI0/XI20/XI7/NET36_XI0/XI20/XI7/MM6_g N_VSS_XI0/XI20/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM7 N_XI0/XI20/XI7/NET36_XI0/XI20/XI7/MM7_d
+ N_XI0/XI20/XI7/NET35_XI0/XI20/XI7/MM7_g N_VSS_XI0/XI20/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM8 N_XI0/XI20/XI7/NET35_XI0/XI20/XI7/MM8_d
+ N_WL<37>_XI0/XI20/XI7/MM8_g N_BLN<8>_XI0/XI20/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI7/MM5 N_XI0/XI20/XI7/NET34_XI0/XI20/XI7/MM5_d
+ N_XI0/XI20/XI7/NET33_XI0/XI20/XI7/MM5_g N_VDD_XI0/XI20/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI7/MM4 N_XI0/XI20/XI7/NET33_XI0/XI20/XI7/MM4_d
+ N_XI0/XI20/XI7/NET34_XI0/XI20/XI7/MM4_g N_VDD_XI0/XI20/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI7/MM10 N_XI0/XI20/XI7/NET35_XI0/XI20/XI7/MM10_d
+ N_XI0/XI20/XI7/NET36_XI0/XI20/XI7/MM10_g N_VDD_XI0/XI20/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI7/MM11 N_XI0/XI20/XI7/NET36_XI0/XI20/XI7/MM11_d
+ N_XI0/XI20/XI7/NET35_XI0/XI20/XI7/MM11_g N_VDD_XI0/XI20/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI8/MM2 N_XI0/XI20/XI8/NET34_XI0/XI20/XI8/MM2_d
+ N_XI0/XI20/XI8/NET33_XI0/XI20/XI8/MM2_g N_VSS_XI0/XI20/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM3 N_XI0/XI20/XI8/NET33_XI0/XI20/XI8/MM3_d
+ N_WL<36>_XI0/XI20/XI8/MM3_g N_BLN<7>_XI0/XI20/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM0 N_XI0/XI20/XI8/NET34_XI0/XI20/XI8/MM0_d
+ N_WL<36>_XI0/XI20/XI8/MM0_g N_BL<7>_XI0/XI20/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM1 N_XI0/XI20/XI8/NET33_XI0/XI20/XI8/MM1_d
+ N_XI0/XI20/XI8/NET34_XI0/XI20/XI8/MM1_g N_VSS_XI0/XI20/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM9 N_XI0/XI20/XI8/NET36_XI0/XI20/XI8/MM9_d
+ N_WL<37>_XI0/XI20/XI8/MM9_g N_BL<7>_XI0/XI20/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM6 N_XI0/XI20/XI8/NET35_XI0/XI20/XI8/MM6_d
+ N_XI0/XI20/XI8/NET36_XI0/XI20/XI8/MM6_g N_VSS_XI0/XI20/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM7 N_XI0/XI20/XI8/NET36_XI0/XI20/XI8/MM7_d
+ N_XI0/XI20/XI8/NET35_XI0/XI20/XI8/MM7_g N_VSS_XI0/XI20/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM8 N_XI0/XI20/XI8/NET35_XI0/XI20/XI8/MM8_d
+ N_WL<37>_XI0/XI20/XI8/MM8_g N_BLN<7>_XI0/XI20/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI8/MM5 N_XI0/XI20/XI8/NET34_XI0/XI20/XI8/MM5_d
+ N_XI0/XI20/XI8/NET33_XI0/XI20/XI8/MM5_g N_VDD_XI0/XI20/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI8/MM4 N_XI0/XI20/XI8/NET33_XI0/XI20/XI8/MM4_d
+ N_XI0/XI20/XI8/NET34_XI0/XI20/XI8/MM4_g N_VDD_XI0/XI20/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI8/MM10 N_XI0/XI20/XI8/NET35_XI0/XI20/XI8/MM10_d
+ N_XI0/XI20/XI8/NET36_XI0/XI20/XI8/MM10_g N_VDD_XI0/XI20/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI8/MM11 N_XI0/XI20/XI8/NET36_XI0/XI20/XI8/MM11_d
+ N_XI0/XI20/XI8/NET35_XI0/XI20/XI8/MM11_g N_VDD_XI0/XI20/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI9/MM2 N_XI0/XI20/XI9/NET34_XI0/XI20/XI9/MM2_d
+ N_XI0/XI20/XI9/NET33_XI0/XI20/XI9/MM2_g N_VSS_XI0/XI20/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM3 N_XI0/XI20/XI9/NET33_XI0/XI20/XI9/MM3_d
+ N_WL<36>_XI0/XI20/XI9/MM3_g N_BLN<6>_XI0/XI20/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM0 N_XI0/XI20/XI9/NET34_XI0/XI20/XI9/MM0_d
+ N_WL<36>_XI0/XI20/XI9/MM0_g N_BL<6>_XI0/XI20/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM1 N_XI0/XI20/XI9/NET33_XI0/XI20/XI9/MM1_d
+ N_XI0/XI20/XI9/NET34_XI0/XI20/XI9/MM1_g N_VSS_XI0/XI20/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM9 N_XI0/XI20/XI9/NET36_XI0/XI20/XI9/MM9_d
+ N_WL<37>_XI0/XI20/XI9/MM9_g N_BL<6>_XI0/XI20/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM6 N_XI0/XI20/XI9/NET35_XI0/XI20/XI9/MM6_d
+ N_XI0/XI20/XI9/NET36_XI0/XI20/XI9/MM6_g N_VSS_XI0/XI20/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM7 N_XI0/XI20/XI9/NET36_XI0/XI20/XI9/MM7_d
+ N_XI0/XI20/XI9/NET35_XI0/XI20/XI9/MM7_g N_VSS_XI0/XI20/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM8 N_XI0/XI20/XI9/NET35_XI0/XI20/XI9/MM8_d
+ N_WL<37>_XI0/XI20/XI9/MM8_g N_BLN<6>_XI0/XI20/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI9/MM5 N_XI0/XI20/XI9/NET34_XI0/XI20/XI9/MM5_d
+ N_XI0/XI20/XI9/NET33_XI0/XI20/XI9/MM5_g N_VDD_XI0/XI20/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI9/MM4 N_XI0/XI20/XI9/NET33_XI0/XI20/XI9/MM4_d
+ N_XI0/XI20/XI9/NET34_XI0/XI20/XI9/MM4_g N_VDD_XI0/XI20/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI9/MM10 N_XI0/XI20/XI9/NET35_XI0/XI20/XI9/MM10_d
+ N_XI0/XI20/XI9/NET36_XI0/XI20/XI9/MM10_g N_VDD_XI0/XI20/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI9/MM11 N_XI0/XI20/XI9/NET36_XI0/XI20/XI9/MM11_d
+ N_XI0/XI20/XI9/NET35_XI0/XI20/XI9/MM11_g N_VDD_XI0/XI20/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI10/MM2 N_XI0/XI20/XI10/NET34_XI0/XI20/XI10/MM2_d
+ N_XI0/XI20/XI10/NET33_XI0/XI20/XI10/MM2_g N_VSS_XI0/XI20/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM3 N_XI0/XI20/XI10/NET33_XI0/XI20/XI10/MM3_d
+ N_WL<36>_XI0/XI20/XI10/MM3_g N_BLN<5>_XI0/XI20/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM0 N_XI0/XI20/XI10/NET34_XI0/XI20/XI10/MM0_d
+ N_WL<36>_XI0/XI20/XI10/MM0_g N_BL<5>_XI0/XI20/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM1 N_XI0/XI20/XI10/NET33_XI0/XI20/XI10/MM1_d
+ N_XI0/XI20/XI10/NET34_XI0/XI20/XI10/MM1_g N_VSS_XI0/XI20/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM9 N_XI0/XI20/XI10/NET36_XI0/XI20/XI10/MM9_d
+ N_WL<37>_XI0/XI20/XI10/MM9_g N_BL<5>_XI0/XI20/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM6 N_XI0/XI20/XI10/NET35_XI0/XI20/XI10/MM6_d
+ N_XI0/XI20/XI10/NET36_XI0/XI20/XI10/MM6_g N_VSS_XI0/XI20/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM7 N_XI0/XI20/XI10/NET36_XI0/XI20/XI10/MM7_d
+ N_XI0/XI20/XI10/NET35_XI0/XI20/XI10/MM7_g N_VSS_XI0/XI20/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM8 N_XI0/XI20/XI10/NET35_XI0/XI20/XI10/MM8_d
+ N_WL<37>_XI0/XI20/XI10/MM8_g N_BLN<5>_XI0/XI20/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI10/MM5 N_XI0/XI20/XI10/NET34_XI0/XI20/XI10/MM5_d
+ N_XI0/XI20/XI10/NET33_XI0/XI20/XI10/MM5_g N_VDD_XI0/XI20/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI10/MM4 N_XI0/XI20/XI10/NET33_XI0/XI20/XI10/MM4_d
+ N_XI0/XI20/XI10/NET34_XI0/XI20/XI10/MM4_g N_VDD_XI0/XI20/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI10/MM10 N_XI0/XI20/XI10/NET35_XI0/XI20/XI10/MM10_d
+ N_XI0/XI20/XI10/NET36_XI0/XI20/XI10/MM10_g N_VDD_XI0/XI20/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI10/MM11 N_XI0/XI20/XI10/NET36_XI0/XI20/XI10/MM11_d
+ N_XI0/XI20/XI10/NET35_XI0/XI20/XI10/MM11_g N_VDD_XI0/XI20/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI11/MM2 N_XI0/XI20/XI11/NET34_XI0/XI20/XI11/MM2_d
+ N_XI0/XI20/XI11/NET33_XI0/XI20/XI11/MM2_g N_VSS_XI0/XI20/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM3 N_XI0/XI20/XI11/NET33_XI0/XI20/XI11/MM3_d
+ N_WL<36>_XI0/XI20/XI11/MM3_g N_BLN<4>_XI0/XI20/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM0 N_XI0/XI20/XI11/NET34_XI0/XI20/XI11/MM0_d
+ N_WL<36>_XI0/XI20/XI11/MM0_g N_BL<4>_XI0/XI20/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM1 N_XI0/XI20/XI11/NET33_XI0/XI20/XI11/MM1_d
+ N_XI0/XI20/XI11/NET34_XI0/XI20/XI11/MM1_g N_VSS_XI0/XI20/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM9 N_XI0/XI20/XI11/NET36_XI0/XI20/XI11/MM9_d
+ N_WL<37>_XI0/XI20/XI11/MM9_g N_BL<4>_XI0/XI20/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM6 N_XI0/XI20/XI11/NET35_XI0/XI20/XI11/MM6_d
+ N_XI0/XI20/XI11/NET36_XI0/XI20/XI11/MM6_g N_VSS_XI0/XI20/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM7 N_XI0/XI20/XI11/NET36_XI0/XI20/XI11/MM7_d
+ N_XI0/XI20/XI11/NET35_XI0/XI20/XI11/MM7_g N_VSS_XI0/XI20/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM8 N_XI0/XI20/XI11/NET35_XI0/XI20/XI11/MM8_d
+ N_WL<37>_XI0/XI20/XI11/MM8_g N_BLN<4>_XI0/XI20/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI11/MM5 N_XI0/XI20/XI11/NET34_XI0/XI20/XI11/MM5_d
+ N_XI0/XI20/XI11/NET33_XI0/XI20/XI11/MM5_g N_VDD_XI0/XI20/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI11/MM4 N_XI0/XI20/XI11/NET33_XI0/XI20/XI11/MM4_d
+ N_XI0/XI20/XI11/NET34_XI0/XI20/XI11/MM4_g N_VDD_XI0/XI20/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI11/MM10 N_XI0/XI20/XI11/NET35_XI0/XI20/XI11/MM10_d
+ N_XI0/XI20/XI11/NET36_XI0/XI20/XI11/MM10_g N_VDD_XI0/XI20/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI11/MM11 N_XI0/XI20/XI11/NET36_XI0/XI20/XI11/MM11_d
+ N_XI0/XI20/XI11/NET35_XI0/XI20/XI11/MM11_g N_VDD_XI0/XI20/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI12/MM2 N_XI0/XI20/XI12/NET34_XI0/XI20/XI12/MM2_d
+ N_XI0/XI20/XI12/NET33_XI0/XI20/XI12/MM2_g N_VSS_XI0/XI20/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM3 N_XI0/XI20/XI12/NET33_XI0/XI20/XI12/MM3_d
+ N_WL<36>_XI0/XI20/XI12/MM3_g N_BLN<3>_XI0/XI20/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM0 N_XI0/XI20/XI12/NET34_XI0/XI20/XI12/MM0_d
+ N_WL<36>_XI0/XI20/XI12/MM0_g N_BL<3>_XI0/XI20/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM1 N_XI0/XI20/XI12/NET33_XI0/XI20/XI12/MM1_d
+ N_XI0/XI20/XI12/NET34_XI0/XI20/XI12/MM1_g N_VSS_XI0/XI20/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM9 N_XI0/XI20/XI12/NET36_XI0/XI20/XI12/MM9_d
+ N_WL<37>_XI0/XI20/XI12/MM9_g N_BL<3>_XI0/XI20/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM6 N_XI0/XI20/XI12/NET35_XI0/XI20/XI12/MM6_d
+ N_XI0/XI20/XI12/NET36_XI0/XI20/XI12/MM6_g N_VSS_XI0/XI20/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM7 N_XI0/XI20/XI12/NET36_XI0/XI20/XI12/MM7_d
+ N_XI0/XI20/XI12/NET35_XI0/XI20/XI12/MM7_g N_VSS_XI0/XI20/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM8 N_XI0/XI20/XI12/NET35_XI0/XI20/XI12/MM8_d
+ N_WL<37>_XI0/XI20/XI12/MM8_g N_BLN<3>_XI0/XI20/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI12/MM5 N_XI0/XI20/XI12/NET34_XI0/XI20/XI12/MM5_d
+ N_XI0/XI20/XI12/NET33_XI0/XI20/XI12/MM5_g N_VDD_XI0/XI20/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI12/MM4 N_XI0/XI20/XI12/NET33_XI0/XI20/XI12/MM4_d
+ N_XI0/XI20/XI12/NET34_XI0/XI20/XI12/MM4_g N_VDD_XI0/XI20/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI12/MM10 N_XI0/XI20/XI12/NET35_XI0/XI20/XI12/MM10_d
+ N_XI0/XI20/XI12/NET36_XI0/XI20/XI12/MM10_g N_VDD_XI0/XI20/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI12/MM11 N_XI0/XI20/XI12/NET36_XI0/XI20/XI12/MM11_d
+ N_XI0/XI20/XI12/NET35_XI0/XI20/XI12/MM11_g N_VDD_XI0/XI20/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI13/MM2 N_XI0/XI20/XI13/NET34_XI0/XI20/XI13/MM2_d
+ N_XI0/XI20/XI13/NET33_XI0/XI20/XI13/MM2_g N_VSS_XI0/XI20/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM3 N_XI0/XI20/XI13/NET33_XI0/XI20/XI13/MM3_d
+ N_WL<36>_XI0/XI20/XI13/MM3_g N_BLN<2>_XI0/XI20/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM0 N_XI0/XI20/XI13/NET34_XI0/XI20/XI13/MM0_d
+ N_WL<36>_XI0/XI20/XI13/MM0_g N_BL<2>_XI0/XI20/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM1 N_XI0/XI20/XI13/NET33_XI0/XI20/XI13/MM1_d
+ N_XI0/XI20/XI13/NET34_XI0/XI20/XI13/MM1_g N_VSS_XI0/XI20/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM9 N_XI0/XI20/XI13/NET36_XI0/XI20/XI13/MM9_d
+ N_WL<37>_XI0/XI20/XI13/MM9_g N_BL<2>_XI0/XI20/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM6 N_XI0/XI20/XI13/NET35_XI0/XI20/XI13/MM6_d
+ N_XI0/XI20/XI13/NET36_XI0/XI20/XI13/MM6_g N_VSS_XI0/XI20/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM7 N_XI0/XI20/XI13/NET36_XI0/XI20/XI13/MM7_d
+ N_XI0/XI20/XI13/NET35_XI0/XI20/XI13/MM7_g N_VSS_XI0/XI20/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM8 N_XI0/XI20/XI13/NET35_XI0/XI20/XI13/MM8_d
+ N_WL<37>_XI0/XI20/XI13/MM8_g N_BLN<2>_XI0/XI20/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI13/MM5 N_XI0/XI20/XI13/NET34_XI0/XI20/XI13/MM5_d
+ N_XI0/XI20/XI13/NET33_XI0/XI20/XI13/MM5_g N_VDD_XI0/XI20/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI13/MM4 N_XI0/XI20/XI13/NET33_XI0/XI20/XI13/MM4_d
+ N_XI0/XI20/XI13/NET34_XI0/XI20/XI13/MM4_g N_VDD_XI0/XI20/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI13/MM10 N_XI0/XI20/XI13/NET35_XI0/XI20/XI13/MM10_d
+ N_XI0/XI20/XI13/NET36_XI0/XI20/XI13/MM10_g N_VDD_XI0/XI20/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI13/MM11 N_XI0/XI20/XI13/NET36_XI0/XI20/XI13/MM11_d
+ N_XI0/XI20/XI13/NET35_XI0/XI20/XI13/MM11_g N_VDD_XI0/XI20/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI14/MM2 N_XI0/XI20/XI14/NET34_XI0/XI20/XI14/MM2_d
+ N_XI0/XI20/XI14/NET33_XI0/XI20/XI14/MM2_g N_VSS_XI0/XI20/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM3 N_XI0/XI20/XI14/NET33_XI0/XI20/XI14/MM3_d
+ N_WL<36>_XI0/XI20/XI14/MM3_g N_BLN<1>_XI0/XI20/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM0 N_XI0/XI20/XI14/NET34_XI0/XI20/XI14/MM0_d
+ N_WL<36>_XI0/XI20/XI14/MM0_g N_BL<1>_XI0/XI20/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM1 N_XI0/XI20/XI14/NET33_XI0/XI20/XI14/MM1_d
+ N_XI0/XI20/XI14/NET34_XI0/XI20/XI14/MM1_g N_VSS_XI0/XI20/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM9 N_XI0/XI20/XI14/NET36_XI0/XI20/XI14/MM9_d
+ N_WL<37>_XI0/XI20/XI14/MM9_g N_BL<1>_XI0/XI20/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM6 N_XI0/XI20/XI14/NET35_XI0/XI20/XI14/MM6_d
+ N_XI0/XI20/XI14/NET36_XI0/XI20/XI14/MM6_g N_VSS_XI0/XI20/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM7 N_XI0/XI20/XI14/NET36_XI0/XI20/XI14/MM7_d
+ N_XI0/XI20/XI14/NET35_XI0/XI20/XI14/MM7_g N_VSS_XI0/XI20/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM8 N_XI0/XI20/XI14/NET35_XI0/XI20/XI14/MM8_d
+ N_WL<37>_XI0/XI20/XI14/MM8_g N_BLN<1>_XI0/XI20/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI14/MM5 N_XI0/XI20/XI14/NET34_XI0/XI20/XI14/MM5_d
+ N_XI0/XI20/XI14/NET33_XI0/XI20/XI14/MM5_g N_VDD_XI0/XI20/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI14/MM4 N_XI0/XI20/XI14/NET33_XI0/XI20/XI14/MM4_d
+ N_XI0/XI20/XI14/NET34_XI0/XI20/XI14/MM4_g N_VDD_XI0/XI20/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI14/MM10 N_XI0/XI20/XI14/NET35_XI0/XI20/XI14/MM10_d
+ N_XI0/XI20/XI14/NET36_XI0/XI20/XI14/MM10_g N_VDD_XI0/XI20/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI14/MM11 N_XI0/XI20/XI14/NET36_XI0/XI20/XI14/MM11_d
+ N_XI0/XI20/XI14/NET35_XI0/XI20/XI14/MM11_g N_VDD_XI0/XI20/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI15/MM2 N_XI0/XI20/XI15/NET34_XI0/XI20/XI15/MM2_d
+ N_XI0/XI20/XI15/NET33_XI0/XI20/XI15/MM2_g N_VSS_XI0/XI20/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM3 N_XI0/XI20/XI15/NET33_XI0/XI20/XI15/MM3_d
+ N_WL<36>_XI0/XI20/XI15/MM3_g N_BLN<0>_XI0/XI20/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM0 N_XI0/XI20/XI15/NET34_XI0/XI20/XI15/MM0_d
+ N_WL<36>_XI0/XI20/XI15/MM0_g N_BL<0>_XI0/XI20/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM1 N_XI0/XI20/XI15/NET33_XI0/XI20/XI15/MM1_d
+ N_XI0/XI20/XI15/NET34_XI0/XI20/XI15/MM1_g N_VSS_XI0/XI20/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM9 N_XI0/XI20/XI15/NET36_XI0/XI20/XI15/MM9_d
+ N_WL<37>_XI0/XI20/XI15/MM9_g N_BL<0>_XI0/XI20/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM6 N_XI0/XI20/XI15/NET35_XI0/XI20/XI15/MM6_d
+ N_XI0/XI20/XI15/NET36_XI0/XI20/XI15/MM6_g N_VSS_XI0/XI20/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM7 N_XI0/XI20/XI15/NET36_XI0/XI20/XI15/MM7_d
+ N_XI0/XI20/XI15/NET35_XI0/XI20/XI15/MM7_g N_VSS_XI0/XI20/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM8 N_XI0/XI20/XI15/NET35_XI0/XI20/XI15/MM8_d
+ N_WL<37>_XI0/XI20/XI15/MM8_g N_BLN<0>_XI0/XI20/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI20/XI15/MM5 N_XI0/XI20/XI15/NET34_XI0/XI20/XI15/MM5_d
+ N_XI0/XI20/XI15/NET33_XI0/XI20/XI15/MM5_g N_VDD_XI0/XI20/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI15/MM4 N_XI0/XI20/XI15/NET33_XI0/XI20/XI15/MM4_d
+ N_XI0/XI20/XI15/NET34_XI0/XI20/XI15/MM4_g N_VDD_XI0/XI20/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI15/MM10 N_XI0/XI20/XI15/NET35_XI0/XI20/XI15/MM10_d
+ N_XI0/XI20/XI15/NET36_XI0/XI20/XI15/MM10_g N_VDD_XI0/XI20/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI20/XI15/MM11 N_XI0/XI20/XI15/NET36_XI0/XI20/XI15/MM11_d
+ N_XI0/XI20/XI15/NET35_XI0/XI20/XI15/MM11_g N_VDD_XI0/XI20/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI0/MM2 N_XI0/XI21/XI0/NET34_XI0/XI21/XI0/MM2_d
+ N_XI0/XI21/XI0/NET33_XI0/XI21/XI0/MM2_g N_VSS_XI0/XI21/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM3 N_XI0/XI21/XI0/NET33_XI0/XI21/XI0/MM3_d
+ N_WL<38>_XI0/XI21/XI0/MM3_g N_BLN<15>_XI0/XI21/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM0 N_XI0/XI21/XI0/NET34_XI0/XI21/XI0/MM0_d
+ N_WL<38>_XI0/XI21/XI0/MM0_g N_BL<15>_XI0/XI21/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM1 N_XI0/XI21/XI0/NET33_XI0/XI21/XI0/MM1_d
+ N_XI0/XI21/XI0/NET34_XI0/XI21/XI0/MM1_g N_VSS_XI0/XI21/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM9 N_XI0/XI21/XI0/NET36_XI0/XI21/XI0/MM9_d
+ N_WL<39>_XI0/XI21/XI0/MM9_g N_BL<15>_XI0/XI21/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM6 N_XI0/XI21/XI0/NET35_XI0/XI21/XI0/MM6_d
+ N_XI0/XI21/XI0/NET36_XI0/XI21/XI0/MM6_g N_VSS_XI0/XI21/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM7 N_XI0/XI21/XI0/NET36_XI0/XI21/XI0/MM7_d
+ N_XI0/XI21/XI0/NET35_XI0/XI21/XI0/MM7_g N_VSS_XI0/XI21/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM8 N_XI0/XI21/XI0/NET35_XI0/XI21/XI0/MM8_d
+ N_WL<39>_XI0/XI21/XI0/MM8_g N_BLN<15>_XI0/XI21/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI0/MM5 N_XI0/XI21/XI0/NET34_XI0/XI21/XI0/MM5_d
+ N_XI0/XI21/XI0/NET33_XI0/XI21/XI0/MM5_g N_VDD_XI0/XI21/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI0/MM4 N_XI0/XI21/XI0/NET33_XI0/XI21/XI0/MM4_d
+ N_XI0/XI21/XI0/NET34_XI0/XI21/XI0/MM4_g N_VDD_XI0/XI21/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI0/MM10 N_XI0/XI21/XI0/NET35_XI0/XI21/XI0/MM10_d
+ N_XI0/XI21/XI0/NET36_XI0/XI21/XI0/MM10_g N_VDD_XI0/XI21/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI0/MM11 N_XI0/XI21/XI0/NET36_XI0/XI21/XI0/MM11_d
+ N_XI0/XI21/XI0/NET35_XI0/XI21/XI0/MM11_g N_VDD_XI0/XI21/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI1/MM2 N_XI0/XI21/XI1/NET34_XI0/XI21/XI1/MM2_d
+ N_XI0/XI21/XI1/NET33_XI0/XI21/XI1/MM2_g N_VSS_XI0/XI21/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM3 N_XI0/XI21/XI1/NET33_XI0/XI21/XI1/MM3_d
+ N_WL<38>_XI0/XI21/XI1/MM3_g N_BLN<14>_XI0/XI21/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM0 N_XI0/XI21/XI1/NET34_XI0/XI21/XI1/MM0_d
+ N_WL<38>_XI0/XI21/XI1/MM0_g N_BL<14>_XI0/XI21/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM1 N_XI0/XI21/XI1/NET33_XI0/XI21/XI1/MM1_d
+ N_XI0/XI21/XI1/NET34_XI0/XI21/XI1/MM1_g N_VSS_XI0/XI21/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM9 N_XI0/XI21/XI1/NET36_XI0/XI21/XI1/MM9_d
+ N_WL<39>_XI0/XI21/XI1/MM9_g N_BL<14>_XI0/XI21/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM6 N_XI0/XI21/XI1/NET35_XI0/XI21/XI1/MM6_d
+ N_XI0/XI21/XI1/NET36_XI0/XI21/XI1/MM6_g N_VSS_XI0/XI21/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM7 N_XI0/XI21/XI1/NET36_XI0/XI21/XI1/MM7_d
+ N_XI0/XI21/XI1/NET35_XI0/XI21/XI1/MM7_g N_VSS_XI0/XI21/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM8 N_XI0/XI21/XI1/NET35_XI0/XI21/XI1/MM8_d
+ N_WL<39>_XI0/XI21/XI1/MM8_g N_BLN<14>_XI0/XI21/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI1/MM5 N_XI0/XI21/XI1/NET34_XI0/XI21/XI1/MM5_d
+ N_XI0/XI21/XI1/NET33_XI0/XI21/XI1/MM5_g N_VDD_XI0/XI21/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI1/MM4 N_XI0/XI21/XI1/NET33_XI0/XI21/XI1/MM4_d
+ N_XI0/XI21/XI1/NET34_XI0/XI21/XI1/MM4_g N_VDD_XI0/XI21/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI1/MM10 N_XI0/XI21/XI1/NET35_XI0/XI21/XI1/MM10_d
+ N_XI0/XI21/XI1/NET36_XI0/XI21/XI1/MM10_g N_VDD_XI0/XI21/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI1/MM11 N_XI0/XI21/XI1/NET36_XI0/XI21/XI1/MM11_d
+ N_XI0/XI21/XI1/NET35_XI0/XI21/XI1/MM11_g N_VDD_XI0/XI21/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI2/MM2 N_XI0/XI21/XI2/NET34_XI0/XI21/XI2/MM2_d
+ N_XI0/XI21/XI2/NET33_XI0/XI21/XI2/MM2_g N_VSS_XI0/XI21/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM3 N_XI0/XI21/XI2/NET33_XI0/XI21/XI2/MM3_d
+ N_WL<38>_XI0/XI21/XI2/MM3_g N_BLN<13>_XI0/XI21/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM0 N_XI0/XI21/XI2/NET34_XI0/XI21/XI2/MM0_d
+ N_WL<38>_XI0/XI21/XI2/MM0_g N_BL<13>_XI0/XI21/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM1 N_XI0/XI21/XI2/NET33_XI0/XI21/XI2/MM1_d
+ N_XI0/XI21/XI2/NET34_XI0/XI21/XI2/MM1_g N_VSS_XI0/XI21/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM9 N_XI0/XI21/XI2/NET36_XI0/XI21/XI2/MM9_d
+ N_WL<39>_XI0/XI21/XI2/MM9_g N_BL<13>_XI0/XI21/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM6 N_XI0/XI21/XI2/NET35_XI0/XI21/XI2/MM6_d
+ N_XI0/XI21/XI2/NET36_XI0/XI21/XI2/MM6_g N_VSS_XI0/XI21/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM7 N_XI0/XI21/XI2/NET36_XI0/XI21/XI2/MM7_d
+ N_XI0/XI21/XI2/NET35_XI0/XI21/XI2/MM7_g N_VSS_XI0/XI21/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM8 N_XI0/XI21/XI2/NET35_XI0/XI21/XI2/MM8_d
+ N_WL<39>_XI0/XI21/XI2/MM8_g N_BLN<13>_XI0/XI21/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI2/MM5 N_XI0/XI21/XI2/NET34_XI0/XI21/XI2/MM5_d
+ N_XI0/XI21/XI2/NET33_XI0/XI21/XI2/MM5_g N_VDD_XI0/XI21/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI2/MM4 N_XI0/XI21/XI2/NET33_XI0/XI21/XI2/MM4_d
+ N_XI0/XI21/XI2/NET34_XI0/XI21/XI2/MM4_g N_VDD_XI0/XI21/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI2/MM10 N_XI0/XI21/XI2/NET35_XI0/XI21/XI2/MM10_d
+ N_XI0/XI21/XI2/NET36_XI0/XI21/XI2/MM10_g N_VDD_XI0/XI21/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI2/MM11 N_XI0/XI21/XI2/NET36_XI0/XI21/XI2/MM11_d
+ N_XI0/XI21/XI2/NET35_XI0/XI21/XI2/MM11_g N_VDD_XI0/XI21/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI3/MM2 N_XI0/XI21/XI3/NET34_XI0/XI21/XI3/MM2_d
+ N_XI0/XI21/XI3/NET33_XI0/XI21/XI3/MM2_g N_VSS_XI0/XI21/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM3 N_XI0/XI21/XI3/NET33_XI0/XI21/XI3/MM3_d
+ N_WL<38>_XI0/XI21/XI3/MM3_g N_BLN<12>_XI0/XI21/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM0 N_XI0/XI21/XI3/NET34_XI0/XI21/XI3/MM0_d
+ N_WL<38>_XI0/XI21/XI3/MM0_g N_BL<12>_XI0/XI21/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM1 N_XI0/XI21/XI3/NET33_XI0/XI21/XI3/MM1_d
+ N_XI0/XI21/XI3/NET34_XI0/XI21/XI3/MM1_g N_VSS_XI0/XI21/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM9 N_XI0/XI21/XI3/NET36_XI0/XI21/XI3/MM9_d
+ N_WL<39>_XI0/XI21/XI3/MM9_g N_BL<12>_XI0/XI21/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM6 N_XI0/XI21/XI3/NET35_XI0/XI21/XI3/MM6_d
+ N_XI0/XI21/XI3/NET36_XI0/XI21/XI3/MM6_g N_VSS_XI0/XI21/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM7 N_XI0/XI21/XI3/NET36_XI0/XI21/XI3/MM7_d
+ N_XI0/XI21/XI3/NET35_XI0/XI21/XI3/MM7_g N_VSS_XI0/XI21/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM8 N_XI0/XI21/XI3/NET35_XI0/XI21/XI3/MM8_d
+ N_WL<39>_XI0/XI21/XI3/MM8_g N_BLN<12>_XI0/XI21/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI3/MM5 N_XI0/XI21/XI3/NET34_XI0/XI21/XI3/MM5_d
+ N_XI0/XI21/XI3/NET33_XI0/XI21/XI3/MM5_g N_VDD_XI0/XI21/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI3/MM4 N_XI0/XI21/XI3/NET33_XI0/XI21/XI3/MM4_d
+ N_XI0/XI21/XI3/NET34_XI0/XI21/XI3/MM4_g N_VDD_XI0/XI21/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI3/MM10 N_XI0/XI21/XI3/NET35_XI0/XI21/XI3/MM10_d
+ N_XI0/XI21/XI3/NET36_XI0/XI21/XI3/MM10_g N_VDD_XI0/XI21/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI3/MM11 N_XI0/XI21/XI3/NET36_XI0/XI21/XI3/MM11_d
+ N_XI0/XI21/XI3/NET35_XI0/XI21/XI3/MM11_g N_VDD_XI0/XI21/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI4/MM2 N_XI0/XI21/XI4/NET34_XI0/XI21/XI4/MM2_d
+ N_XI0/XI21/XI4/NET33_XI0/XI21/XI4/MM2_g N_VSS_XI0/XI21/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM3 N_XI0/XI21/XI4/NET33_XI0/XI21/XI4/MM3_d
+ N_WL<38>_XI0/XI21/XI4/MM3_g N_BLN<11>_XI0/XI21/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM0 N_XI0/XI21/XI4/NET34_XI0/XI21/XI4/MM0_d
+ N_WL<38>_XI0/XI21/XI4/MM0_g N_BL<11>_XI0/XI21/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM1 N_XI0/XI21/XI4/NET33_XI0/XI21/XI4/MM1_d
+ N_XI0/XI21/XI4/NET34_XI0/XI21/XI4/MM1_g N_VSS_XI0/XI21/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM9 N_XI0/XI21/XI4/NET36_XI0/XI21/XI4/MM9_d
+ N_WL<39>_XI0/XI21/XI4/MM9_g N_BL<11>_XI0/XI21/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM6 N_XI0/XI21/XI4/NET35_XI0/XI21/XI4/MM6_d
+ N_XI0/XI21/XI4/NET36_XI0/XI21/XI4/MM6_g N_VSS_XI0/XI21/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM7 N_XI0/XI21/XI4/NET36_XI0/XI21/XI4/MM7_d
+ N_XI0/XI21/XI4/NET35_XI0/XI21/XI4/MM7_g N_VSS_XI0/XI21/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM8 N_XI0/XI21/XI4/NET35_XI0/XI21/XI4/MM8_d
+ N_WL<39>_XI0/XI21/XI4/MM8_g N_BLN<11>_XI0/XI21/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI4/MM5 N_XI0/XI21/XI4/NET34_XI0/XI21/XI4/MM5_d
+ N_XI0/XI21/XI4/NET33_XI0/XI21/XI4/MM5_g N_VDD_XI0/XI21/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI4/MM4 N_XI0/XI21/XI4/NET33_XI0/XI21/XI4/MM4_d
+ N_XI0/XI21/XI4/NET34_XI0/XI21/XI4/MM4_g N_VDD_XI0/XI21/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI4/MM10 N_XI0/XI21/XI4/NET35_XI0/XI21/XI4/MM10_d
+ N_XI0/XI21/XI4/NET36_XI0/XI21/XI4/MM10_g N_VDD_XI0/XI21/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI4/MM11 N_XI0/XI21/XI4/NET36_XI0/XI21/XI4/MM11_d
+ N_XI0/XI21/XI4/NET35_XI0/XI21/XI4/MM11_g N_VDD_XI0/XI21/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI5/MM2 N_XI0/XI21/XI5/NET34_XI0/XI21/XI5/MM2_d
+ N_XI0/XI21/XI5/NET33_XI0/XI21/XI5/MM2_g N_VSS_XI0/XI21/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM3 N_XI0/XI21/XI5/NET33_XI0/XI21/XI5/MM3_d
+ N_WL<38>_XI0/XI21/XI5/MM3_g N_BLN<10>_XI0/XI21/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM0 N_XI0/XI21/XI5/NET34_XI0/XI21/XI5/MM0_d
+ N_WL<38>_XI0/XI21/XI5/MM0_g N_BL<10>_XI0/XI21/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM1 N_XI0/XI21/XI5/NET33_XI0/XI21/XI5/MM1_d
+ N_XI0/XI21/XI5/NET34_XI0/XI21/XI5/MM1_g N_VSS_XI0/XI21/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM9 N_XI0/XI21/XI5/NET36_XI0/XI21/XI5/MM9_d
+ N_WL<39>_XI0/XI21/XI5/MM9_g N_BL<10>_XI0/XI21/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM6 N_XI0/XI21/XI5/NET35_XI0/XI21/XI5/MM6_d
+ N_XI0/XI21/XI5/NET36_XI0/XI21/XI5/MM6_g N_VSS_XI0/XI21/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM7 N_XI0/XI21/XI5/NET36_XI0/XI21/XI5/MM7_d
+ N_XI0/XI21/XI5/NET35_XI0/XI21/XI5/MM7_g N_VSS_XI0/XI21/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM8 N_XI0/XI21/XI5/NET35_XI0/XI21/XI5/MM8_d
+ N_WL<39>_XI0/XI21/XI5/MM8_g N_BLN<10>_XI0/XI21/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI5/MM5 N_XI0/XI21/XI5/NET34_XI0/XI21/XI5/MM5_d
+ N_XI0/XI21/XI5/NET33_XI0/XI21/XI5/MM5_g N_VDD_XI0/XI21/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI5/MM4 N_XI0/XI21/XI5/NET33_XI0/XI21/XI5/MM4_d
+ N_XI0/XI21/XI5/NET34_XI0/XI21/XI5/MM4_g N_VDD_XI0/XI21/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI5/MM10 N_XI0/XI21/XI5/NET35_XI0/XI21/XI5/MM10_d
+ N_XI0/XI21/XI5/NET36_XI0/XI21/XI5/MM10_g N_VDD_XI0/XI21/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI5/MM11 N_XI0/XI21/XI5/NET36_XI0/XI21/XI5/MM11_d
+ N_XI0/XI21/XI5/NET35_XI0/XI21/XI5/MM11_g N_VDD_XI0/XI21/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI6/MM2 N_XI0/XI21/XI6/NET34_XI0/XI21/XI6/MM2_d
+ N_XI0/XI21/XI6/NET33_XI0/XI21/XI6/MM2_g N_VSS_XI0/XI21/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM3 N_XI0/XI21/XI6/NET33_XI0/XI21/XI6/MM3_d
+ N_WL<38>_XI0/XI21/XI6/MM3_g N_BLN<9>_XI0/XI21/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM0 N_XI0/XI21/XI6/NET34_XI0/XI21/XI6/MM0_d
+ N_WL<38>_XI0/XI21/XI6/MM0_g N_BL<9>_XI0/XI21/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM1 N_XI0/XI21/XI6/NET33_XI0/XI21/XI6/MM1_d
+ N_XI0/XI21/XI6/NET34_XI0/XI21/XI6/MM1_g N_VSS_XI0/XI21/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM9 N_XI0/XI21/XI6/NET36_XI0/XI21/XI6/MM9_d
+ N_WL<39>_XI0/XI21/XI6/MM9_g N_BL<9>_XI0/XI21/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM6 N_XI0/XI21/XI6/NET35_XI0/XI21/XI6/MM6_d
+ N_XI0/XI21/XI6/NET36_XI0/XI21/XI6/MM6_g N_VSS_XI0/XI21/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM7 N_XI0/XI21/XI6/NET36_XI0/XI21/XI6/MM7_d
+ N_XI0/XI21/XI6/NET35_XI0/XI21/XI6/MM7_g N_VSS_XI0/XI21/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM8 N_XI0/XI21/XI6/NET35_XI0/XI21/XI6/MM8_d
+ N_WL<39>_XI0/XI21/XI6/MM8_g N_BLN<9>_XI0/XI21/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI6/MM5 N_XI0/XI21/XI6/NET34_XI0/XI21/XI6/MM5_d
+ N_XI0/XI21/XI6/NET33_XI0/XI21/XI6/MM5_g N_VDD_XI0/XI21/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI6/MM4 N_XI0/XI21/XI6/NET33_XI0/XI21/XI6/MM4_d
+ N_XI0/XI21/XI6/NET34_XI0/XI21/XI6/MM4_g N_VDD_XI0/XI21/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI6/MM10 N_XI0/XI21/XI6/NET35_XI0/XI21/XI6/MM10_d
+ N_XI0/XI21/XI6/NET36_XI0/XI21/XI6/MM10_g N_VDD_XI0/XI21/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI6/MM11 N_XI0/XI21/XI6/NET36_XI0/XI21/XI6/MM11_d
+ N_XI0/XI21/XI6/NET35_XI0/XI21/XI6/MM11_g N_VDD_XI0/XI21/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI7/MM2 N_XI0/XI21/XI7/NET34_XI0/XI21/XI7/MM2_d
+ N_XI0/XI21/XI7/NET33_XI0/XI21/XI7/MM2_g N_VSS_XI0/XI21/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM3 N_XI0/XI21/XI7/NET33_XI0/XI21/XI7/MM3_d
+ N_WL<38>_XI0/XI21/XI7/MM3_g N_BLN<8>_XI0/XI21/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM0 N_XI0/XI21/XI7/NET34_XI0/XI21/XI7/MM0_d
+ N_WL<38>_XI0/XI21/XI7/MM0_g N_BL<8>_XI0/XI21/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM1 N_XI0/XI21/XI7/NET33_XI0/XI21/XI7/MM1_d
+ N_XI0/XI21/XI7/NET34_XI0/XI21/XI7/MM1_g N_VSS_XI0/XI21/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM9 N_XI0/XI21/XI7/NET36_XI0/XI21/XI7/MM9_d
+ N_WL<39>_XI0/XI21/XI7/MM9_g N_BL<8>_XI0/XI21/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM6 N_XI0/XI21/XI7/NET35_XI0/XI21/XI7/MM6_d
+ N_XI0/XI21/XI7/NET36_XI0/XI21/XI7/MM6_g N_VSS_XI0/XI21/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM7 N_XI0/XI21/XI7/NET36_XI0/XI21/XI7/MM7_d
+ N_XI0/XI21/XI7/NET35_XI0/XI21/XI7/MM7_g N_VSS_XI0/XI21/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM8 N_XI0/XI21/XI7/NET35_XI0/XI21/XI7/MM8_d
+ N_WL<39>_XI0/XI21/XI7/MM8_g N_BLN<8>_XI0/XI21/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI7/MM5 N_XI0/XI21/XI7/NET34_XI0/XI21/XI7/MM5_d
+ N_XI0/XI21/XI7/NET33_XI0/XI21/XI7/MM5_g N_VDD_XI0/XI21/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI7/MM4 N_XI0/XI21/XI7/NET33_XI0/XI21/XI7/MM4_d
+ N_XI0/XI21/XI7/NET34_XI0/XI21/XI7/MM4_g N_VDD_XI0/XI21/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI7/MM10 N_XI0/XI21/XI7/NET35_XI0/XI21/XI7/MM10_d
+ N_XI0/XI21/XI7/NET36_XI0/XI21/XI7/MM10_g N_VDD_XI0/XI21/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI7/MM11 N_XI0/XI21/XI7/NET36_XI0/XI21/XI7/MM11_d
+ N_XI0/XI21/XI7/NET35_XI0/XI21/XI7/MM11_g N_VDD_XI0/XI21/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI8/MM2 N_XI0/XI21/XI8/NET34_XI0/XI21/XI8/MM2_d
+ N_XI0/XI21/XI8/NET33_XI0/XI21/XI8/MM2_g N_VSS_XI0/XI21/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM3 N_XI0/XI21/XI8/NET33_XI0/XI21/XI8/MM3_d
+ N_WL<38>_XI0/XI21/XI8/MM3_g N_BLN<7>_XI0/XI21/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM0 N_XI0/XI21/XI8/NET34_XI0/XI21/XI8/MM0_d
+ N_WL<38>_XI0/XI21/XI8/MM0_g N_BL<7>_XI0/XI21/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM1 N_XI0/XI21/XI8/NET33_XI0/XI21/XI8/MM1_d
+ N_XI0/XI21/XI8/NET34_XI0/XI21/XI8/MM1_g N_VSS_XI0/XI21/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM9 N_XI0/XI21/XI8/NET36_XI0/XI21/XI8/MM9_d
+ N_WL<39>_XI0/XI21/XI8/MM9_g N_BL<7>_XI0/XI21/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM6 N_XI0/XI21/XI8/NET35_XI0/XI21/XI8/MM6_d
+ N_XI0/XI21/XI8/NET36_XI0/XI21/XI8/MM6_g N_VSS_XI0/XI21/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM7 N_XI0/XI21/XI8/NET36_XI0/XI21/XI8/MM7_d
+ N_XI0/XI21/XI8/NET35_XI0/XI21/XI8/MM7_g N_VSS_XI0/XI21/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM8 N_XI0/XI21/XI8/NET35_XI0/XI21/XI8/MM8_d
+ N_WL<39>_XI0/XI21/XI8/MM8_g N_BLN<7>_XI0/XI21/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI8/MM5 N_XI0/XI21/XI8/NET34_XI0/XI21/XI8/MM5_d
+ N_XI0/XI21/XI8/NET33_XI0/XI21/XI8/MM5_g N_VDD_XI0/XI21/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI8/MM4 N_XI0/XI21/XI8/NET33_XI0/XI21/XI8/MM4_d
+ N_XI0/XI21/XI8/NET34_XI0/XI21/XI8/MM4_g N_VDD_XI0/XI21/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI8/MM10 N_XI0/XI21/XI8/NET35_XI0/XI21/XI8/MM10_d
+ N_XI0/XI21/XI8/NET36_XI0/XI21/XI8/MM10_g N_VDD_XI0/XI21/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI8/MM11 N_XI0/XI21/XI8/NET36_XI0/XI21/XI8/MM11_d
+ N_XI0/XI21/XI8/NET35_XI0/XI21/XI8/MM11_g N_VDD_XI0/XI21/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI9/MM2 N_XI0/XI21/XI9/NET34_XI0/XI21/XI9/MM2_d
+ N_XI0/XI21/XI9/NET33_XI0/XI21/XI9/MM2_g N_VSS_XI0/XI21/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM3 N_XI0/XI21/XI9/NET33_XI0/XI21/XI9/MM3_d
+ N_WL<38>_XI0/XI21/XI9/MM3_g N_BLN<6>_XI0/XI21/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM0 N_XI0/XI21/XI9/NET34_XI0/XI21/XI9/MM0_d
+ N_WL<38>_XI0/XI21/XI9/MM0_g N_BL<6>_XI0/XI21/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM1 N_XI0/XI21/XI9/NET33_XI0/XI21/XI9/MM1_d
+ N_XI0/XI21/XI9/NET34_XI0/XI21/XI9/MM1_g N_VSS_XI0/XI21/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM9 N_XI0/XI21/XI9/NET36_XI0/XI21/XI9/MM9_d
+ N_WL<39>_XI0/XI21/XI9/MM9_g N_BL<6>_XI0/XI21/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM6 N_XI0/XI21/XI9/NET35_XI0/XI21/XI9/MM6_d
+ N_XI0/XI21/XI9/NET36_XI0/XI21/XI9/MM6_g N_VSS_XI0/XI21/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM7 N_XI0/XI21/XI9/NET36_XI0/XI21/XI9/MM7_d
+ N_XI0/XI21/XI9/NET35_XI0/XI21/XI9/MM7_g N_VSS_XI0/XI21/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM8 N_XI0/XI21/XI9/NET35_XI0/XI21/XI9/MM8_d
+ N_WL<39>_XI0/XI21/XI9/MM8_g N_BLN<6>_XI0/XI21/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI9/MM5 N_XI0/XI21/XI9/NET34_XI0/XI21/XI9/MM5_d
+ N_XI0/XI21/XI9/NET33_XI0/XI21/XI9/MM5_g N_VDD_XI0/XI21/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI9/MM4 N_XI0/XI21/XI9/NET33_XI0/XI21/XI9/MM4_d
+ N_XI0/XI21/XI9/NET34_XI0/XI21/XI9/MM4_g N_VDD_XI0/XI21/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI9/MM10 N_XI0/XI21/XI9/NET35_XI0/XI21/XI9/MM10_d
+ N_XI0/XI21/XI9/NET36_XI0/XI21/XI9/MM10_g N_VDD_XI0/XI21/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI9/MM11 N_XI0/XI21/XI9/NET36_XI0/XI21/XI9/MM11_d
+ N_XI0/XI21/XI9/NET35_XI0/XI21/XI9/MM11_g N_VDD_XI0/XI21/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI10/MM2 N_XI0/XI21/XI10/NET34_XI0/XI21/XI10/MM2_d
+ N_XI0/XI21/XI10/NET33_XI0/XI21/XI10/MM2_g N_VSS_XI0/XI21/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM3 N_XI0/XI21/XI10/NET33_XI0/XI21/XI10/MM3_d
+ N_WL<38>_XI0/XI21/XI10/MM3_g N_BLN<5>_XI0/XI21/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM0 N_XI0/XI21/XI10/NET34_XI0/XI21/XI10/MM0_d
+ N_WL<38>_XI0/XI21/XI10/MM0_g N_BL<5>_XI0/XI21/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM1 N_XI0/XI21/XI10/NET33_XI0/XI21/XI10/MM1_d
+ N_XI0/XI21/XI10/NET34_XI0/XI21/XI10/MM1_g N_VSS_XI0/XI21/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM9 N_XI0/XI21/XI10/NET36_XI0/XI21/XI10/MM9_d
+ N_WL<39>_XI0/XI21/XI10/MM9_g N_BL<5>_XI0/XI21/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM6 N_XI0/XI21/XI10/NET35_XI0/XI21/XI10/MM6_d
+ N_XI0/XI21/XI10/NET36_XI0/XI21/XI10/MM6_g N_VSS_XI0/XI21/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM7 N_XI0/XI21/XI10/NET36_XI0/XI21/XI10/MM7_d
+ N_XI0/XI21/XI10/NET35_XI0/XI21/XI10/MM7_g N_VSS_XI0/XI21/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM8 N_XI0/XI21/XI10/NET35_XI0/XI21/XI10/MM8_d
+ N_WL<39>_XI0/XI21/XI10/MM8_g N_BLN<5>_XI0/XI21/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI10/MM5 N_XI0/XI21/XI10/NET34_XI0/XI21/XI10/MM5_d
+ N_XI0/XI21/XI10/NET33_XI0/XI21/XI10/MM5_g N_VDD_XI0/XI21/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI10/MM4 N_XI0/XI21/XI10/NET33_XI0/XI21/XI10/MM4_d
+ N_XI0/XI21/XI10/NET34_XI0/XI21/XI10/MM4_g N_VDD_XI0/XI21/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI10/MM10 N_XI0/XI21/XI10/NET35_XI0/XI21/XI10/MM10_d
+ N_XI0/XI21/XI10/NET36_XI0/XI21/XI10/MM10_g N_VDD_XI0/XI21/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI10/MM11 N_XI0/XI21/XI10/NET36_XI0/XI21/XI10/MM11_d
+ N_XI0/XI21/XI10/NET35_XI0/XI21/XI10/MM11_g N_VDD_XI0/XI21/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI11/MM2 N_XI0/XI21/XI11/NET34_XI0/XI21/XI11/MM2_d
+ N_XI0/XI21/XI11/NET33_XI0/XI21/XI11/MM2_g N_VSS_XI0/XI21/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM3 N_XI0/XI21/XI11/NET33_XI0/XI21/XI11/MM3_d
+ N_WL<38>_XI0/XI21/XI11/MM3_g N_BLN<4>_XI0/XI21/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM0 N_XI0/XI21/XI11/NET34_XI0/XI21/XI11/MM0_d
+ N_WL<38>_XI0/XI21/XI11/MM0_g N_BL<4>_XI0/XI21/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM1 N_XI0/XI21/XI11/NET33_XI0/XI21/XI11/MM1_d
+ N_XI0/XI21/XI11/NET34_XI0/XI21/XI11/MM1_g N_VSS_XI0/XI21/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM9 N_XI0/XI21/XI11/NET36_XI0/XI21/XI11/MM9_d
+ N_WL<39>_XI0/XI21/XI11/MM9_g N_BL<4>_XI0/XI21/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM6 N_XI0/XI21/XI11/NET35_XI0/XI21/XI11/MM6_d
+ N_XI0/XI21/XI11/NET36_XI0/XI21/XI11/MM6_g N_VSS_XI0/XI21/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM7 N_XI0/XI21/XI11/NET36_XI0/XI21/XI11/MM7_d
+ N_XI0/XI21/XI11/NET35_XI0/XI21/XI11/MM7_g N_VSS_XI0/XI21/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM8 N_XI0/XI21/XI11/NET35_XI0/XI21/XI11/MM8_d
+ N_WL<39>_XI0/XI21/XI11/MM8_g N_BLN<4>_XI0/XI21/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI11/MM5 N_XI0/XI21/XI11/NET34_XI0/XI21/XI11/MM5_d
+ N_XI0/XI21/XI11/NET33_XI0/XI21/XI11/MM5_g N_VDD_XI0/XI21/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI11/MM4 N_XI0/XI21/XI11/NET33_XI0/XI21/XI11/MM4_d
+ N_XI0/XI21/XI11/NET34_XI0/XI21/XI11/MM4_g N_VDD_XI0/XI21/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI11/MM10 N_XI0/XI21/XI11/NET35_XI0/XI21/XI11/MM10_d
+ N_XI0/XI21/XI11/NET36_XI0/XI21/XI11/MM10_g N_VDD_XI0/XI21/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI11/MM11 N_XI0/XI21/XI11/NET36_XI0/XI21/XI11/MM11_d
+ N_XI0/XI21/XI11/NET35_XI0/XI21/XI11/MM11_g N_VDD_XI0/XI21/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI12/MM2 N_XI0/XI21/XI12/NET34_XI0/XI21/XI12/MM2_d
+ N_XI0/XI21/XI12/NET33_XI0/XI21/XI12/MM2_g N_VSS_XI0/XI21/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM3 N_XI0/XI21/XI12/NET33_XI0/XI21/XI12/MM3_d
+ N_WL<38>_XI0/XI21/XI12/MM3_g N_BLN<3>_XI0/XI21/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM0 N_XI0/XI21/XI12/NET34_XI0/XI21/XI12/MM0_d
+ N_WL<38>_XI0/XI21/XI12/MM0_g N_BL<3>_XI0/XI21/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM1 N_XI0/XI21/XI12/NET33_XI0/XI21/XI12/MM1_d
+ N_XI0/XI21/XI12/NET34_XI0/XI21/XI12/MM1_g N_VSS_XI0/XI21/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM9 N_XI0/XI21/XI12/NET36_XI0/XI21/XI12/MM9_d
+ N_WL<39>_XI0/XI21/XI12/MM9_g N_BL<3>_XI0/XI21/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM6 N_XI0/XI21/XI12/NET35_XI0/XI21/XI12/MM6_d
+ N_XI0/XI21/XI12/NET36_XI0/XI21/XI12/MM6_g N_VSS_XI0/XI21/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM7 N_XI0/XI21/XI12/NET36_XI0/XI21/XI12/MM7_d
+ N_XI0/XI21/XI12/NET35_XI0/XI21/XI12/MM7_g N_VSS_XI0/XI21/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM8 N_XI0/XI21/XI12/NET35_XI0/XI21/XI12/MM8_d
+ N_WL<39>_XI0/XI21/XI12/MM8_g N_BLN<3>_XI0/XI21/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI12/MM5 N_XI0/XI21/XI12/NET34_XI0/XI21/XI12/MM5_d
+ N_XI0/XI21/XI12/NET33_XI0/XI21/XI12/MM5_g N_VDD_XI0/XI21/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI12/MM4 N_XI0/XI21/XI12/NET33_XI0/XI21/XI12/MM4_d
+ N_XI0/XI21/XI12/NET34_XI0/XI21/XI12/MM4_g N_VDD_XI0/XI21/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI12/MM10 N_XI0/XI21/XI12/NET35_XI0/XI21/XI12/MM10_d
+ N_XI0/XI21/XI12/NET36_XI0/XI21/XI12/MM10_g N_VDD_XI0/XI21/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI12/MM11 N_XI0/XI21/XI12/NET36_XI0/XI21/XI12/MM11_d
+ N_XI0/XI21/XI12/NET35_XI0/XI21/XI12/MM11_g N_VDD_XI0/XI21/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI13/MM2 N_XI0/XI21/XI13/NET34_XI0/XI21/XI13/MM2_d
+ N_XI0/XI21/XI13/NET33_XI0/XI21/XI13/MM2_g N_VSS_XI0/XI21/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM3 N_XI0/XI21/XI13/NET33_XI0/XI21/XI13/MM3_d
+ N_WL<38>_XI0/XI21/XI13/MM3_g N_BLN<2>_XI0/XI21/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM0 N_XI0/XI21/XI13/NET34_XI0/XI21/XI13/MM0_d
+ N_WL<38>_XI0/XI21/XI13/MM0_g N_BL<2>_XI0/XI21/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM1 N_XI0/XI21/XI13/NET33_XI0/XI21/XI13/MM1_d
+ N_XI0/XI21/XI13/NET34_XI0/XI21/XI13/MM1_g N_VSS_XI0/XI21/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM9 N_XI0/XI21/XI13/NET36_XI0/XI21/XI13/MM9_d
+ N_WL<39>_XI0/XI21/XI13/MM9_g N_BL<2>_XI0/XI21/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM6 N_XI0/XI21/XI13/NET35_XI0/XI21/XI13/MM6_d
+ N_XI0/XI21/XI13/NET36_XI0/XI21/XI13/MM6_g N_VSS_XI0/XI21/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM7 N_XI0/XI21/XI13/NET36_XI0/XI21/XI13/MM7_d
+ N_XI0/XI21/XI13/NET35_XI0/XI21/XI13/MM7_g N_VSS_XI0/XI21/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM8 N_XI0/XI21/XI13/NET35_XI0/XI21/XI13/MM8_d
+ N_WL<39>_XI0/XI21/XI13/MM8_g N_BLN<2>_XI0/XI21/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI13/MM5 N_XI0/XI21/XI13/NET34_XI0/XI21/XI13/MM5_d
+ N_XI0/XI21/XI13/NET33_XI0/XI21/XI13/MM5_g N_VDD_XI0/XI21/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI13/MM4 N_XI0/XI21/XI13/NET33_XI0/XI21/XI13/MM4_d
+ N_XI0/XI21/XI13/NET34_XI0/XI21/XI13/MM4_g N_VDD_XI0/XI21/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI13/MM10 N_XI0/XI21/XI13/NET35_XI0/XI21/XI13/MM10_d
+ N_XI0/XI21/XI13/NET36_XI0/XI21/XI13/MM10_g N_VDD_XI0/XI21/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI13/MM11 N_XI0/XI21/XI13/NET36_XI0/XI21/XI13/MM11_d
+ N_XI0/XI21/XI13/NET35_XI0/XI21/XI13/MM11_g N_VDD_XI0/XI21/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI14/MM2 N_XI0/XI21/XI14/NET34_XI0/XI21/XI14/MM2_d
+ N_XI0/XI21/XI14/NET33_XI0/XI21/XI14/MM2_g N_VSS_XI0/XI21/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM3 N_XI0/XI21/XI14/NET33_XI0/XI21/XI14/MM3_d
+ N_WL<38>_XI0/XI21/XI14/MM3_g N_BLN<1>_XI0/XI21/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM0 N_XI0/XI21/XI14/NET34_XI0/XI21/XI14/MM0_d
+ N_WL<38>_XI0/XI21/XI14/MM0_g N_BL<1>_XI0/XI21/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM1 N_XI0/XI21/XI14/NET33_XI0/XI21/XI14/MM1_d
+ N_XI0/XI21/XI14/NET34_XI0/XI21/XI14/MM1_g N_VSS_XI0/XI21/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM9 N_XI0/XI21/XI14/NET36_XI0/XI21/XI14/MM9_d
+ N_WL<39>_XI0/XI21/XI14/MM9_g N_BL<1>_XI0/XI21/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM6 N_XI0/XI21/XI14/NET35_XI0/XI21/XI14/MM6_d
+ N_XI0/XI21/XI14/NET36_XI0/XI21/XI14/MM6_g N_VSS_XI0/XI21/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM7 N_XI0/XI21/XI14/NET36_XI0/XI21/XI14/MM7_d
+ N_XI0/XI21/XI14/NET35_XI0/XI21/XI14/MM7_g N_VSS_XI0/XI21/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM8 N_XI0/XI21/XI14/NET35_XI0/XI21/XI14/MM8_d
+ N_WL<39>_XI0/XI21/XI14/MM8_g N_BLN<1>_XI0/XI21/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI14/MM5 N_XI0/XI21/XI14/NET34_XI0/XI21/XI14/MM5_d
+ N_XI0/XI21/XI14/NET33_XI0/XI21/XI14/MM5_g N_VDD_XI0/XI21/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI14/MM4 N_XI0/XI21/XI14/NET33_XI0/XI21/XI14/MM4_d
+ N_XI0/XI21/XI14/NET34_XI0/XI21/XI14/MM4_g N_VDD_XI0/XI21/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI14/MM10 N_XI0/XI21/XI14/NET35_XI0/XI21/XI14/MM10_d
+ N_XI0/XI21/XI14/NET36_XI0/XI21/XI14/MM10_g N_VDD_XI0/XI21/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI14/MM11 N_XI0/XI21/XI14/NET36_XI0/XI21/XI14/MM11_d
+ N_XI0/XI21/XI14/NET35_XI0/XI21/XI14/MM11_g N_VDD_XI0/XI21/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI15/MM2 N_XI0/XI21/XI15/NET34_XI0/XI21/XI15/MM2_d
+ N_XI0/XI21/XI15/NET33_XI0/XI21/XI15/MM2_g N_VSS_XI0/XI21/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM3 N_XI0/XI21/XI15/NET33_XI0/XI21/XI15/MM3_d
+ N_WL<38>_XI0/XI21/XI15/MM3_g N_BLN<0>_XI0/XI21/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM0 N_XI0/XI21/XI15/NET34_XI0/XI21/XI15/MM0_d
+ N_WL<38>_XI0/XI21/XI15/MM0_g N_BL<0>_XI0/XI21/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM1 N_XI0/XI21/XI15/NET33_XI0/XI21/XI15/MM1_d
+ N_XI0/XI21/XI15/NET34_XI0/XI21/XI15/MM1_g N_VSS_XI0/XI21/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM9 N_XI0/XI21/XI15/NET36_XI0/XI21/XI15/MM9_d
+ N_WL<39>_XI0/XI21/XI15/MM9_g N_BL<0>_XI0/XI21/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM6 N_XI0/XI21/XI15/NET35_XI0/XI21/XI15/MM6_d
+ N_XI0/XI21/XI15/NET36_XI0/XI21/XI15/MM6_g N_VSS_XI0/XI21/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM7 N_XI0/XI21/XI15/NET36_XI0/XI21/XI15/MM7_d
+ N_XI0/XI21/XI15/NET35_XI0/XI21/XI15/MM7_g N_VSS_XI0/XI21/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM8 N_XI0/XI21/XI15/NET35_XI0/XI21/XI15/MM8_d
+ N_WL<39>_XI0/XI21/XI15/MM8_g N_BLN<0>_XI0/XI21/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI21/XI15/MM5 N_XI0/XI21/XI15/NET34_XI0/XI21/XI15/MM5_d
+ N_XI0/XI21/XI15/NET33_XI0/XI21/XI15/MM5_g N_VDD_XI0/XI21/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI15/MM4 N_XI0/XI21/XI15/NET33_XI0/XI21/XI15/MM4_d
+ N_XI0/XI21/XI15/NET34_XI0/XI21/XI15/MM4_g N_VDD_XI0/XI21/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI15/MM10 N_XI0/XI21/XI15/NET35_XI0/XI21/XI15/MM10_d
+ N_XI0/XI21/XI15/NET36_XI0/XI21/XI15/MM10_g N_VDD_XI0/XI21/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI21/XI15/MM11 N_XI0/XI21/XI15/NET36_XI0/XI21/XI15/MM11_d
+ N_XI0/XI21/XI15/NET35_XI0/XI21/XI15/MM11_g N_VDD_XI0/XI21/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI0/MM2 N_XI0/XI22/XI0/NET34_XI0/XI22/XI0/MM2_d
+ N_XI0/XI22/XI0/NET33_XI0/XI22/XI0/MM2_g N_VSS_XI0/XI22/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM3 N_XI0/XI22/XI0/NET33_XI0/XI22/XI0/MM3_d
+ N_WL<40>_XI0/XI22/XI0/MM3_g N_BLN<15>_XI0/XI22/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM0 N_XI0/XI22/XI0/NET34_XI0/XI22/XI0/MM0_d
+ N_WL<40>_XI0/XI22/XI0/MM0_g N_BL<15>_XI0/XI22/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM1 N_XI0/XI22/XI0/NET33_XI0/XI22/XI0/MM1_d
+ N_XI0/XI22/XI0/NET34_XI0/XI22/XI0/MM1_g N_VSS_XI0/XI22/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM9 N_XI0/XI22/XI0/NET36_XI0/XI22/XI0/MM9_d
+ N_WL<41>_XI0/XI22/XI0/MM9_g N_BL<15>_XI0/XI22/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM6 N_XI0/XI22/XI0/NET35_XI0/XI22/XI0/MM6_d
+ N_XI0/XI22/XI0/NET36_XI0/XI22/XI0/MM6_g N_VSS_XI0/XI22/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM7 N_XI0/XI22/XI0/NET36_XI0/XI22/XI0/MM7_d
+ N_XI0/XI22/XI0/NET35_XI0/XI22/XI0/MM7_g N_VSS_XI0/XI22/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM8 N_XI0/XI22/XI0/NET35_XI0/XI22/XI0/MM8_d
+ N_WL<41>_XI0/XI22/XI0/MM8_g N_BLN<15>_XI0/XI22/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI0/MM5 N_XI0/XI22/XI0/NET34_XI0/XI22/XI0/MM5_d
+ N_XI0/XI22/XI0/NET33_XI0/XI22/XI0/MM5_g N_VDD_XI0/XI22/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI0/MM4 N_XI0/XI22/XI0/NET33_XI0/XI22/XI0/MM4_d
+ N_XI0/XI22/XI0/NET34_XI0/XI22/XI0/MM4_g N_VDD_XI0/XI22/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI0/MM10 N_XI0/XI22/XI0/NET35_XI0/XI22/XI0/MM10_d
+ N_XI0/XI22/XI0/NET36_XI0/XI22/XI0/MM10_g N_VDD_XI0/XI22/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI0/MM11 N_XI0/XI22/XI0/NET36_XI0/XI22/XI0/MM11_d
+ N_XI0/XI22/XI0/NET35_XI0/XI22/XI0/MM11_g N_VDD_XI0/XI22/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI1/MM2 N_XI0/XI22/XI1/NET34_XI0/XI22/XI1/MM2_d
+ N_XI0/XI22/XI1/NET33_XI0/XI22/XI1/MM2_g N_VSS_XI0/XI22/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM3 N_XI0/XI22/XI1/NET33_XI0/XI22/XI1/MM3_d
+ N_WL<40>_XI0/XI22/XI1/MM3_g N_BLN<14>_XI0/XI22/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM0 N_XI0/XI22/XI1/NET34_XI0/XI22/XI1/MM0_d
+ N_WL<40>_XI0/XI22/XI1/MM0_g N_BL<14>_XI0/XI22/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM1 N_XI0/XI22/XI1/NET33_XI0/XI22/XI1/MM1_d
+ N_XI0/XI22/XI1/NET34_XI0/XI22/XI1/MM1_g N_VSS_XI0/XI22/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM9 N_XI0/XI22/XI1/NET36_XI0/XI22/XI1/MM9_d
+ N_WL<41>_XI0/XI22/XI1/MM9_g N_BL<14>_XI0/XI22/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM6 N_XI0/XI22/XI1/NET35_XI0/XI22/XI1/MM6_d
+ N_XI0/XI22/XI1/NET36_XI0/XI22/XI1/MM6_g N_VSS_XI0/XI22/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM7 N_XI0/XI22/XI1/NET36_XI0/XI22/XI1/MM7_d
+ N_XI0/XI22/XI1/NET35_XI0/XI22/XI1/MM7_g N_VSS_XI0/XI22/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM8 N_XI0/XI22/XI1/NET35_XI0/XI22/XI1/MM8_d
+ N_WL<41>_XI0/XI22/XI1/MM8_g N_BLN<14>_XI0/XI22/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI1/MM5 N_XI0/XI22/XI1/NET34_XI0/XI22/XI1/MM5_d
+ N_XI0/XI22/XI1/NET33_XI0/XI22/XI1/MM5_g N_VDD_XI0/XI22/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI1/MM4 N_XI0/XI22/XI1/NET33_XI0/XI22/XI1/MM4_d
+ N_XI0/XI22/XI1/NET34_XI0/XI22/XI1/MM4_g N_VDD_XI0/XI22/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI1/MM10 N_XI0/XI22/XI1/NET35_XI0/XI22/XI1/MM10_d
+ N_XI0/XI22/XI1/NET36_XI0/XI22/XI1/MM10_g N_VDD_XI0/XI22/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI1/MM11 N_XI0/XI22/XI1/NET36_XI0/XI22/XI1/MM11_d
+ N_XI0/XI22/XI1/NET35_XI0/XI22/XI1/MM11_g N_VDD_XI0/XI22/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI2/MM2 N_XI0/XI22/XI2/NET34_XI0/XI22/XI2/MM2_d
+ N_XI0/XI22/XI2/NET33_XI0/XI22/XI2/MM2_g N_VSS_XI0/XI22/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM3 N_XI0/XI22/XI2/NET33_XI0/XI22/XI2/MM3_d
+ N_WL<40>_XI0/XI22/XI2/MM3_g N_BLN<13>_XI0/XI22/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM0 N_XI0/XI22/XI2/NET34_XI0/XI22/XI2/MM0_d
+ N_WL<40>_XI0/XI22/XI2/MM0_g N_BL<13>_XI0/XI22/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM1 N_XI0/XI22/XI2/NET33_XI0/XI22/XI2/MM1_d
+ N_XI0/XI22/XI2/NET34_XI0/XI22/XI2/MM1_g N_VSS_XI0/XI22/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM9 N_XI0/XI22/XI2/NET36_XI0/XI22/XI2/MM9_d
+ N_WL<41>_XI0/XI22/XI2/MM9_g N_BL<13>_XI0/XI22/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM6 N_XI0/XI22/XI2/NET35_XI0/XI22/XI2/MM6_d
+ N_XI0/XI22/XI2/NET36_XI0/XI22/XI2/MM6_g N_VSS_XI0/XI22/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM7 N_XI0/XI22/XI2/NET36_XI0/XI22/XI2/MM7_d
+ N_XI0/XI22/XI2/NET35_XI0/XI22/XI2/MM7_g N_VSS_XI0/XI22/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM8 N_XI0/XI22/XI2/NET35_XI0/XI22/XI2/MM8_d
+ N_WL<41>_XI0/XI22/XI2/MM8_g N_BLN<13>_XI0/XI22/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI2/MM5 N_XI0/XI22/XI2/NET34_XI0/XI22/XI2/MM5_d
+ N_XI0/XI22/XI2/NET33_XI0/XI22/XI2/MM5_g N_VDD_XI0/XI22/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI2/MM4 N_XI0/XI22/XI2/NET33_XI0/XI22/XI2/MM4_d
+ N_XI0/XI22/XI2/NET34_XI0/XI22/XI2/MM4_g N_VDD_XI0/XI22/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI2/MM10 N_XI0/XI22/XI2/NET35_XI0/XI22/XI2/MM10_d
+ N_XI0/XI22/XI2/NET36_XI0/XI22/XI2/MM10_g N_VDD_XI0/XI22/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI2/MM11 N_XI0/XI22/XI2/NET36_XI0/XI22/XI2/MM11_d
+ N_XI0/XI22/XI2/NET35_XI0/XI22/XI2/MM11_g N_VDD_XI0/XI22/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI3/MM2 N_XI0/XI22/XI3/NET34_XI0/XI22/XI3/MM2_d
+ N_XI0/XI22/XI3/NET33_XI0/XI22/XI3/MM2_g N_VSS_XI0/XI22/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM3 N_XI0/XI22/XI3/NET33_XI0/XI22/XI3/MM3_d
+ N_WL<40>_XI0/XI22/XI3/MM3_g N_BLN<12>_XI0/XI22/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM0 N_XI0/XI22/XI3/NET34_XI0/XI22/XI3/MM0_d
+ N_WL<40>_XI0/XI22/XI3/MM0_g N_BL<12>_XI0/XI22/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM1 N_XI0/XI22/XI3/NET33_XI0/XI22/XI3/MM1_d
+ N_XI0/XI22/XI3/NET34_XI0/XI22/XI3/MM1_g N_VSS_XI0/XI22/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM9 N_XI0/XI22/XI3/NET36_XI0/XI22/XI3/MM9_d
+ N_WL<41>_XI0/XI22/XI3/MM9_g N_BL<12>_XI0/XI22/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM6 N_XI0/XI22/XI3/NET35_XI0/XI22/XI3/MM6_d
+ N_XI0/XI22/XI3/NET36_XI0/XI22/XI3/MM6_g N_VSS_XI0/XI22/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM7 N_XI0/XI22/XI3/NET36_XI0/XI22/XI3/MM7_d
+ N_XI0/XI22/XI3/NET35_XI0/XI22/XI3/MM7_g N_VSS_XI0/XI22/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM8 N_XI0/XI22/XI3/NET35_XI0/XI22/XI3/MM8_d
+ N_WL<41>_XI0/XI22/XI3/MM8_g N_BLN<12>_XI0/XI22/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI3/MM5 N_XI0/XI22/XI3/NET34_XI0/XI22/XI3/MM5_d
+ N_XI0/XI22/XI3/NET33_XI0/XI22/XI3/MM5_g N_VDD_XI0/XI22/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI3/MM4 N_XI0/XI22/XI3/NET33_XI0/XI22/XI3/MM4_d
+ N_XI0/XI22/XI3/NET34_XI0/XI22/XI3/MM4_g N_VDD_XI0/XI22/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI3/MM10 N_XI0/XI22/XI3/NET35_XI0/XI22/XI3/MM10_d
+ N_XI0/XI22/XI3/NET36_XI0/XI22/XI3/MM10_g N_VDD_XI0/XI22/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI3/MM11 N_XI0/XI22/XI3/NET36_XI0/XI22/XI3/MM11_d
+ N_XI0/XI22/XI3/NET35_XI0/XI22/XI3/MM11_g N_VDD_XI0/XI22/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI4/MM2 N_XI0/XI22/XI4/NET34_XI0/XI22/XI4/MM2_d
+ N_XI0/XI22/XI4/NET33_XI0/XI22/XI4/MM2_g N_VSS_XI0/XI22/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM3 N_XI0/XI22/XI4/NET33_XI0/XI22/XI4/MM3_d
+ N_WL<40>_XI0/XI22/XI4/MM3_g N_BLN<11>_XI0/XI22/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM0 N_XI0/XI22/XI4/NET34_XI0/XI22/XI4/MM0_d
+ N_WL<40>_XI0/XI22/XI4/MM0_g N_BL<11>_XI0/XI22/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM1 N_XI0/XI22/XI4/NET33_XI0/XI22/XI4/MM1_d
+ N_XI0/XI22/XI4/NET34_XI0/XI22/XI4/MM1_g N_VSS_XI0/XI22/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM9 N_XI0/XI22/XI4/NET36_XI0/XI22/XI4/MM9_d
+ N_WL<41>_XI0/XI22/XI4/MM9_g N_BL<11>_XI0/XI22/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM6 N_XI0/XI22/XI4/NET35_XI0/XI22/XI4/MM6_d
+ N_XI0/XI22/XI4/NET36_XI0/XI22/XI4/MM6_g N_VSS_XI0/XI22/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM7 N_XI0/XI22/XI4/NET36_XI0/XI22/XI4/MM7_d
+ N_XI0/XI22/XI4/NET35_XI0/XI22/XI4/MM7_g N_VSS_XI0/XI22/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM8 N_XI0/XI22/XI4/NET35_XI0/XI22/XI4/MM8_d
+ N_WL<41>_XI0/XI22/XI4/MM8_g N_BLN<11>_XI0/XI22/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI4/MM5 N_XI0/XI22/XI4/NET34_XI0/XI22/XI4/MM5_d
+ N_XI0/XI22/XI4/NET33_XI0/XI22/XI4/MM5_g N_VDD_XI0/XI22/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI4/MM4 N_XI0/XI22/XI4/NET33_XI0/XI22/XI4/MM4_d
+ N_XI0/XI22/XI4/NET34_XI0/XI22/XI4/MM4_g N_VDD_XI0/XI22/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI4/MM10 N_XI0/XI22/XI4/NET35_XI0/XI22/XI4/MM10_d
+ N_XI0/XI22/XI4/NET36_XI0/XI22/XI4/MM10_g N_VDD_XI0/XI22/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI4/MM11 N_XI0/XI22/XI4/NET36_XI0/XI22/XI4/MM11_d
+ N_XI0/XI22/XI4/NET35_XI0/XI22/XI4/MM11_g N_VDD_XI0/XI22/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI5/MM2 N_XI0/XI22/XI5/NET34_XI0/XI22/XI5/MM2_d
+ N_XI0/XI22/XI5/NET33_XI0/XI22/XI5/MM2_g N_VSS_XI0/XI22/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM3 N_XI0/XI22/XI5/NET33_XI0/XI22/XI5/MM3_d
+ N_WL<40>_XI0/XI22/XI5/MM3_g N_BLN<10>_XI0/XI22/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM0 N_XI0/XI22/XI5/NET34_XI0/XI22/XI5/MM0_d
+ N_WL<40>_XI0/XI22/XI5/MM0_g N_BL<10>_XI0/XI22/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM1 N_XI0/XI22/XI5/NET33_XI0/XI22/XI5/MM1_d
+ N_XI0/XI22/XI5/NET34_XI0/XI22/XI5/MM1_g N_VSS_XI0/XI22/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM9 N_XI0/XI22/XI5/NET36_XI0/XI22/XI5/MM9_d
+ N_WL<41>_XI0/XI22/XI5/MM9_g N_BL<10>_XI0/XI22/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM6 N_XI0/XI22/XI5/NET35_XI0/XI22/XI5/MM6_d
+ N_XI0/XI22/XI5/NET36_XI0/XI22/XI5/MM6_g N_VSS_XI0/XI22/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM7 N_XI0/XI22/XI5/NET36_XI0/XI22/XI5/MM7_d
+ N_XI0/XI22/XI5/NET35_XI0/XI22/XI5/MM7_g N_VSS_XI0/XI22/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM8 N_XI0/XI22/XI5/NET35_XI0/XI22/XI5/MM8_d
+ N_WL<41>_XI0/XI22/XI5/MM8_g N_BLN<10>_XI0/XI22/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI5/MM5 N_XI0/XI22/XI5/NET34_XI0/XI22/XI5/MM5_d
+ N_XI0/XI22/XI5/NET33_XI0/XI22/XI5/MM5_g N_VDD_XI0/XI22/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI5/MM4 N_XI0/XI22/XI5/NET33_XI0/XI22/XI5/MM4_d
+ N_XI0/XI22/XI5/NET34_XI0/XI22/XI5/MM4_g N_VDD_XI0/XI22/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI5/MM10 N_XI0/XI22/XI5/NET35_XI0/XI22/XI5/MM10_d
+ N_XI0/XI22/XI5/NET36_XI0/XI22/XI5/MM10_g N_VDD_XI0/XI22/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI5/MM11 N_XI0/XI22/XI5/NET36_XI0/XI22/XI5/MM11_d
+ N_XI0/XI22/XI5/NET35_XI0/XI22/XI5/MM11_g N_VDD_XI0/XI22/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI6/MM2 N_XI0/XI22/XI6/NET34_XI0/XI22/XI6/MM2_d
+ N_XI0/XI22/XI6/NET33_XI0/XI22/XI6/MM2_g N_VSS_XI0/XI22/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM3 N_XI0/XI22/XI6/NET33_XI0/XI22/XI6/MM3_d
+ N_WL<40>_XI0/XI22/XI6/MM3_g N_BLN<9>_XI0/XI22/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM0 N_XI0/XI22/XI6/NET34_XI0/XI22/XI6/MM0_d
+ N_WL<40>_XI0/XI22/XI6/MM0_g N_BL<9>_XI0/XI22/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM1 N_XI0/XI22/XI6/NET33_XI0/XI22/XI6/MM1_d
+ N_XI0/XI22/XI6/NET34_XI0/XI22/XI6/MM1_g N_VSS_XI0/XI22/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM9 N_XI0/XI22/XI6/NET36_XI0/XI22/XI6/MM9_d
+ N_WL<41>_XI0/XI22/XI6/MM9_g N_BL<9>_XI0/XI22/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM6 N_XI0/XI22/XI6/NET35_XI0/XI22/XI6/MM6_d
+ N_XI0/XI22/XI6/NET36_XI0/XI22/XI6/MM6_g N_VSS_XI0/XI22/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM7 N_XI0/XI22/XI6/NET36_XI0/XI22/XI6/MM7_d
+ N_XI0/XI22/XI6/NET35_XI0/XI22/XI6/MM7_g N_VSS_XI0/XI22/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM8 N_XI0/XI22/XI6/NET35_XI0/XI22/XI6/MM8_d
+ N_WL<41>_XI0/XI22/XI6/MM8_g N_BLN<9>_XI0/XI22/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI6/MM5 N_XI0/XI22/XI6/NET34_XI0/XI22/XI6/MM5_d
+ N_XI0/XI22/XI6/NET33_XI0/XI22/XI6/MM5_g N_VDD_XI0/XI22/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI6/MM4 N_XI0/XI22/XI6/NET33_XI0/XI22/XI6/MM4_d
+ N_XI0/XI22/XI6/NET34_XI0/XI22/XI6/MM4_g N_VDD_XI0/XI22/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI6/MM10 N_XI0/XI22/XI6/NET35_XI0/XI22/XI6/MM10_d
+ N_XI0/XI22/XI6/NET36_XI0/XI22/XI6/MM10_g N_VDD_XI0/XI22/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI6/MM11 N_XI0/XI22/XI6/NET36_XI0/XI22/XI6/MM11_d
+ N_XI0/XI22/XI6/NET35_XI0/XI22/XI6/MM11_g N_VDD_XI0/XI22/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI7/MM2 N_XI0/XI22/XI7/NET34_XI0/XI22/XI7/MM2_d
+ N_XI0/XI22/XI7/NET33_XI0/XI22/XI7/MM2_g N_VSS_XI0/XI22/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM3 N_XI0/XI22/XI7/NET33_XI0/XI22/XI7/MM3_d
+ N_WL<40>_XI0/XI22/XI7/MM3_g N_BLN<8>_XI0/XI22/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM0 N_XI0/XI22/XI7/NET34_XI0/XI22/XI7/MM0_d
+ N_WL<40>_XI0/XI22/XI7/MM0_g N_BL<8>_XI0/XI22/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM1 N_XI0/XI22/XI7/NET33_XI0/XI22/XI7/MM1_d
+ N_XI0/XI22/XI7/NET34_XI0/XI22/XI7/MM1_g N_VSS_XI0/XI22/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM9 N_XI0/XI22/XI7/NET36_XI0/XI22/XI7/MM9_d
+ N_WL<41>_XI0/XI22/XI7/MM9_g N_BL<8>_XI0/XI22/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM6 N_XI0/XI22/XI7/NET35_XI0/XI22/XI7/MM6_d
+ N_XI0/XI22/XI7/NET36_XI0/XI22/XI7/MM6_g N_VSS_XI0/XI22/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM7 N_XI0/XI22/XI7/NET36_XI0/XI22/XI7/MM7_d
+ N_XI0/XI22/XI7/NET35_XI0/XI22/XI7/MM7_g N_VSS_XI0/XI22/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM8 N_XI0/XI22/XI7/NET35_XI0/XI22/XI7/MM8_d
+ N_WL<41>_XI0/XI22/XI7/MM8_g N_BLN<8>_XI0/XI22/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI7/MM5 N_XI0/XI22/XI7/NET34_XI0/XI22/XI7/MM5_d
+ N_XI0/XI22/XI7/NET33_XI0/XI22/XI7/MM5_g N_VDD_XI0/XI22/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI7/MM4 N_XI0/XI22/XI7/NET33_XI0/XI22/XI7/MM4_d
+ N_XI0/XI22/XI7/NET34_XI0/XI22/XI7/MM4_g N_VDD_XI0/XI22/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI7/MM10 N_XI0/XI22/XI7/NET35_XI0/XI22/XI7/MM10_d
+ N_XI0/XI22/XI7/NET36_XI0/XI22/XI7/MM10_g N_VDD_XI0/XI22/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI7/MM11 N_XI0/XI22/XI7/NET36_XI0/XI22/XI7/MM11_d
+ N_XI0/XI22/XI7/NET35_XI0/XI22/XI7/MM11_g N_VDD_XI0/XI22/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI8/MM2 N_XI0/XI22/XI8/NET34_XI0/XI22/XI8/MM2_d
+ N_XI0/XI22/XI8/NET33_XI0/XI22/XI8/MM2_g N_VSS_XI0/XI22/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM3 N_XI0/XI22/XI8/NET33_XI0/XI22/XI8/MM3_d
+ N_WL<40>_XI0/XI22/XI8/MM3_g N_BLN<7>_XI0/XI22/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM0 N_XI0/XI22/XI8/NET34_XI0/XI22/XI8/MM0_d
+ N_WL<40>_XI0/XI22/XI8/MM0_g N_BL<7>_XI0/XI22/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM1 N_XI0/XI22/XI8/NET33_XI0/XI22/XI8/MM1_d
+ N_XI0/XI22/XI8/NET34_XI0/XI22/XI8/MM1_g N_VSS_XI0/XI22/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM9 N_XI0/XI22/XI8/NET36_XI0/XI22/XI8/MM9_d
+ N_WL<41>_XI0/XI22/XI8/MM9_g N_BL<7>_XI0/XI22/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM6 N_XI0/XI22/XI8/NET35_XI0/XI22/XI8/MM6_d
+ N_XI0/XI22/XI8/NET36_XI0/XI22/XI8/MM6_g N_VSS_XI0/XI22/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM7 N_XI0/XI22/XI8/NET36_XI0/XI22/XI8/MM7_d
+ N_XI0/XI22/XI8/NET35_XI0/XI22/XI8/MM7_g N_VSS_XI0/XI22/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM8 N_XI0/XI22/XI8/NET35_XI0/XI22/XI8/MM8_d
+ N_WL<41>_XI0/XI22/XI8/MM8_g N_BLN<7>_XI0/XI22/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI8/MM5 N_XI0/XI22/XI8/NET34_XI0/XI22/XI8/MM5_d
+ N_XI0/XI22/XI8/NET33_XI0/XI22/XI8/MM5_g N_VDD_XI0/XI22/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI8/MM4 N_XI0/XI22/XI8/NET33_XI0/XI22/XI8/MM4_d
+ N_XI0/XI22/XI8/NET34_XI0/XI22/XI8/MM4_g N_VDD_XI0/XI22/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI8/MM10 N_XI0/XI22/XI8/NET35_XI0/XI22/XI8/MM10_d
+ N_XI0/XI22/XI8/NET36_XI0/XI22/XI8/MM10_g N_VDD_XI0/XI22/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI8/MM11 N_XI0/XI22/XI8/NET36_XI0/XI22/XI8/MM11_d
+ N_XI0/XI22/XI8/NET35_XI0/XI22/XI8/MM11_g N_VDD_XI0/XI22/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI9/MM2 N_XI0/XI22/XI9/NET34_XI0/XI22/XI9/MM2_d
+ N_XI0/XI22/XI9/NET33_XI0/XI22/XI9/MM2_g N_VSS_XI0/XI22/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM3 N_XI0/XI22/XI9/NET33_XI0/XI22/XI9/MM3_d
+ N_WL<40>_XI0/XI22/XI9/MM3_g N_BLN<6>_XI0/XI22/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM0 N_XI0/XI22/XI9/NET34_XI0/XI22/XI9/MM0_d
+ N_WL<40>_XI0/XI22/XI9/MM0_g N_BL<6>_XI0/XI22/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM1 N_XI0/XI22/XI9/NET33_XI0/XI22/XI9/MM1_d
+ N_XI0/XI22/XI9/NET34_XI0/XI22/XI9/MM1_g N_VSS_XI0/XI22/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM9 N_XI0/XI22/XI9/NET36_XI0/XI22/XI9/MM9_d
+ N_WL<41>_XI0/XI22/XI9/MM9_g N_BL<6>_XI0/XI22/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM6 N_XI0/XI22/XI9/NET35_XI0/XI22/XI9/MM6_d
+ N_XI0/XI22/XI9/NET36_XI0/XI22/XI9/MM6_g N_VSS_XI0/XI22/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM7 N_XI0/XI22/XI9/NET36_XI0/XI22/XI9/MM7_d
+ N_XI0/XI22/XI9/NET35_XI0/XI22/XI9/MM7_g N_VSS_XI0/XI22/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM8 N_XI0/XI22/XI9/NET35_XI0/XI22/XI9/MM8_d
+ N_WL<41>_XI0/XI22/XI9/MM8_g N_BLN<6>_XI0/XI22/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI9/MM5 N_XI0/XI22/XI9/NET34_XI0/XI22/XI9/MM5_d
+ N_XI0/XI22/XI9/NET33_XI0/XI22/XI9/MM5_g N_VDD_XI0/XI22/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI9/MM4 N_XI0/XI22/XI9/NET33_XI0/XI22/XI9/MM4_d
+ N_XI0/XI22/XI9/NET34_XI0/XI22/XI9/MM4_g N_VDD_XI0/XI22/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI9/MM10 N_XI0/XI22/XI9/NET35_XI0/XI22/XI9/MM10_d
+ N_XI0/XI22/XI9/NET36_XI0/XI22/XI9/MM10_g N_VDD_XI0/XI22/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI9/MM11 N_XI0/XI22/XI9/NET36_XI0/XI22/XI9/MM11_d
+ N_XI0/XI22/XI9/NET35_XI0/XI22/XI9/MM11_g N_VDD_XI0/XI22/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI10/MM2 N_XI0/XI22/XI10/NET34_XI0/XI22/XI10/MM2_d
+ N_XI0/XI22/XI10/NET33_XI0/XI22/XI10/MM2_g N_VSS_XI0/XI22/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM3 N_XI0/XI22/XI10/NET33_XI0/XI22/XI10/MM3_d
+ N_WL<40>_XI0/XI22/XI10/MM3_g N_BLN<5>_XI0/XI22/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM0 N_XI0/XI22/XI10/NET34_XI0/XI22/XI10/MM0_d
+ N_WL<40>_XI0/XI22/XI10/MM0_g N_BL<5>_XI0/XI22/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM1 N_XI0/XI22/XI10/NET33_XI0/XI22/XI10/MM1_d
+ N_XI0/XI22/XI10/NET34_XI0/XI22/XI10/MM1_g N_VSS_XI0/XI22/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM9 N_XI0/XI22/XI10/NET36_XI0/XI22/XI10/MM9_d
+ N_WL<41>_XI0/XI22/XI10/MM9_g N_BL<5>_XI0/XI22/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM6 N_XI0/XI22/XI10/NET35_XI0/XI22/XI10/MM6_d
+ N_XI0/XI22/XI10/NET36_XI0/XI22/XI10/MM6_g N_VSS_XI0/XI22/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM7 N_XI0/XI22/XI10/NET36_XI0/XI22/XI10/MM7_d
+ N_XI0/XI22/XI10/NET35_XI0/XI22/XI10/MM7_g N_VSS_XI0/XI22/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM8 N_XI0/XI22/XI10/NET35_XI0/XI22/XI10/MM8_d
+ N_WL<41>_XI0/XI22/XI10/MM8_g N_BLN<5>_XI0/XI22/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI10/MM5 N_XI0/XI22/XI10/NET34_XI0/XI22/XI10/MM5_d
+ N_XI0/XI22/XI10/NET33_XI0/XI22/XI10/MM5_g N_VDD_XI0/XI22/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI10/MM4 N_XI0/XI22/XI10/NET33_XI0/XI22/XI10/MM4_d
+ N_XI0/XI22/XI10/NET34_XI0/XI22/XI10/MM4_g N_VDD_XI0/XI22/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI10/MM10 N_XI0/XI22/XI10/NET35_XI0/XI22/XI10/MM10_d
+ N_XI0/XI22/XI10/NET36_XI0/XI22/XI10/MM10_g N_VDD_XI0/XI22/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI10/MM11 N_XI0/XI22/XI10/NET36_XI0/XI22/XI10/MM11_d
+ N_XI0/XI22/XI10/NET35_XI0/XI22/XI10/MM11_g N_VDD_XI0/XI22/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI11/MM2 N_XI0/XI22/XI11/NET34_XI0/XI22/XI11/MM2_d
+ N_XI0/XI22/XI11/NET33_XI0/XI22/XI11/MM2_g N_VSS_XI0/XI22/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM3 N_XI0/XI22/XI11/NET33_XI0/XI22/XI11/MM3_d
+ N_WL<40>_XI0/XI22/XI11/MM3_g N_BLN<4>_XI0/XI22/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM0 N_XI0/XI22/XI11/NET34_XI0/XI22/XI11/MM0_d
+ N_WL<40>_XI0/XI22/XI11/MM0_g N_BL<4>_XI0/XI22/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM1 N_XI0/XI22/XI11/NET33_XI0/XI22/XI11/MM1_d
+ N_XI0/XI22/XI11/NET34_XI0/XI22/XI11/MM1_g N_VSS_XI0/XI22/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM9 N_XI0/XI22/XI11/NET36_XI0/XI22/XI11/MM9_d
+ N_WL<41>_XI0/XI22/XI11/MM9_g N_BL<4>_XI0/XI22/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM6 N_XI0/XI22/XI11/NET35_XI0/XI22/XI11/MM6_d
+ N_XI0/XI22/XI11/NET36_XI0/XI22/XI11/MM6_g N_VSS_XI0/XI22/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM7 N_XI0/XI22/XI11/NET36_XI0/XI22/XI11/MM7_d
+ N_XI0/XI22/XI11/NET35_XI0/XI22/XI11/MM7_g N_VSS_XI0/XI22/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM8 N_XI0/XI22/XI11/NET35_XI0/XI22/XI11/MM8_d
+ N_WL<41>_XI0/XI22/XI11/MM8_g N_BLN<4>_XI0/XI22/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI11/MM5 N_XI0/XI22/XI11/NET34_XI0/XI22/XI11/MM5_d
+ N_XI0/XI22/XI11/NET33_XI0/XI22/XI11/MM5_g N_VDD_XI0/XI22/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI11/MM4 N_XI0/XI22/XI11/NET33_XI0/XI22/XI11/MM4_d
+ N_XI0/XI22/XI11/NET34_XI0/XI22/XI11/MM4_g N_VDD_XI0/XI22/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI11/MM10 N_XI0/XI22/XI11/NET35_XI0/XI22/XI11/MM10_d
+ N_XI0/XI22/XI11/NET36_XI0/XI22/XI11/MM10_g N_VDD_XI0/XI22/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI11/MM11 N_XI0/XI22/XI11/NET36_XI0/XI22/XI11/MM11_d
+ N_XI0/XI22/XI11/NET35_XI0/XI22/XI11/MM11_g N_VDD_XI0/XI22/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI12/MM2 N_XI0/XI22/XI12/NET34_XI0/XI22/XI12/MM2_d
+ N_XI0/XI22/XI12/NET33_XI0/XI22/XI12/MM2_g N_VSS_XI0/XI22/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM3 N_XI0/XI22/XI12/NET33_XI0/XI22/XI12/MM3_d
+ N_WL<40>_XI0/XI22/XI12/MM3_g N_BLN<3>_XI0/XI22/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM0 N_XI0/XI22/XI12/NET34_XI0/XI22/XI12/MM0_d
+ N_WL<40>_XI0/XI22/XI12/MM0_g N_BL<3>_XI0/XI22/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM1 N_XI0/XI22/XI12/NET33_XI0/XI22/XI12/MM1_d
+ N_XI0/XI22/XI12/NET34_XI0/XI22/XI12/MM1_g N_VSS_XI0/XI22/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM9 N_XI0/XI22/XI12/NET36_XI0/XI22/XI12/MM9_d
+ N_WL<41>_XI0/XI22/XI12/MM9_g N_BL<3>_XI0/XI22/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM6 N_XI0/XI22/XI12/NET35_XI0/XI22/XI12/MM6_d
+ N_XI0/XI22/XI12/NET36_XI0/XI22/XI12/MM6_g N_VSS_XI0/XI22/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM7 N_XI0/XI22/XI12/NET36_XI0/XI22/XI12/MM7_d
+ N_XI0/XI22/XI12/NET35_XI0/XI22/XI12/MM7_g N_VSS_XI0/XI22/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM8 N_XI0/XI22/XI12/NET35_XI0/XI22/XI12/MM8_d
+ N_WL<41>_XI0/XI22/XI12/MM8_g N_BLN<3>_XI0/XI22/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI12/MM5 N_XI0/XI22/XI12/NET34_XI0/XI22/XI12/MM5_d
+ N_XI0/XI22/XI12/NET33_XI0/XI22/XI12/MM5_g N_VDD_XI0/XI22/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI12/MM4 N_XI0/XI22/XI12/NET33_XI0/XI22/XI12/MM4_d
+ N_XI0/XI22/XI12/NET34_XI0/XI22/XI12/MM4_g N_VDD_XI0/XI22/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI12/MM10 N_XI0/XI22/XI12/NET35_XI0/XI22/XI12/MM10_d
+ N_XI0/XI22/XI12/NET36_XI0/XI22/XI12/MM10_g N_VDD_XI0/XI22/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI12/MM11 N_XI0/XI22/XI12/NET36_XI0/XI22/XI12/MM11_d
+ N_XI0/XI22/XI12/NET35_XI0/XI22/XI12/MM11_g N_VDD_XI0/XI22/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI13/MM2 N_XI0/XI22/XI13/NET34_XI0/XI22/XI13/MM2_d
+ N_XI0/XI22/XI13/NET33_XI0/XI22/XI13/MM2_g N_VSS_XI0/XI22/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM3 N_XI0/XI22/XI13/NET33_XI0/XI22/XI13/MM3_d
+ N_WL<40>_XI0/XI22/XI13/MM3_g N_BLN<2>_XI0/XI22/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM0 N_XI0/XI22/XI13/NET34_XI0/XI22/XI13/MM0_d
+ N_WL<40>_XI0/XI22/XI13/MM0_g N_BL<2>_XI0/XI22/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM1 N_XI0/XI22/XI13/NET33_XI0/XI22/XI13/MM1_d
+ N_XI0/XI22/XI13/NET34_XI0/XI22/XI13/MM1_g N_VSS_XI0/XI22/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM9 N_XI0/XI22/XI13/NET36_XI0/XI22/XI13/MM9_d
+ N_WL<41>_XI0/XI22/XI13/MM9_g N_BL<2>_XI0/XI22/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM6 N_XI0/XI22/XI13/NET35_XI0/XI22/XI13/MM6_d
+ N_XI0/XI22/XI13/NET36_XI0/XI22/XI13/MM6_g N_VSS_XI0/XI22/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM7 N_XI0/XI22/XI13/NET36_XI0/XI22/XI13/MM7_d
+ N_XI0/XI22/XI13/NET35_XI0/XI22/XI13/MM7_g N_VSS_XI0/XI22/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM8 N_XI0/XI22/XI13/NET35_XI0/XI22/XI13/MM8_d
+ N_WL<41>_XI0/XI22/XI13/MM8_g N_BLN<2>_XI0/XI22/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI13/MM5 N_XI0/XI22/XI13/NET34_XI0/XI22/XI13/MM5_d
+ N_XI0/XI22/XI13/NET33_XI0/XI22/XI13/MM5_g N_VDD_XI0/XI22/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI13/MM4 N_XI0/XI22/XI13/NET33_XI0/XI22/XI13/MM4_d
+ N_XI0/XI22/XI13/NET34_XI0/XI22/XI13/MM4_g N_VDD_XI0/XI22/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI13/MM10 N_XI0/XI22/XI13/NET35_XI0/XI22/XI13/MM10_d
+ N_XI0/XI22/XI13/NET36_XI0/XI22/XI13/MM10_g N_VDD_XI0/XI22/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI13/MM11 N_XI0/XI22/XI13/NET36_XI0/XI22/XI13/MM11_d
+ N_XI0/XI22/XI13/NET35_XI0/XI22/XI13/MM11_g N_VDD_XI0/XI22/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI14/MM2 N_XI0/XI22/XI14/NET34_XI0/XI22/XI14/MM2_d
+ N_XI0/XI22/XI14/NET33_XI0/XI22/XI14/MM2_g N_VSS_XI0/XI22/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM3 N_XI0/XI22/XI14/NET33_XI0/XI22/XI14/MM3_d
+ N_WL<40>_XI0/XI22/XI14/MM3_g N_BLN<1>_XI0/XI22/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM0 N_XI0/XI22/XI14/NET34_XI0/XI22/XI14/MM0_d
+ N_WL<40>_XI0/XI22/XI14/MM0_g N_BL<1>_XI0/XI22/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM1 N_XI0/XI22/XI14/NET33_XI0/XI22/XI14/MM1_d
+ N_XI0/XI22/XI14/NET34_XI0/XI22/XI14/MM1_g N_VSS_XI0/XI22/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM9 N_XI0/XI22/XI14/NET36_XI0/XI22/XI14/MM9_d
+ N_WL<41>_XI0/XI22/XI14/MM9_g N_BL<1>_XI0/XI22/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM6 N_XI0/XI22/XI14/NET35_XI0/XI22/XI14/MM6_d
+ N_XI0/XI22/XI14/NET36_XI0/XI22/XI14/MM6_g N_VSS_XI0/XI22/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM7 N_XI0/XI22/XI14/NET36_XI0/XI22/XI14/MM7_d
+ N_XI0/XI22/XI14/NET35_XI0/XI22/XI14/MM7_g N_VSS_XI0/XI22/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM8 N_XI0/XI22/XI14/NET35_XI0/XI22/XI14/MM8_d
+ N_WL<41>_XI0/XI22/XI14/MM8_g N_BLN<1>_XI0/XI22/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI14/MM5 N_XI0/XI22/XI14/NET34_XI0/XI22/XI14/MM5_d
+ N_XI0/XI22/XI14/NET33_XI0/XI22/XI14/MM5_g N_VDD_XI0/XI22/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI14/MM4 N_XI0/XI22/XI14/NET33_XI0/XI22/XI14/MM4_d
+ N_XI0/XI22/XI14/NET34_XI0/XI22/XI14/MM4_g N_VDD_XI0/XI22/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI14/MM10 N_XI0/XI22/XI14/NET35_XI0/XI22/XI14/MM10_d
+ N_XI0/XI22/XI14/NET36_XI0/XI22/XI14/MM10_g N_VDD_XI0/XI22/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI14/MM11 N_XI0/XI22/XI14/NET36_XI0/XI22/XI14/MM11_d
+ N_XI0/XI22/XI14/NET35_XI0/XI22/XI14/MM11_g N_VDD_XI0/XI22/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI15/MM2 N_XI0/XI22/XI15/NET34_XI0/XI22/XI15/MM2_d
+ N_XI0/XI22/XI15/NET33_XI0/XI22/XI15/MM2_g N_VSS_XI0/XI22/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM3 N_XI0/XI22/XI15/NET33_XI0/XI22/XI15/MM3_d
+ N_WL<40>_XI0/XI22/XI15/MM3_g N_BLN<0>_XI0/XI22/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM0 N_XI0/XI22/XI15/NET34_XI0/XI22/XI15/MM0_d
+ N_WL<40>_XI0/XI22/XI15/MM0_g N_BL<0>_XI0/XI22/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM1 N_XI0/XI22/XI15/NET33_XI0/XI22/XI15/MM1_d
+ N_XI0/XI22/XI15/NET34_XI0/XI22/XI15/MM1_g N_VSS_XI0/XI22/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM9 N_XI0/XI22/XI15/NET36_XI0/XI22/XI15/MM9_d
+ N_WL<41>_XI0/XI22/XI15/MM9_g N_BL<0>_XI0/XI22/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM6 N_XI0/XI22/XI15/NET35_XI0/XI22/XI15/MM6_d
+ N_XI0/XI22/XI15/NET36_XI0/XI22/XI15/MM6_g N_VSS_XI0/XI22/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM7 N_XI0/XI22/XI15/NET36_XI0/XI22/XI15/MM7_d
+ N_XI0/XI22/XI15/NET35_XI0/XI22/XI15/MM7_g N_VSS_XI0/XI22/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM8 N_XI0/XI22/XI15/NET35_XI0/XI22/XI15/MM8_d
+ N_WL<41>_XI0/XI22/XI15/MM8_g N_BLN<0>_XI0/XI22/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI22/XI15/MM5 N_XI0/XI22/XI15/NET34_XI0/XI22/XI15/MM5_d
+ N_XI0/XI22/XI15/NET33_XI0/XI22/XI15/MM5_g N_VDD_XI0/XI22/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI15/MM4 N_XI0/XI22/XI15/NET33_XI0/XI22/XI15/MM4_d
+ N_XI0/XI22/XI15/NET34_XI0/XI22/XI15/MM4_g N_VDD_XI0/XI22/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI15/MM10 N_XI0/XI22/XI15/NET35_XI0/XI22/XI15/MM10_d
+ N_XI0/XI22/XI15/NET36_XI0/XI22/XI15/MM10_g N_VDD_XI0/XI22/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI22/XI15/MM11 N_XI0/XI22/XI15/NET36_XI0/XI22/XI15/MM11_d
+ N_XI0/XI22/XI15/NET35_XI0/XI22/XI15/MM11_g N_VDD_XI0/XI22/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI0/MM2 N_XI0/XI23/XI0/NET34_XI0/XI23/XI0/MM2_d
+ N_XI0/XI23/XI0/NET33_XI0/XI23/XI0/MM2_g N_VSS_XI0/XI23/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM3 N_XI0/XI23/XI0/NET33_XI0/XI23/XI0/MM3_d
+ N_WL<42>_XI0/XI23/XI0/MM3_g N_BLN<15>_XI0/XI23/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM0 N_XI0/XI23/XI0/NET34_XI0/XI23/XI0/MM0_d
+ N_WL<42>_XI0/XI23/XI0/MM0_g N_BL<15>_XI0/XI23/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM1 N_XI0/XI23/XI0/NET33_XI0/XI23/XI0/MM1_d
+ N_XI0/XI23/XI0/NET34_XI0/XI23/XI0/MM1_g N_VSS_XI0/XI23/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM9 N_XI0/XI23/XI0/NET36_XI0/XI23/XI0/MM9_d
+ N_WL<43>_XI0/XI23/XI0/MM9_g N_BL<15>_XI0/XI23/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM6 N_XI0/XI23/XI0/NET35_XI0/XI23/XI0/MM6_d
+ N_XI0/XI23/XI0/NET36_XI0/XI23/XI0/MM6_g N_VSS_XI0/XI23/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM7 N_XI0/XI23/XI0/NET36_XI0/XI23/XI0/MM7_d
+ N_XI0/XI23/XI0/NET35_XI0/XI23/XI0/MM7_g N_VSS_XI0/XI23/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM8 N_XI0/XI23/XI0/NET35_XI0/XI23/XI0/MM8_d
+ N_WL<43>_XI0/XI23/XI0/MM8_g N_BLN<15>_XI0/XI23/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI0/MM5 N_XI0/XI23/XI0/NET34_XI0/XI23/XI0/MM5_d
+ N_XI0/XI23/XI0/NET33_XI0/XI23/XI0/MM5_g N_VDD_XI0/XI23/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI0/MM4 N_XI0/XI23/XI0/NET33_XI0/XI23/XI0/MM4_d
+ N_XI0/XI23/XI0/NET34_XI0/XI23/XI0/MM4_g N_VDD_XI0/XI23/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI0/MM10 N_XI0/XI23/XI0/NET35_XI0/XI23/XI0/MM10_d
+ N_XI0/XI23/XI0/NET36_XI0/XI23/XI0/MM10_g N_VDD_XI0/XI23/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI0/MM11 N_XI0/XI23/XI0/NET36_XI0/XI23/XI0/MM11_d
+ N_XI0/XI23/XI0/NET35_XI0/XI23/XI0/MM11_g N_VDD_XI0/XI23/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI1/MM2 N_XI0/XI23/XI1/NET34_XI0/XI23/XI1/MM2_d
+ N_XI0/XI23/XI1/NET33_XI0/XI23/XI1/MM2_g N_VSS_XI0/XI23/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM3 N_XI0/XI23/XI1/NET33_XI0/XI23/XI1/MM3_d
+ N_WL<42>_XI0/XI23/XI1/MM3_g N_BLN<14>_XI0/XI23/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM0 N_XI0/XI23/XI1/NET34_XI0/XI23/XI1/MM0_d
+ N_WL<42>_XI0/XI23/XI1/MM0_g N_BL<14>_XI0/XI23/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM1 N_XI0/XI23/XI1/NET33_XI0/XI23/XI1/MM1_d
+ N_XI0/XI23/XI1/NET34_XI0/XI23/XI1/MM1_g N_VSS_XI0/XI23/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM9 N_XI0/XI23/XI1/NET36_XI0/XI23/XI1/MM9_d
+ N_WL<43>_XI0/XI23/XI1/MM9_g N_BL<14>_XI0/XI23/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM6 N_XI0/XI23/XI1/NET35_XI0/XI23/XI1/MM6_d
+ N_XI0/XI23/XI1/NET36_XI0/XI23/XI1/MM6_g N_VSS_XI0/XI23/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM7 N_XI0/XI23/XI1/NET36_XI0/XI23/XI1/MM7_d
+ N_XI0/XI23/XI1/NET35_XI0/XI23/XI1/MM7_g N_VSS_XI0/XI23/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM8 N_XI0/XI23/XI1/NET35_XI0/XI23/XI1/MM8_d
+ N_WL<43>_XI0/XI23/XI1/MM8_g N_BLN<14>_XI0/XI23/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI1/MM5 N_XI0/XI23/XI1/NET34_XI0/XI23/XI1/MM5_d
+ N_XI0/XI23/XI1/NET33_XI0/XI23/XI1/MM5_g N_VDD_XI0/XI23/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI1/MM4 N_XI0/XI23/XI1/NET33_XI0/XI23/XI1/MM4_d
+ N_XI0/XI23/XI1/NET34_XI0/XI23/XI1/MM4_g N_VDD_XI0/XI23/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI1/MM10 N_XI0/XI23/XI1/NET35_XI0/XI23/XI1/MM10_d
+ N_XI0/XI23/XI1/NET36_XI0/XI23/XI1/MM10_g N_VDD_XI0/XI23/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI1/MM11 N_XI0/XI23/XI1/NET36_XI0/XI23/XI1/MM11_d
+ N_XI0/XI23/XI1/NET35_XI0/XI23/XI1/MM11_g N_VDD_XI0/XI23/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI2/MM2 N_XI0/XI23/XI2/NET34_XI0/XI23/XI2/MM2_d
+ N_XI0/XI23/XI2/NET33_XI0/XI23/XI2/MM2_g N_VSS_XI0/XI23/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM3 N_XI0/XI23/XI2/NET33_XI0/XI23/XI2/MM3_d
+ N_WL<42>_XI0/XI23/XI2/MM3_g N_BLN<13>_XI0/XI23/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM0 N_XI0/XI23/XI2/NET34_XI0/XI23/XI2/MM0_d
+ N_WL<42>_XI0/XI23/XI2/MM0_g N_BL<13>_XI0/XI23/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM1 N_XI0/XI23/XI2/NET33_XI0/XI23/XI2/MM1_d
+ N_XI0/XI23/XI2/NET34_XI0/XI23/XI2/MM1_g N_VSS_XI0/XI23/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM9 N_XI0/XI23/XI2/NET36_XI0/XI23/XI2/MM9_d
+ N_WL<43>_XI0/XI23/XI2/MM9_g N_BL<13>_XI0/XI23/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM6 N_XI0/XI23/XI2/NET35_XI0/XI23/XI2/MM6_d
+ N_XI0/XI23/XI2/NET36_XI0/XI23/XI2/MM6_g N_VSS_XI0/XI23/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM7 N_XI0/XI23/XI2/NET36_XI0/XI23/XI2/MM7_d
+ N_XI0/XI23/XI2/NET35_XI0/XI23/XI2/MM7_g N_VSS_XI0/XI23/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM8 N_XI0/XI23/XI2/NET35_XI0/XI23/XI2/MM8_d
+ N_WL<43>_XI0/XI23/XI2/MM8_g N_BLN<13>_XI0/XI23/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI2/MM5 N_XI0/XI23/XI2/NET34_XI0/XI23/XI2/MM5_d
+ N_XI0/XI23/XI2/NET33_XI0/XI23/XI2/MM5_g N_VDD_XI0/XI23/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI2/MM4 N_XI0/XI23/XI2/NET33_XI0/XI23/XI2/MM4_d
+ N_XI0/XI23/XI2/NET34_XI0/XI23/XI2/MM4_g N_VDD_XI0/XI23/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI2/MM10 N_XI0/XI23/XI2/NET35_XI0/XI23/XI2/MM10_d
+ N_XI0/XI23/XI2/NET36_XI0/XI23/XI2/MM10_g N_VDD_XI0/XI23/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI2/MM11 N_XI0/XI23/XI2/NET36_XI0/XI23/XI2/MM11_d
+ N_XI0/XI23/XI2/NET35_XI0/XI23/XI2/MM11_g N_VDD_XI0/XI23/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI3/MM2 N_XI0/XI23/XI3/NET34_XI0/XI23/XI3/MM2_d
+ N_XI0/XI23/XI3/NET33_XI0/XI23/XI3/MM2_g N_VSS_XI0/XI23/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM3 N_XI0/XI23/XI3/NET33_XI0/XI23/XI3/MM3_d
+ N_WL<42>_XI0/XI23/XI3/MM3_g N_BLN<12>_XI0/XI23/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM0 N_XI0/XI23/XI3/NET34_XI0/XI23/XI3/MM0_d
+ N_WL<42>_XI0/XI23/XI3/MM0_g N_BL<12>_XI0/XI23/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM1 N_XI0/XI23/XI3/NET33_XI0/XI23/XI3/MM1_d
+ N_XI0/XI23/XI3/NET34_XI0/XI23/XI3/MM1_g N_VSS_XI0/XI23/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM9 N_XI0/XI23/XI3/NET36_XI0/XI23/XI3/MM9_d
+ N_WL<43>_XI0/XI23/XI3/MM9_g N_BL<12>_XI0/XI23/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM6 N_XI0/XI23/XI3/NET35_XI0/XI23/XI3/MM6_d
+ N_XI0/XI23/XI3/NET36_XI0/XI23/XI3/MM6_g N_VSS_XI0/XI23/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM7 N_XI0/XI23/XI3/NET36_XI0/XI23/XI3/MM7_d
+ N_XI0/XI23/XI3/NET35_XI0/XI23/XI3/MM7_g N_VSS_XI0/XI23/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM8 N_XI0/XI23/XI3/NET35_XI0/XI23/XI3/MM8_d
+ N_WL<43>_XI0/XI23/XI3/MM8_g N_BLN<12>_XI0/XI23/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI3/MM5 N_XI0/XI23/XI3/NET34_XI0/XI23/XI3/MM5_d
+ N_XI0/XI23/XI3/NET33_XI0/XI23/XI3/MM5_g N_VDD_XI0/XI23/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI3/MM4 N_XI0/XI23/XI3/NET33_XI0/XI23/XI3/MM4_d
+ N_XI0/XI23/XI3/NET34_XI0/XI23/XI3/MM4_g N_VDD_XI0/XI23/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI3/MM10 N_XI0/XI23/XI3/NET35_XI0/XI23/XI3/MM10_d
+ N_XI0/XI23/XI3/NET36_XI0/XI23/XI3/MM10_g N_VDD_XI0/XI23/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI3/MM11 N_XI0/XI23/XI3/NET36_XI0/XI23/XI3/MM11_d
+ N_XI0/XI23/XI3/NET35_XI0/XI23/XI3/MM11_g N_VDD_XI0/XI23/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI4/MM2 N_XI0/XI23/XI4/NET34_XI0/XI23/XI4/MM2_d
+ N_XI0/XI23/XI4/NET33_XI0/XI23/XI4/MM2_g N_VSS_XI0/XI23/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM3 N_XI0/XI23/XI4/NET33_XI0/XI23/XI4/MM3_d
+ N_WL<42>_XI0/XI23/XI4/MM3_g N_BLN<11>_XI0/XI23/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM0 N_XI0/XI23/XI4/NET34_XI0/XI23/XI4/MM0_d
+ N_WL<42>_XI0/XI23/XI4/MM0_g N_BL<11>_XI0/XI23/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM1 N_XI0/XI23/XI4/NET33_XI0/XI23/XI4/MM1_d
+ N_XI0/XI23/XI4/NET34_XI0/XI23/XI4/MM1_g N_VSS_XI0/XI23/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM9 N_XI0/XI23/XI4/NET36_XI0/XI23/XI4/MM9_d
+ N_WL<43>_XI0/XI23/XI4/MM9_g N_BL<11>_XI0/XI23/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM6 N_XI0/XI23/XI4/NET35_XI0/XI23/XI4/MM6_d
+ N_XI0/XI23/XI4/NET36_XI0/XI23/XI4/MM6_g N_VSS_XI0/XI23/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM7 N_XI0/XI23/XI4/NET36_XI0/XI23/XI4/MM7_d
+ N_XI0/XI23/XI4/NET35_XI0/XI23/XI4/MM7_g N_VSS_XI0/XI23/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM8 N_XI0/XI23/XI4/NET35_XI0/XI23/XI4/MM8_d
+ N_WL<43>_XI0/XI23/XI4/MM8_g N_BLN<11>_XI0/XI23/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI4/MM5 N_XI0/XI23/XI4/NET34_XI0/XI23/XI4/MM5_d
+ N_XI0/XI23/XI4/NET33_XI0/XI23/XI4/MM5_g N_VDD_XI0/XI23/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI4/MM4 N_XI0/XI23/XI4/NET33_XI0/XI23/XI4/MM4_d
+ N_XI0/XI23/XI4/NET34_XI0/XI23/XI4/MM4_g N_VDD_XI0/XI23/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI4/MM10 N_XI0/XI23/XI4/NET35_XI0/XI23/XI4/MM10_d
+ N_XI0/XI23/XI4/NET36_XI0/XI23/XI4/MM10_g N_VDD_XI0/XI23/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI4/MM11 N_XI0/XI23/XI4/NET36_XI0/XI23/XI4/MM11_d
+ N_XI0/XI23/XI4/NET35_XI0/XI23/XI4/MM11_g N_VDD_XI0/XI23/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI5/MM2 N_XI0/XI23/XI5/NET34_XI0/XI23/XI5/MM2_d
+ N_XI0/XI23/XI5/NET33_XI0/XI23/XI5/MM2_g N_VSS_XI0/XI23/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM3 N_XI0/XI23/XI5/NET33_XI0/XI23/XI5/MM3_d
+ N_WL<42>_XI0/XI23/XI5/MM3_g N_BLN<10>_XI0/XI23/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM0 N_XI0/XI23/XI5/NET34_XI0/XI23/XI5/MM0_d
+ N_WL<42>_XI0/XI23/XI5/MM0_g N_BL<10>_XI0/XI23/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM1 N_XI0/XI23/XI5/NET33_XI0/XI23/XI5/MM1_d
+ N_XI0/XI23/XI5/NET34_XI0/XI23/XI5/MM1_g N_VSS_XI0/XI23/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM9 N_XI0/XI23/XI5/NET36_XI0/XI23/XI5/MM9_d
+ N_WL<43>_XI0/XI23/XI5/MM9_g N_BL<10>_XI0/XI23/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM6 N_XI0/XI23/XI5/NET35_XI0/XI23/XI5/MM6_d
+ N_XI0/XI23/XI5/NET36_XI0/XI23/XI5/MM6_g N_VSS_XI0/XI23/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM7 N_XI0/XI23/XI5/NET36_XI0/XI23/XI5/MM7_d
+ N_XI0/XI23/XI5/NET35_XI0/XI23/XI5/MM7_g N_VSS_XI0/XI23/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM8 N_XI0/XI23/XI5/NET35_XI0/XI23/XI5/MM8_d
+ N_WL<43>_XI0/XI23/XI5/MM8_g N_BLN<10>_XI0/XI23/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI5/MM5 N_XI0/XI23/XI5/NET34_XI0/XI23/XI5/MM5_d
+ N_XI0/XI23/XI5/NET33_XI0/XI23/XI5/MM5_g N_VDD_XI0/XI23/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI5/MM4 N_XI0/XI23/XI5/NET33_XI0/XI23/XI5/MM4_d
+ N_XI0/XI23/XI5/NET34_XI0/XI23/XI5/MM4_g N_VDD_XI0/XI23/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI5/MM10 N_XI0/XI23/XI5/NET35_XI0/XI23/XI5/MM10_d
+ N_XI0/XI23/XI5/NET36_XI0/XI23/XI5/MM10_g N_VDD_XI0/XI23/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI5/MM11 N_XI0/XI23/XI5/NET36_XI0/XI23/XI5/MM11_d
+ N_XI0/XI23/XI5/NET35_XI0/XI23/XI5/MM11_g N_VDD_XI0/XI23/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI6/MM2 N_XI0/XI23/XI6/NET34_XI0/XI23/XI6/MM2_d
+ N_XI0/XI23/XI6/NET33_XI0/XI23/XI6/MM2_g N_VSS_XI0/XI23/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM3 N_XI0/XI23/XI6/NET33_XI0/XI23/XI6/MM3_d
+ N_WL<42>_XI0/XI23/XI6/MM3_g N_BLN<9>_XI0/XI23/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM0 N_XI0/XI23/XI6/NET34_XI0/XI23/XI6/MM0_d
+ N_WL<42>_XI0/XI23/XI6/MM0_g N_BL<9>_XI0/XI23/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM1 N_XI0/XI23/XI6/NET33_XI0/XI23/XI6/MM1_d
+ N_XI0/XI23/XI6/NET34_XI0/XI23/XI6/MM1_g N_VSS_XI0/XI23/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM9 N_XI0/XI23/XI6/NET36_XI0/XI23/XI6/MM9_d
+ N_WL<43>_XI0/XI23/XI6/MM9_g N_BL<9>_XI0/XI23/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM6 N_XI0/XI23/XI6/NET35_XI0/XI23/XI6/MM6_d
+ N_XI0/XI23/XI6/NET36_XI0/XI23/XI6/MM6_g N_VSS_XI0/XI23/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM7 N_XI0/XI23/XI6/NET36_XI0/XI23/XI6/MM7_d
+ N_XI0/XI23/XI6/NET35_XI0/XI23/XI6/MM7_g N_VSS_XI0/XI23/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM8 N_XI0/XI23/XI6/NET35_XI0/XI23/XI6/MM8_d
+ N_WL<43>_XI0/XI23/XI6/MM8_g N_BLN<9>_XI0/XI23/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI6/MM5 N_XI0/XI23/XI6/NET34_XI0/XI23/XI6/MM5_d
+ N_XI0/XI23/XI6/NET33_XI0/XI23/XI6/MM5_g N_VDD_XI0/XI23/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI6/MM4 N_XI0/XI23/XI6/NET33_XI0/XI23/XI6/MM4_d
+ N_XI0/XI23/XI6/NET34_XI0/XI23/XI6/MM4_g N_VDD_XI0/XI23/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI6/MM10 N_XI0/XI23/XI6/NET35_XI0/XI23/XI6/MM10_d
+ N_XI0/XI23/XI6/NET36_XI0/XI23/XI6/MM10_g N_VDD_XI0/XI23/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI6/MM11 N_XI0/XI23/XI6/NET36_XI0/XI23/XI6/MM11_d
+ N_XI0/XI23/XI6/NET35_XI0/XI23/XI6/MM11_g N_VDD_XI0/XI23/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI7/MM2 N_XI0/XI23/XI7/NET34_XI0/XI23/XI7/MM2_d
+ N_XI0/XI23/XI7/NET33_XI0/XI23/XI7/MM2_g N_VSS_XI0/XI23/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM3 N_XI0/XI23/XI7/NET33_XI0/XI23/XI7/MM3_d
+ N_WL<42>_XI0/XI23/XI7/MM3_g N_BLN<8>_XI0/XI23/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM0 N_XI0/XI23/XI7/NET34_XI0/XI23/XI7/MM0_d
+ N_WL<42>_XI0/XI23/XI7/MM0_g N_BL<8>_XI0/XI23/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM1 N_XI0/XI23/XI7/NET33_XI0/XI23/XI7/MM1_d
+ N_XI0/XI23/XI7/NET34_XI0/XI23/XI7/MM1_g N_VSS_XI0/XI23/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM9 N_XI0/XI23/XI7/NET36_XI0/XI23/XI7/MM9_d
+ N_WL<43>_XI0/XI23/XI7/MM9_g N_BL<8>_XI0/XI23/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM6 N_XI0/XI23/XI7/NET35_XI0/XI23/XI7/MM6_d
+ N_XI0/XI23/XI7/NET36_XI0/XI23/XI7/MM6_g N_VSS_XI0/XI23/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM7 N_XI0/XI23/XI7/NET36_XI0/XI23/XI7/MM7_d
+ N_XI0/XI23/XI7/NET35_XI0/XI23/XI7/MM7_g N_VSS_XI0/XI23/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM8 N_XI0/XI23/XI7/NET35_XI0/XI23/XI7/MM8_d
+ N_WL<43>_XI0/XI23/XI7/MM8_g N_BLN<8>_XI0/XI23/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI7/MM5 N_XI0/XI23/XI7/NET34_XI0/XI23/XI7/MM5_d
+ N_XI0/XI23/XI7/NET33_XI0/XI23/XI7/MM5_g N_VDD_XI0/XI23/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI7/MM4 N_XI0/XI23/XI7/NET33_XI0/XI23/XI7/MM4_d
+ N_XI0/XI23/XI7/NET34_XI0/XI23/XI7/MM4_g N_VDD_XI0/XI23/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI7/MM10 N_XI0/XI23/XI7/NET35_XI0/XI23/XI7/MM10_d
+ N_XI0/XI23/XI7/NET36_XI0/XI23/XI7/MM10_g N_VDD_XI0/XI23/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI7/MM11 N_XI0/XI23/XI7/NET36_XI0/XI23/XI7/MM11_d
+ N_XI0/XI23/XI7/NET35_XI0/XI23/XI7/MM11_g N_VDD_XI0/XI23/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI8/MM2 N_XI0/XI23/XI8/NET34_XI0/XI23/XI8/MM2_d
+ N_XI0/XI23/XI8/NET33_XI0/XI23/XI8/MM2_g N_VSS_XI0/XI23/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM3 N_XI0/XI23/XI8/NET33_XI0/XI23/XI8/MM3_d
+ N_WL<42>_XI0/XI23/XI8/MM3_g N_BLN<7>_XI0/XI23/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM0 N_XI0/XI23/XI8/NET34_XI0/XI23/XI8/MM0_d
+ N_WL<42>_XI0/XI23/XI8/MM0_g N_BL<7>_XI0/XI23/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM1 N_XI0/XI23/XI8/NET33_XI0/XI23/XI8/MM1_d
+ N_XI0/XI23/XI8/NET34_XI0/XI23/XI8/MM1_g N_VSS_XI0/XI23/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM9 N_XI0/XI23/XI8/NET36_XI0/XI23/XI8/MM9_d
+ N_WL<43>_XI0/XI23/XI8/MM9_g N_BL<7>_XI0/XI23/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM6 N_XI0/XI23/XI8/NET35_XI0/XI23/XI8/MM6_d
+ N_XI0/XI23/XI8/NET36_XI0/XI23/XI8/MM6_g N_VSS_XI0/XI23/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM7 N_XI0/XI23/XI8/NET36_XI0/XI23/XI8/MM7_d
+ N_XI0/XI23/XI8/NET35_XI0/XI23/XI8/MM7_g N_VSS_XI0/XI23/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM8 N_XI0/XI23/XI8/NET35_XI0/XI23/XI8/MM8_d
+ N_WL<43>_XI0/XI23/XI8/MM8_g N_BLN<7>_XI0/XI23/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI8/MM5 N_XI0/XI23/XI8/NET34_XI0/XI23/XI8/MM5_d
+ N_XI0/XI23/XI8/NET33_XI0/XI23/XI8/MM5_g N_VDD_XI0/XI23/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI8/MM4 N_XI0/XI23/XI8/NET33_XI0/XI23/XI8/MM4_d
+ N_XI0/XI23/XI8/NET34_XI0/XI23/XI8/MM4_g N_VDD_XI0/XI23/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI8/MM10 N_XI0/XI23/XI8/NET35_XI0/XI23/XI8/MM10_d
+ N_XI0/XI23/XI8/NET36_XI0/XI23/XI8/MM10_g N_VDD_XI0/XI23/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI8/MM11 N_XI0/XI23/XI8/NET36_XI0/XI23/XI8/MM11_d
+ N_XI0/XI23/XI8/NET35_XI0/XI23/XI8/MM11_g N_VDD_XI0/XI23/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI9/MM2 N_XI0/XI23/XI9/NET34_XI0/XI23/XI9/MM2_d
+ N_XI0/XI23/XI9/NET33_XI0/XI23/XI9/MM2_g N_VSS_XI0/XI23/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM3 N_XI0/XI23/XI9/NET33_XI0/XI23/XI9/MM3_d
+ N_WL<42>_XI0/XI23/XI9/MM3_g N_BLN<6>_XI0/XI23/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM0 N_XI0/XI23/XI9/NET34_XI0/XI23/XI9/MM0_d
+ N_WL<42>_XI0/XI23/XI9/MM0_g N_BL<6>_XI0/XI23/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM1 N_XI0/XI23/XI9/NET33_XI0/XI23/XI9/MM1_d
+ N_XI0/XI23/XI9/NET34_XI0/XI23/XI9/MM1_g N_VSS_XI0/XI23/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM9 N_XI0/XI23/XI9/NET36_XI0/XI23/XI9/MM9_d
+ N_WL<43>_XI0/XI23/XI9/MM9_g N_BL<6>_XI0/XI23/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM6 N_XI0/XI23/XI9/NET35_XI0/XI23/XI9/MM6_d
+ N_XI0/XI23/XI9/NET36_XI0/XI23/XI9/MM6_g N_VSS_XI0/XI23/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM7 N_XI0/XI23/XI9/NET36_XI0/XI23/XI9/MM7_d
+ N_XI0/XI23/XI9/NET35_XI0/XI23/XI9/MM7_g N_VSS_XI0/XI23/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM8 N_XI0/XI23/XI9/NET35_XI0/XI23/XI9/MM8_d
+ N_WL<43>_XI0/XI23/XI9/MM8_g N_BLN<6>_XI0/XI23/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI9/MM5 N_XI0/XI23/XI9/NET34_XI0/XI23/XI9/MM5_d
+ N_XI0/XI23/XI9/NET33_XI0/XI23/XI9/MM5_g N_VDD_XI0/XI23/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI9/MM4 N_XI0/XI23/XI9/NET33_XI0/XI23/XI9/MM4_d
+ N_XI0/XI23/XI9/NET34_XI0/XI23/XI9/MM4_g N_VDD_XI0/XI23/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI9/MM10 N_XI0/XI23/XI9/NET35_XI0/XI23/XI9/MM10_d
+ N_XI0/XI23/XI9/NET36_XI0/XI23/XI9/MM10_g N_VDD_XI0/XI23/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI9/MM11 N_XI0/XI23/XI9/NET36_XI0/XI23/XI9/MM11_d
+ N_XI0/XI23/XI9/NET35_XI0/XI23/XI9/MM11_g N_VDD_XI0/XI23/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI10/MM2 N_XI0/XI23/XI10/NET34_XI0/XI23/XI10/MM2_d
+ N_XI0/XI23/XI10/NET33_XI0/XI23/XI10/MM2_g N_VSS_XI0/XI23/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM3 N_XI0/XI23/XI10/NET33_XI0/XI23/XI10/MM3_d
+ N_WL<42>_XI0/XI23/XI10/MM3_g N_BLN<5>_XI0/XI23/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM0 N_XI0/XI23/XI10/NET34_XI0/XI23/XI10/MM0_d
+ N_WL<42>_XI0/XI23/XI10/MM0_g N_BL<5>_XI0/XI23/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM1 N_XI0/XI23/XI10/NET33_XI0/XI23/XI10/MM1_d
+ N_XI0/XI23/XI10/NET34_XI0/XI23/XI10/MM1_g N_VSS_XI0/XI23/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM9 N_XI0/XI23/XI10/NET36_XI0/XI23/XI10/MM9_d
+ N_WL<43>_XI0/XI23/XI10/MM9_g N_BL<5>_XI0/XI23/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM6 N_XI0/XI23/XI10/NET35_XI0/XI23/XI10/MM6_d
+ N_XI0/XI23/XI10/NET36_XI0/XI23/XI10/MM6_g N_VSS_XI0/XI23/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM7 N_XI0/XI23/XI10/NET36_XI0/XI23/XI10/MM7_d
+ N_XI0/XI23/XI10/NET35_XI0/XI23/XI10/MM7_g N_VSS_XI0/XI23/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM8 N_XI0/XI23/XI10/NET35_XI0/XI23/XI10/MM8_d
+ N_WL<43>_XI0/XI23/XI10/MM8_g N_BLN<5>_XI0/XI23/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI10/MM5 N_XI0/XI23/XI10/NET34_XI0/XI23/XI10/MM5_d
+ N_XI0/XI23/XI10/NET33_XI0/XI23/XI10/MM5_g N_VDD_XI0/XI23/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI10/MM4 N_XI0/XI23/XI10/NET33_XI0/XI23/XI10/MM4_d
+ N_XI0/XI23/XI10/NET34_XI0/XI23/XI10/MM4_g N_VDD_XI0/XI23/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI10/MM10 N_XI0/XI23/XI10/NET35_XI0/XI23/XI10/MM10_d
+ N_XI0/XI23/XI10/NET36_XI0/XI23/XI10/MM10_g N_VDD_XI0/XI23/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI10/MM11 N_XI0/XI23/XI10/NET36_XI0/XI23/XI10/MM11_d
+ N_XI0/XI23/XI10/NET35_XI0/XI23/XI10/MM11_g N_VDD_XI0/XI23/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI11/MM2 N_XI0/XI23/XI11/NET34_XI0/XI23/XI11/MM2_d
+ N_XI0/XI23/XI11/NET33_XI0/XI23/XI11/MM2_g N_VSS_XI0/XI23/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM3 N_XI0/XI23/XI11/NET33_XI0/XI23/XI11/MM3_d
+ N_WL<42>_XI0/XI23/XI11/MM3_g N_BLN<4>_XI0/XI23/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM0 N_XI0/XI23/XI11/NET34_XI0/XI23/XI11/MM0_d
+ N_WL<42>_XI0/XI23/XI11/MM0_g N_BL<4>_XI0/XI23/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM1 N_XI0/XI23/XI11/NET33_XI0/XI23/XI11/MM1_d
+ N_XI0/XI23/XI11/NET34_XI0/XI23/XI11/MM1_g N_VSS_XI0/XI23/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM9 N_XI0/XI23/XI11/NET36_XI0/XI23/XI11/MM9_d
+ N_WL<43>_XI0/XI23/XI11/MM9_g N_BL<4>_XI0/XI23/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM6 N_XI0/XI23/XI11/NET35_XI0/XI23/XI11/MM6_d
+ N_XI0/XI23/XI11/NET36_XI0/XI23/XI11/MM6_g N_VSS_XI0/XI23/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM7 N_XI0/XI23/XI11/NET36_XI0/XI23/XI11/MM7_d
+ N_XI0/XI23/XI11/NET35_XI0/XI23/XI11/MM7_g N_VSS_XI0/XI23/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM8 N_XI0/XI23/XI11/NET35_XI0/XI23/XI11/MM8_d
+ N_WL<43>_XI0/XI23/XI11/MM8_g N_BLN<4>_XI0/XI23/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI11/MM5 N_XI0/XI23/XI11/NET34_XI0/XI23/XI11/MM5_d
+ N_XI0/XI23/XI11/NET33_XI0/XI23/XI11/MM5_g N_VDD_XI0/XI23/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI11/MM4 N_XI0/XI23/XI11/NET33_XI0/XI23/XI11/MM4_d
+ N_XI0/XI23/XI11/NET34_XI0/XI23/XI11/MM4_g N_VDD_XI0/XI23/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI11/MM10 N_XI0/XI23/XI11/NET35_XI0/XI23/XI11/MM10_d
+ N_XI0/XI23/XI11/NET36_XI0/XI23/XI11/MM10_g N_VDD_XI0/XI23/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI11/MM11 N_XI0/XI23/XI11/NET36_XI0/XI23/XI11/MM11_d
+ N_XI0/XI23/XI11/NET35_XI0/XI23/XI11/MM11_g N_VDD_XI0/XI23/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI12/MM2 N_XI0/XI23/XI12/NET34_XI0/XI23/XI12/MM2_d
+ N_XI0/XI23/XI12/NET33_XI0/XI23/XI12/MM2_g N_VSS_XI0/XI23/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM3 N_XI0/XI23/XI12/NET33_XI0/XI23/XI12/MM3_d
+ N_WL<42>_XI0/XI23/XI12/MM3_g N_BLN<3>_XI0/XI23/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM0 N_XI0/XI23/XI12/NET34_XI0/XI23/XI12/MM0_d
+ N_WL<42>_XI0/XI23/XI12/MM0_g N_BL<3>_XI0/XI23/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM1 N_XI0/XI23/XI12/NET33_XI0/XI23/XI12/MM1_d
+ N_XI0/XI23/XI12/NET34_XI0/XI23/XI12/MM1_g N_VSS_XI0/XI23/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM9 N_XI0/XI23/XI12/NET36_XI0/XI23/XI12/MM9_d
+ N_WL<43>_XI0/XI23/XI12/MM9_g N_BL<3>_XI0/XI23/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM6 N_XI0/XI23/XI12/NET35_XI0/XI23/XI12/MM6_d
+ N_XI0/XI23/XI12/NET36_XI0/XI23/XI12/MM6_g N_VSS_XI0/XI23/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM7 N_XI0/XI23/XI12/NET36_XI0/XI23/XI12/MM7_d
+ N_XI0/XI23/XI12/NET35_XI0/XI23/XI12/MM7_g N_VSS_XI0/XI23/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM8 N_XI0/XI23/XI12/NET35_XI0/XI23/XI12/MM8_d
+ N_WL<43>_XI0/XI23/XI12/MM8_g N_BLN<3>_XI0/XI23/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI12/MM5 N_XI0/XI23/XI12/NET34_XI0/XI23/XI12/MM5_d
+ N_XI0/XI23/XI12/NET33_XI0/XI23/XI12/MM5_g N_VDD_XI0/XI23/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI12/MM4 N_XI0/XI23/XI12/NET33_XI0/XI23/XI12/MM4_d
+ N_XI0/XI23/XI12/NET34_XI0/XI23/XI12/MM4_g N_VDD_XI0/XI23/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI12/MM10 N_XI0/XI23/XI12/NET35_XI0/XI23/XI12/MM10_d
+ N_XI0/XI23/XI12/NET36_XI0/XI23/XI12/MM10_g N_VDD_XI0/XI23/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI12/MM11 N_XI0/XI23/XI12/NET36_XI0/XI23/XI12/MM11_d
+ N_XI0/XI23/XI12/NET35_XI0/XI23/XI12/MM11_g N_VDD_XI0/XI23/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI13/MM2 N_XI0/XI23/XI13/NET34_XI0/XI23/XI13/MM2_d
+ N_XI0/XI23/XI13/NET33_XI0/XI23/XI13/MM2_g N_VSS_XI0/XI23/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM3 N_XI0/XI23/XI13/NET33_XI0/XI23/XI13/MM3_d
+ N_WL<42>_XI0/XI23/XI13/MM3_g N_BLN<2>_XI0/XI23/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM0 N_XI0/XI23/XI13/NET34_XI0/XI23/XI13/MM0_d
+ N_WL<42>_XI0/XI23/XI13/MM0_g N_BL<2>_XI0/XI23/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM1 N_XI0/XI23/XI13/NET33_XI0/XI23/XI13/MM1_d
+ N_XI0/XI23/XI13/NET34_XI0/XI23/XI13/MM1_g N_VSS_XI0/XI23/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM9 N_XI0/XI23/XI13/NET36_XI0/XI23/XI13/MM9_d
+ N_WL<43>_XI0/XI23/XI13/MM9_g N_BL<2>_XI0/XI23/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM6 N_XI0/XI23/XI13/NET35_XI0/XI23/XI13/MM6_d
+ N_XI0/XI23/XI13/NET36_XI0/XI23/XI13/MM6_g N_VSS_XI0/XI23/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM7 N_XI0/XI23/XI13/NET36_XI0/XI23/XI13/MM7_d
+ N_XI0/XI23/XI13/NET35_XI0/XI23/XI13/MM7_g N_VSS_XI0/XI23/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM8 N_XI0/XI23/XI13/NET35_XI0/XI23/XI13/MM8_d
+ N_WL<43>_XI0/XI23/XI13/MM8_g N_BLN<2>_XI0/XI23/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI13/MM5 N_XI0/XI23/XI13/NET34_XI0/XI23/XI13/MM5_d
+ N_XI0/XI23/XI13/NET33_XI0/XI23/XI13/MM5_g N_VDD_XI0/XI23/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI13/MM4 N_XI0/XI23/XI13/NET33_XI0/XI23/XI13/MM4_d
+ N_XI0/XI23/XI13/NET34_XI0/XI23/XI13/MM4_g N_VDD_XI0/XI23/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI13/MM10 N_XI0/XI23/XI13/NET35_XI0/XI23/XI13/MM10_d
+ N_XI0/XI23/XI13/NET36_XI0/XI23/XI13/MM10_g N_VDD_XI0/XI23/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI13/MM11 N_XI0/XI23/XI13/NET36_XI0/XI23/XI13/MM11_d
+ N_XI0/XI23/XI13/NET35_XI0/XI23/XI13/MM11_g N_VDD_XI0/XI23/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI14/MM2 N_XI0/XI23/XI14/NET34_XI0/XI23/XI14/MM2_d
+ N_XI0/XI23/XI14/NET33_XI0/XI23/XI14/MM2_g N_VSS_XI0/XI23/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM3 N_XI0/XI23/XI14/NET33_XI0/XI23/XI14/MM3_d
+ N_WL<42>_XI0/XI23/XI14/MM3_g N_BLN<1>_XI0/XI23/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM0 N_XI0/XI23/XI14/NET34_XI0/XI23/XI14/MM0_d
+ N_WL<42>_XI0/XI23/XI14/MM0_g N_BL<1>_XI0/XI23/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM1 N_XI0/XI23/XI14/NET33_XI0/XI23/XI14/MM1_d
+ N_XI0/XI23/XI14/NET34_XI0/XI23/XI14/MM1_g N_VSS_XI0/XI23/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM9 N_XI0/XI23/XI14/NET36_XI0/XI23/XI14/MM9_d
+ N_WL<43>_XI0/XI23/XI14/MM9_g N_BL<1>_XI0/XI23/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM6 N_XI0/XI23/XI14/NET35_XI0/XI23/XI14/MM6_d
+ N_XI0/XI23/XI14/NET36_XI0/XI23/XI14/MM6_g N_VSS_XI0/XI23/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM7 N_XI0/XI23/XI14/NET36_XI0/XI23/XI14/MM7_d
+ N_XI0/XI23/XI14/NET35_XI0/XI23/XI14/MM7_g N_VSS_XI0/XI23/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM8 N_XI0/XI23/XI14/NET35_XI0/XI23/XI14/MM8_d
+ N_WL<43>_XI0/XI23/XI14/MM8_g N_BLN<1>_XI0/XI23/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI14/MM5 N_XI0/XI23/XI14/NET34_XI0/XI23/XI14/MM5_d
+ N_XI0/XI23/XI14/NET33_XI0/XI23/XI14/MM5_g N_VDD_XI0/XI23/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI14/MM4 N_XI0/XI23/XI14/NET33_XI0/XI23/XI14/MM4_d
+ N_XI0/XI23/XI14/NET34_XI0/XI23/XI14/MM4_g N_VDD_XI0/XI23/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI14/MM10 N_XI0/XI23/XI14/NET35_XI0/XI23/XI14/MM10_d
+ N_XI0/XI23/XI14/NET36_XI0/XI23/XI14/MM10_g N_VDD_XI0/XI23/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI14/MM11 N_XI0/XI23/XI14/NET36_XI0/XI23/XI14/MM11_d
+ N_XI0/XI23/XI14/NET35_XI0/XI23/XI14/MM11_g N_VDD_XI0/XI23/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI15/MM2 N_XI0/XI23/XI15/NET34_XI0/XI23/XI15/MM2_d
+ N_XI0/XI23/XI15/NET33_XI0/XI23/XI15/MM2_g N_VSS_XI0/XI23/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM3 N_XI0/XI23/XI15/NET33_XI0/XI23/XI15/MM3_d
+ N_WL<42>_XI0/XI23/XI15/MM3_g N_BLN<0>_XI0/XI23/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM0 N_XI0/XI23/XI15/NET34_XI0/XI23/XI15/MM0_d
+ N_WL<42>_XI0/XI23/XI15/MM0_g N_BL<0>_XI0/XI23/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM1 N_XI0/XI23/XI15/NET33_XI0/XI23/XI15/MM1_d
+ N_XI0/XI23/XI15/NET34_XI0/XI23/XI15/MM1_g N_VSS_XI0/XI23/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM9 N_XI0/XI23/XI15/NET36_XI0/XI23/XI15/MM9_d
+ N_WL<43>_XI0/XI23/XI15/MM9_g N_BL<0>_XI0/XI23/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM6 N_XI0/XI23/XI15/NET35_XI0/XI23/XI15/MM6_d
+ N_XI0/XI23/XI15/NET36_XI0/XI23/XI15/MM6_g N_VSS_XI0/XI23/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM7 N_XI0/XI23/XI15/NET36_XI0/XI23/XI15/MM7_d
+ N_XI0/XI23/XI15/NET35_XI0/XI23/XI15/MM7_g N_VSS_XI0/XI23/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM8 N_XI0/XI23/XI15/NET35_XI0/XI23/XI15/MM8_d
+ N_WL<43>_XI0/XI23/XI15/MM8_g N_BLN<0>_XI0/XI23/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI23/XI15/MM5 N_XI0/XI23/XI15/NET34_XI0/XI23/XI15/MM5_d
+ N_XI0/XI23/XI15/NET33_XI0/XI23/XI15/MM5_g N_VDD_XI0/XI23/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI15/MM4 N_XI0/XI23/XI15/NET33_XI0/XI23/XI15/MM4_d
+ N_XI0/XI23/XI15/NET34_XI0/XI23/XI15/MM4_g N_VDD_XI0/XI23/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI15/MM10 N_XI0/XI23/XI15/NET35_XI0/XI23/XI15/MM10_d
+ N_XI0/XI23/XI15/NET36_XI0/XI23/XI15/MM10_g N_VDD_XI0/XI23/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI23/XI15/MM11 N_XI0/XI23/XI15/NET36_XI0/XI23/XI15/MM11_d
+ N_XI0/XI23/XI15/NET35_XI0/XI23/XI15/MM11_g N_VDD_XI0/XI23/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI0/MM2 N_XI0/XI24/XI0/NET34_XI0/XI24/XI0/MM2_d
+ N_XI0/XI24/XI0/NET33_XI0/XI24/XI0/MM2_g N_VSS_XI0/XI24/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM3 N_XI0/XI24/XI0/NET33_XI0/XI24/XI0/MM3_d
+ N_WL<44>_XI0/XI24/XI0/MM3_g N_BLN<15>_XI0/XI24/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM0 N_XI0/XI24/XI0/NET34_XI0/XI24/XI0/MM0_d
+ N_WL<44>_XI0/XI24/XI0/MM0_g N_BL<15>_XI0/XI24/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM1 N_XI0/XI24/XI0/NET33_XI0/XI24/XI0/MM1_d
+ N_XI0/XI24/XI0/NET34_XI0/XI24/XI0/MM1_g N_VSS_XI0/XI24/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM9 N_XI0/XI24/XI0/NET36_XI0/XI24/XI0/MM9_d
+ N_WL<45>_XI0/XI24/XI0/MM9_g N_BL<15>_XI0/XI24/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM6 N_XI0/XI24/XI0/NET35_XI0/XI24/XI0/MM6_d
+ N_XI0/XI24/XI0/NET36_XI0/XI24/XI0/MM6_g N_VSS_XI0/XI24/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM7 N_XI0/XI24/XI0/NET36_XI0/XI24/XI0/MM7_d
+ N_XI0/XI24/XI0/NET35_XI0/XI24/XI0/MM7_g N_VSS_XI0/XI24/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM8 N_XI0/XI24/XI0/NET35_XI0/XI24/XI0/MM8_d
+ N_WL<45>_XI0/XI24/XI0/MM8_g N_BLN<15>_XI0/XI24/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI0/MM5 N_XI0/XI24/XI0/NET34_XI0/XI24/XI0/MM5_d
+ N_XI0/XI24/XI0/NET33_XI0/XI24/XI0/MM5_g N_VDD_XI0/XI24/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI0/MM4 N_XI0/XI24/XI0/NET33_XI0/XI24/XI0/MM4_d
+ N_XI0/XI24/XI0/NET34_XI0/XI24/XI0/MM4_g N_VDD_XI0/XI24/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI0/MM10 N_XI0/XI24/XI0/NET35_XI0/XI24/XI0/MM10_d
+ N_XI0/XI24/XI0/NET36_XI0/XI24/XI0/MM10_g N_VDD_XI0/XI24/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI0/MM11 N_XI0/XI24/XI0/NET36_XI0/XI24/XI0/MM11_d
+ N_XI0/XI24/XI0/NET35_XI0/XI24/XI0/MM11_g N_VDD_XI0/XI24/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI1/MM2 N_XI0/XI24/XI1/NET34_XI0/XI24/XI1/MM2_d
+ N_XI0/XI24/XI1/NET33_XI0/XI24/XI1/MM2_g N_VSS_XI0/XI24/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM3 N_XI0/XI24/XI1/NET33_XI0/XI24/XI1/MM3_d
+ N_WL<44>_XI0/XI24/XI1/MM3_g N_BLN<14>_XI0/XI24/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM0 N_XI0/XI24/XI1/NET34_XI0/XI24/XI1/MM0_d
+ N_WL<44>_XI0/XI24/XI1/MM0_g N_BL<14>_XI0/XI24/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM1 N_XI0/XI24/XI1/NET33_XI0/XI24/XI1/MM1_d
+ N_XI0/XI24/XI1/NET34_XI0/XI24/XI1/MM1_g N_VSS_XI0/XI24/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM9 N_XI0/XI24/XI1/NET36_XI0/XI24/XI1/MM9_d
+ N_WL<45>_XI0/XI24/XI1/MM9_g N_BL<14>_XI0/XI24/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM6 N_XI0/XI24/XI1/NET35_XI0/XI24/XI1/MM6_d
+ N_XI0/XI24/XI1/NET36_XI0/XI24/XI1/MM6_g N_VSS_XI0/XI24/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM7 N_XI0/XI24/XI1/NET36_XI0/XI24/XI1/MM7_d
+ N_XI0/XI24/XI1/NET35_XI0/XI24/XI1/MM7_g N_VSS_XI0/XI24/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM8 N_XI0/XI24/XI1/NET35_XI0/XI24/XI1/MM8_d
+ N_WL<45>_XI0/XI24/XI1/MM8_g N_BLN<14>_XI0/XI24/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI1/MM5 N_XI0/XI24/XI1/NET34_XI0/XI24/XI1/MM5_d
+ N_XI0/XI24/XI1/NET33_XI0/XI24/XI1/MM5_g N_VDD_XI0/XI24/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI1/MM4 N_XI0/XI24/XI1/NET33_XI0/XI24/XI1/MM4_d
+ N_XI0/XI24/XI1/NET34_XI0/XI24/XI1/MM4_g N_VDD_XI0/XI24/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI1/MM10 N_XI0/XI24/XI1/NET35_XI0/XI24/XI1/MM10_d
+ N_XI0/XI24/XI1/NET36_XI0/XI24/XI1/MM10_g N_VDD_XI0/XI24/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI1/MM11 N_XI0/XI24/XI1/NET36_XI0/XI24/XI1/MM11_d
+ N_XI0/XI24/XI1/NET35_XI0/XI24/XI1/MM11_g N_VDD_XI0/XI24/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI2/MM2 N_XI0/XI24/XI2/NET34_XI0/XI24/XI2/MM2_d
+ N_XI0/XI24/XI2/NET33_XI0/XI24/XI2/MM2_g N_VSS_XI0/XI24/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM3 N_XI0/XI24/XI2/NET33_XI0/XI24/XI2/MM3_d
+ N_WL<44>_XI0/XI24/XI2/MM3_g N_BLN<13>_XI0/XI24/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM0 N_XI0/XI24/XI2/NET34_XI0/XI24/XI2/MM0_d
+ N_WL<44>_XI0/XI24/XI2/MM0_g N_BL<13>_XI0/XI24/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM1 N_XI0/XI24/XI2/NET33_XI0/XI24/XI2/MM1_d
+ N_XI0/XI24/XI2/NET34_XI0/XI24/XI2/MM1_g N_VSS_XI0/XI24/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM9 N_XI0/XI24/XI2/NET36_XI0/XI24/XI2/MM9_d
+ N_WL<45>_XI0/XI24/XI2/MM9_g N_BL<13>_XI0/XI24/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM6 N_XI0/XI24/XI2/NET35_XI0/XI24/XI2/MM6_d
+ N_XI0/XI24/XI2/NET36_XI0/XI24/XI2/MM6_g N_VSS_XI0/XI24/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM7 N_XI0/XI24/XI2/NET36_XI0/XI24/XI2/MM7_d
+ N_XI0/XI24/XI2/NET35_XI0/XI24/XI2/MM7_g N_VSS_XI0/XI24/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM8 N_XI0/XI24/XI2/NET35_XI0/XI24/XI2/MM8_d
+ N_WL<45>_XI0/XI24/XI2/MM8_g N_BLN<13>_XI0/XI24/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI2/MM5 N_XI0/XI24/XI2/NET34_XI0/XI24/XI2/MM5_d
+ N_XI0/XI24/XI2/NET33_XI0/XI24/XI2/MM5_g N_VDD_XI0/XI24/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI2/MM4 N_XI0/XI24/XI2/NET33_XI0/XI24/XI2/MM4_d
+ N_XI0/XI24/XI2/NET34_XI0/XI24/XI2/MM4_g N_VDD_XI0/XI24/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI2/MM10 N_XI0/XI24/XI2/NET35_XI0/XI24/XI2/MM10_d
+ N_XI0/XI24/XI2/NET36_XI0/XI24/XI2/MM10_g N_VDD_XI0/XI24/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI2/MM11 N_XI0/XI24/XI2/NET36_XI0/XI24/XI2/MM11_d
+ N_XI0/XI24/XI2/NET35_XI0/XI24/XI2/MM11_g N_VDD_XI0/XI24/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI3/MM2 N_XI0/XI24/XI3/NET34_XI0/XI24/XI3/MM2_d
+ N_XI0/XI24/XI3/NET33_XI0/XI24/XI3/MM2_g N_VSS_XI0/XI24/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM3 N_XI0/XI24/XI3/NET33_XI0/XI24/XI3/MM3_d
+ N_WL<44>_XI0/XI24/XI3/MM3_g N_BLN<12>_XI0/XI24/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM0 N_XI0/XI24/XI3/NET34_XI0/XI24/XI3/MM0_d
+ N_WL<44>_XI0/XI24/XI3/MM0_g N_BL<12>_XI0/XI24/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM1 N_XI0/XI24/XI3/NET33_XI0/XI24/XI3/MM1_d
+ N_XI0/XI24/XI3/NET34_XI0/XI24/XI3/MM1_g N_VSS_XI0/XI24/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM9 N_XI0/XI24/XI3/NET36_XI0/XI24/XI3/MM9_d
+ N_WL<45>_XI0/XI24/XI3/MM9_g N_BL<12>_XI0/XI24/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM6 N_XI0/XI24/XI3/NET35_XI0/XI24/XI3/MM6_d
+ N_XI0/XI24/XI3/NET36_XI0/XI24/XI3/MM6_g N_VSS_XI0/XI24/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM7 N_XI0/XI24/XI3/NET36_XI0/XI24/XI3/MM7_d
+ N_XI0/XI24/XI3/NET35_XI0/XI24/XI3/MM7_g N_VSS_XI0/XI24/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM8 N_XI0/XI24/XI3/NET35_XI0/XI24/XI3/MM8_d
+ N_WL<45>_XI0/XI24/XI3/MM8_g N_BLN<12>_XI0/XI24/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI3/MM5 N_XI0/XI24/XI3/NET34_XI0/XI24/XI3/MM5_d
+ N_XI0/XI24/XI3/NET33_XI0/XI24/XI3/MM5_g N_VDD_XI0/XI24/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI3/MM4 N_XI0/XI24/XI3/NET33_XI0/XI24/XI3/MM4_d
+ N_XI0/XI24/XI3/NET34_XI0/XI24/XI3/MM4_g N_VDD_XI0/XI24/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI3/MM10 N_XI0/XI24/XI3/NET35_XI0/XI24/XI3/MM10_d
+ N_XI0/XI24/XI3/NET36_XI0/XI24/XI3/MM10_g N_VDD_XI0/XI24/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI3/MM11 N_XI0/XI24/XI3/NET36_XI0/XI24/XI3/MM11_d
+ N_XI0/XI24/XI3/NET35_XI0/XI24/XI3/MM11_g N_VDD_XI0/XI24/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI4/MM2 N_XI0/XI24/XI4/NET34_XI0/XI24/XI4/MM2_d
+ N_XI0/XI24/XI4/NET33_XI0/XI24/XI4/MM2_g N_VSS_XI0/XI24/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM3 N_XI0/XI24/XI4/NET33_XI0/XI24/XI4/MM3_d
+ N_WL<44>_XI0/XI24/XI4/MM3_g N_BLN<11>_XI0/XI24/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM0 N_XI0/XI24/XI4/NET34_XI0/XI24/XI4/MM0_d
+ N_WL<44>_XI0/XI24/XI4/MM0_g N_BL<11>_XI0/XI24/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM1 N_XI0/XI24/XI4/NET33_XI0/XI24/XI4/MM1_d
+ N_XI0/XI24/XI4/NET34_XI0/XI24/XI4/MM1_g N_VSS_XI0/XI24/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM9 N_XI0/XI24/XI4/NET36_XI0/XI24/XI4/MM9_d
+ N_WL<45>_XI0/XI24/XI4/MM9_g N_BL<11>_XI0/XI24/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM6 N_XI0/XI24/XI4/NET35_XI0/XI24/XI4/MM6_d
+ N_XI0/XI24/XI4/NET36_XI0/XI24/XI4/MM6_g N_VSS_XI0/XI24/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM7 N_XI0/XI24/XI4/NET36_XI0/XI24/XI4/MM7_d
+ N_XI0/XI24/XI4/NET35_XI0/XI24/XI4/MM7_g N_VSS_XI0/XI24/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM8 N_XI0/XI24/XI4/NET35_XI0/XI24/XI4/MM8_d
+ N_WL<45>_XI0/XI24/XI4/MM8_g N_BLN<11>_XI0/XI24/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI4/MM5 N_XI0/XI24/XI4/NET34_XI0/XI24/XI4/MM5_d
+ N_XI0/XI24/XI4/NET33_XI0/XI24/XI4/MM5_g N_VDD_XI0/XI24/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI4/MM4 N_XI0/XI24/XI4/NET33_XI0/XI24/XI4/MM4_d
+ N_XI0/XI24/XI4/NET34_XI0/XI24/XI4/MM4_g N_VDD_XI0/XI24/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI4/MM10 N_XI0/XI24/XI4/NET35_XI0/XI24/XI4/MM10_d
+ N_XI0/XI24/XI4/NET36_XI0/XI24/XI4/MM10_g N_VDD_XI0/XI24/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI4/MM11 N_XI0/XI24/XI4/NET36_XI0/XI24/XI4/MM11_d
+ N_XI0/XI24/XI4/NET35_XI0/XI24/XI4/MM11_g N_VDD_XI0/XI24/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI5/MM2 N_XI0/XI24/XI5/NET34_XI0/XI24/XI5/MM2_d
+ N_XI0/XI24/XI5/NET33_XI0/XI24/XI5/MM2_g N_VSS_XI0/XI24/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM3 N_XI0/XI24/XI5/NET33_XI0/XI24/XI5/MM3_d
+ N_WL<44>_XI0/XI24/XI5/MM3_g N_BLN<10>_XI0/XI24/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM0 N_XI0/XI24/XI5/NET34_XI0/XI24/XI5/MM0_d
+ N_WL<44>_XI0/XI24/XI5/MM0_g N_BL<10>_XI0/XI24/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM1 N_XI0/XI24/XI5/NET33_XI0/XI24/XI5/MM1_d
+ N_XI0/XI24/XI5/NET34_XI0/XI24/XI5/MM1_g N_VSS_XI0/XI24/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM9 N_XI0/XI24/XI5/NET36_XI0/XI24/XI5/MM9_d
+ N_WL<45>_XI0/XI24/XI5/MM9_g N_BL<10>_XI0/XI24/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM6 N_XI0/XI24/XI5/NET35_XI0/XI24/XI5/MM6_d
+ N_XI0/XI24/XI5/NET36_XI0/XI24/XI5/MM6_g N_VSS_XI0/XI24/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM7 N_XI0/XI24/XI5/NET36_XI0/XI24/XI5/MM7_d
+ N_XI0/XI24/XI5/NET35_XI0/XI24/XI5/MM7_g N_VSS_XI0/XI24/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM8 N_XI0/XI24/XI5/NET35_XI0/XI24/XI5/MM8_d
+ N_WL<45>_XI0/XI24/XI5/MM8_g N_BLN<10>_XI0/XI24/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI5/MM5 N_XI0/XI24/XI5/NET34_XI0/XI24/XI5/MM5_d
+ N_XI0/XI24/XI5/NET33_XI0/XI24/XI5/MM5_g N_VDD_XI0/XI24/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI5/MM4 N_XI0/XI24/XI5/NET33_XI0/XI24/XI5/MM4_d
+ N_XI0/XI24/XI5/NET34_XI0/XI24/XI5/MM4_g N_VDD_XI0/XI24/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI5/MM10 N_XI0/XI24/XI5/NET35_XI0/XI24/XI5/MM10_d
+ N_XI0/XI24/XI5/NET36_XI0/XI24/XI5/MM10_g N_VDD_XI0/XI24/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI5/MM11 N_XI0/XI24/XI5/NET36_XI0/XI24/XI5/MM11_d
+ N_XI0/XI24/XI5/NET35_XI0/XI24/XI5/MM11_g N_VDD_XI0/XI24/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI6/MM2 N_XI0/XI24/XI6/NET34_XI0/XI24/XI6/MM2_d
+ N_XI0/XI24/XI6/NET33_XI0/XI24/XI6/MM2_g N_VSS_XI0/XI24/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM3 N_XI0/XI24/XI6/NET33_XI0/XI24/XI6/MM3_d
+ N_WL<44>_XI0/XI24/XI6/MM3_g N_BLN<9>_XI0/XI24/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM0 N_XI0/XI24/XI6/NET34_XI0/XI24/XI6/MM0_d
+ N_WL<44>_XI0/XI24/XI6/MM0_g N_BL<9>_XI0/XI24/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM1 N_XI0/XI24/XI6/NET33_XI0/XI24/XI6/MM1_d
+ N_XI0/XI24/XI6/NET34_XI0/XI24/XI6/MM1_g N_VSS_XI0/XI24/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM9 N_XI0/XI24/XI6/NET36_XI0/XI24/XI6/MM9_d
+ N_WL<45>_XI0/XI24/XI6/MM9_g N_BL<9>_XI0/XI24/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM6 N_XI0/XI24/XI6/NET35_XI0/XI24/XI6/MM6_d
+ N_XI0/XI24/XI6/NET36_XI0/XI24/XI6/MM6_g N_VSS_XI0/XI24/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM7 N_XI0/XI24/XI6/NET36_XI0/XI24/XI6/MM7_d
+ N_XI0/XI24/XI6/NET35_XI0/XI24/XI6/MM7_g N_VSS_XI0/XI24/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM8 N_XI0/XI24/XI6/NET35_XI0/XI24/XI6/MM8_d
+ N_WL<45>_XI0/XI24/XI6/MM8_g N_BLN<9>_XI0/XI24/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI6/MM5 N_XI0/XI24/XI6/NET34_XI0/XI24/XI6/MM5_d
+ N_XI0/XI24/XI6/NET33_XI0/XI24/XI6/MM5_g N_VDD_XI0/XI24/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI6/MM4 N_XI0/XI24/XI6/NET33_XI0/XI24/XI6/MM4_d
+ N_XI0/XI24/XI6/NET34_XI0/XI24/XI6/MM4_g N_VDD_XI0/XI24/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI6/MM10 N_XI0/XI24/XI6/NET35_XI0/XI24/XI6/MM10_d
+ N_XI0/XI24/XI6/NET36_XI0/XI24/XI6/MM10_g N_VDD_XI0/XI24/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI6/MM11 N_XI0/XI24/XI6/NET36_XI0/XI24/XI6/MM11_d
+ N_XI0/XI24/XI6/NET35_XI0/XI24/XI6/MM11_g N_VDD_XI0/XI24/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI7/MM2 N_XI0/XI24/XI7/NET34_XI0/XI24/XI7/MM2_d
+ N_XI0/XI24/XI7/NET33_XI0/XI24/XI7/MM2_g N_VSS_XI0/XI24/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM3 N_XI0/XI24/XI7/NET33_XI0/XI24/XI7/MM3_d
+ N_WL<44>_XI0/XI24/XI7/MM3_g N_BLN<8>_XI0/XI24/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM0 N_XI0/XI24/XI7/NET34_XI0/XI24/XI7/MM0_d
+ N_WL<44>_XI0/XI24/XI7/MM0_g N_BL<8>_XI0/XI24/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM1 N_XI0/XI24/XI7/NET33_XI0/XI24/XI7/MM1_d
+ N_XI0/XI24/XI7/NET34_XI0/XI24/XI7/MM1_g N_VSS_XI0/XI24/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM9 N_XI0/XI24/XI7/NET36_XI0/XI24/XI7/MM9_d
+ N_WL<45>_XI0/XI24/XI7/MM9_g N_BL<8>_XI0/XI24/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM6 N_XI0/XI24/XI7/NET35_XI0/XI24/XI7/MM6_d
+ N_XI0/XI24/XI7/NET36_XI0/XI24/XI7/MM6_g N_VSS_XI0/XI24/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM7 N_XI0/XI24/XI7/NET36_XI0/XI24/XI7/MM7_d
+ N_XI0/XI24/XI7/NET35_XI0/XI24/XI7/MM7_g N_VSS_XI0/XI24/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM8 N_XI0/XI24/XI7/NET35_XI0/XI24/XI7/MM8_d
+ N_WL<45>_XI0/XI24/XI7/MM8_g N_BLN<8>_XI0/XI24/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI7/MM5 N_XI0/XI24/XI7/NET34_XI0/XI24/XI7/MM5_d
+ N_XI0/XI24/XI7/NET33_XI0/XI24/XI7/MM5_g N_VDD_XI0/XI24/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI7/MM4 N_XI0/XI24/XI7/NET33_XI0/XI24/XI7/MM4_d
+ N_XI0/XI24/XI7/NET34_XI0/XI24/XI7/MM4_g N_VDD_XI0/XI24/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI7/MM10 N_XI0/XI24/XI7/NET35_XI0/XI24/XI7/MM10_d
+ N_XI0/XI24/XI7/NET36_XI0/XI24/XI7/MM10_g N_VDD_XI0/XI24/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI7/MM11 N_XI0/XI24/XI7/NET36_XI0/XI24/XI7/MM11_d
+ N_XI0/XI24/XI7/NET35_XI0/XI24/XI7/MM11_g N_VDD_XI0/XI24/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI8/MM2 N_XI0/XI24/XI8/NET34_XI0/XI24/XI8/MM2_d
+ N_XI0/XI24/XI8/NET33_XI0/XI24/XI8/MM2_g N_VSS_XI0/XI24/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM3 N_XI0/XI24/XI8/NET33_XI0/XI24/XI8/MM3_d
+ N_WL<44>_XI0/XI24/XI8/MM3_g N_BLN<7>_XI0/XI24/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM0 N_XI0/XI24/XI8/NET34_XI0/XI24/XI8/MM0_d
+ N_WL<44>_XI0/XI24/XI8/MM0_g N_BL<7>_XI0/XI24/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM1 N_XI0/XI24/XI8/NET33_XI0/XI24/XI8/MM1_d
+ N_XI0/XI24/XI8/NET34_XI0/XI24/XI8/MM1_g N_VSS_XI0/XI24/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM9 N_XI0/XI24/XI8/NET36_XI0/XI24/XI8/MM9_d
+ N_WL<45>_XI0/XI24/XI8/MM9_g N_BL<7>_XI0/XI24/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM6 N_XI0/XI24/XI8/NET35_XI0/XI24/XI8/MM6_d
+ N_XI0/XI24/XI8/NET36_XI0/XI24/XI8/MM6_g N_VSS_XI0/XI24/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM7 N_XI0/XI24/XI8/NET36_XI0/XI24/XI8/MM7_d
+ N_XI0/XI24/XI8/NET35_XI0/XI24/XI8/MM7_g N_VSS_XI0/XI24/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM8 N_XI0/XI24/XI8/NET35_XI0/XI24/XI8/MM8_d
+ N_WL<45>_XI0/XI24/XI8/MM8_g N_BLN<7>_XI0/XI24/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI8/MM5 N_XI0/XI24/XI8/NET34_XI0/XI24/XI8/MM5_d
+ N_XI0/XI24/XI8/NET33_XI0/XI24/XI8/MM5_g N_VDD_XI0/XI24/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI8/MM4 N_XI0/XI24/XI8/NET33_XI0/XI24/XI8/MM4_d
+ N_XI0/XI24/XI8/NET34_XI0/XI24/XI8/MM4_g N_VDD_XI0/XI24/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI8/MM10 N_XI0/XI24/XI8/NET35_XI0/XI24/XI8/MM10_d
+ N_XI0/XI24/XI8/NET36_XI0/XI24/XI8/MM10_g N_VDD_XI0/XI24/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI8/MM11 N_XI0/XI24/XI8/NET36_XI0/XI24/XI8/MM11_d
+ N_XI0/XI24/XI8/NET35_XI0/XI24/XI8/MM11_g N_VDD_XI0/XI24/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI9/MM2 N_XI0/XI24/XI9/NET34_XI0/XI24/XI9/MM2_d
+ N_XI0/XI24/XI9/NET33_XI0/XI24/XI9/MM2_g N_VSS_XI0/XI24/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM3 N_XI0/XI24/XI9/NET33_XI0/XI24/XI9/MM3_d
+ N_WL<44>_XI0/XI24/XI9/MM3_g N_BLN<6>_XI0/XI24/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM0 N_XI0/XI24/XI9/NET34_XI0/XI24/XI9/MM0_d
+ N_WL<44>_XI0/XI24/XI9/MM0_g N_BL<6>_XI0/XI24/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM1 N_XI0/XI24/XI9/NET33_XI0/XI24/XI9/MM1_d
+ N_XI0/XI24/XI9/NET34_XI0/XI24/XI9/MM1_g N_VSS_XI0/XI24/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM9 N_XI0/XI24/XI9/NET36_XI0/XI24/XI9/MM9_d
+ N_WL<45>_XI0/XI24/XI9/MM9_g N_BL<6>_XI0/XI24/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM6 N_XI0/XI24/XI9/NET35_XI0/XI24/XI9/MM6_d
+ N_XI0/XI24/XI9/NET36_XI0/XI24/XI9/MM6_g N_VSS_XI0/XI24/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM7 N_XI0/XI24/XI9/NET36_XI0/XI24/XI9/MM7_d
+ N_XI0/XI24/XI9/NET35_XI0/XI24/XI9/MM7_g N_VSS_XI0/XI24/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM8 N_XI0/XI24/XI9/NET35_XI0/XI24/XI9/MM8_d
+ N_WL<45>_XI0/XI24/XI9/MM8_g N_BLN<6>_XI0/XI24/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI9/MM5 N_XI0/XI24/XI9/NET34_XI0/XI24/XI9/MM5_d
+ N_XI0/XI24/XI9/NET33_XI0/XI24/XI9/MM5_g N_VDD_XI0/XI24/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI9/MM4 N_XI0/XI24/XI9/NET33_XI0/XI24/XI9/MM4_d
+ N_XI0/XI24/XI9/NET34_XI0/XI24/XI9/MM4_g N_VDD_XI0/XI24/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI9/MM10 N_XI0/XI24/XI9/NET35_XI0/XI24/XI9/MM10_d
+ N_XI0/XI24/XI9/NET36_XI0/XI24/XI9/MM10_g N_VDD_XI0/XI24/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI9/MM11 N_XI0/XI24/XI9/NET36_XI0/XI24/XI9/MM11_d
+ N_XI0/XI24/XI9/NET35_XI0/XI24/XI9/MM11_g N_VDD_XI0/XI24/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI10/MM2 N_XI0/XI24/XI10/NET34_XI0/XI24/XI10/MM2_d
+ N_XI0/XI24/XI10/NET33_XI0/XI24/XI10/MM2_g N_VSS_XI0/XI24/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM3 N_XI0/XI24/XI10/NET33_XI0/XI24/XI10/MM3_d
+ N_WL<44>_XI0/XI24/XI10/MM3_g N_BLN<5>_XI0/XI24/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM0 N_XI0/XI24/XI10/NET34_XI0/XI24/XI10/MM0_d
+ N_WL<44>_XI0/XI24/XI10/MM0_g N_BL<5>_XI0/XI24/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM1 N_XI0/XI24/XI10/NET33_XI0/XI24/XI10/MM1_d
+ N_XI0/XI24/XI10/NET34_XI0/XI24/XI10/MM1_g N_VSS_XI0/XI24/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM9 N_XI0/XI24/XI10/NET36_XI0/XI24/XI10/MM9_d
+ N_WL<45>_XI0/XI24/XI10/MM9_g N_BL<5>_XI0/XI24/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM6 N_XI0/XI24/XI10/NET35_XI0/XI24/XI10/MM6_d
+ N_XI0/XI24/XI10/NET36_XI0/XI24/XI10/MM6_g N_VSS_XI0/XI24/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM7 N_XI0/XI24/XI10/NET36_XI0/XI24/XI10/MM7_d
+ N_XI0/XI24/XI10/NET35_XI0/XI24/XI10/MM7_g N_VSS_XI0/XI24/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM8 N_XI0/XI24/XI10/NET35_XI0/XI24/XI10/MM8_d
+ N_WL<45>_XI0/XI24/XI10/MM8_g N_BLN<5>_XI0/XI24/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI10/MM5 N_XI0/XI24/XI10/NET34_XI0/XI24/XI10/MM5_d
+ N_XI0/XI24/XI10/NET33_XI0/XI24/XI10/MM5_g N_VDD_XI0/XI24/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI10/MM4 N_XI0/XI24/XI10/NET33_XI0/XI24/XI10/MM4_d
+ N_XI0/XI24/XI10/NET34_XI0/XI24/XI10/MM4_g N_VDD_XI0/XI24/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI10/MM10 N_XI0/XI24/XI10/NET35_XI0/XI24/XI10/MM10_d
+ N_XI0/XI24/XI10/NET36_XI0/XI24/XI10/MM10_g N_VDD_XI0/XI24/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI10/MM11 N_XI0/XI24/XI10/NET36_XI0/XI24/XI10/MM11_d
+ N_XI0/XI24/XI10/NET35_XI0/XI24/XI10/MM11_g N_VDD_XI0/XI24/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI11/MM2 N_XI0/XI24/XI11/NET34_XI0/XI24/XI11/MM2_d
+ N_XI0/XI24/XI11/NET33_XI0/XI24/XI11/MM2_g N_VSS_XI0/XI24/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM3 N_XI0/XI24/XI11/NET33_XI0/XI24/XI11/MM3_d
+ N_WL<44>_XI0/XI24/XI11/MM3_g N_BLN<4>_XI0/XI24/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM0 N_XI0/XI24/XI11/NET34_XI0/XI24/XI11/MM0_d
+ N_WL<44>_XI0/XI24/XI11/MM0_g N_BL<4>_XI0/XI24/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM1 N_XI0/XI24/XI11/NET33_XI0/XI24/XI11/MM1_d
+ N_XI0/XI24/XI11/NET34_XI0/XI24/XI11/MM1_g N_VSS_XI0/XI24/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM9 N_XI0/XI24/XI11/NET36_XI0/XI24/XI11/MM9_d
+ N_WL<45>_XI0/XI24/XI11/MM9_g N_BL<4>_XI0/XI24/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM6 N_XI0/XI24/XI11/NET35_XI0/XI24/XI11/MM6_d
+ N_XI0/XI24/XI11/NET36_XI0/XI24/XI11/MM6_g N_VSS_XI0/XI24/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM7 N_XI0/XI24/XI11/NET36_XI0/XI24/XI11/MM7_d
+ N_XI0/XI24/XI11/NET35_XI0/XI24/XI11/MM7_g N_VSS_XI0/XI24/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM8 N_XI0/XI24/XI11/NET35_XI0/XI24/XI11/MM8_d
+ N_WL<45>_XI0/XI24/XI11/MM8_g N_BLN<4>_XI0/XI24/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI11/MM5 N_XI0/XI24/XI11/NET34_XI0/XI24/XI11/MM5_d
+ N_XI0/XI24/XI11/NET33_XI0/XI24/XI11/MM5_g N_VDD_XI0/XI24/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI11/MM4 N_XI0/XI24/XI11/NET33_XI0/XI24/XI11/MM4_d
+ N_XI0/XI24/XI11/NET34_XI0/XI24/XI11/MM4_g N_VDD_XI0/XI24/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI11/MM10 N_XI0/XI24/XI11/NET35_XI0/XI24/XI11/MM10_d
+ N_XI0/XI24/XI11/NET36_XI0/XI24/XI11/MM10_g N_VDD_XI0/XI24/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI11/MM11 N_XI0/XI24/XI11/NET36_XI0/XI24/XI11/MM11_d
+ N_XI0/XI24/XI11/NET35_XI0/XI24/XI11/MM11_g N_VDD_XI0/XI24/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI12/MM2 N_XI0/XI24/XI12/NET34_XI0/XI24/XI12/MM2_d
+ N_XI0/XI24/XI12/NET33_XI0/XI24/XI12/MM2_g N_VSS_XI0/XI24/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM3 N_XI0/XI24/XI12/NET33_XI0/XI24/XI12/MM3_d
+ N_WL<44>_XI0/XI24/XI12/MM3_g N_BLN<3>_XI0/XI24/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM0 N_XI0/XI24/XI12/NET34_XI0/XI24/XI12/MM0_d
+ N_WL<44>_XI0/XI24/XI12/MM0_g N_BL<3>_XI0/XI24/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM1 N_XI0/XI24/XI12/NET33_XI0/XI24/XI12/MM1_d
+ N_XI0/XI24/XI12/NET34_XI0/XI24/XI12/MM1_g N_VSS_XI0/XI24/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM9 N_XI0/XI24/XI12/NET36_XI0/XI24/XI12/MM9_d
+ N_WL<45>_XI0/XI24/XI12/MM9_g N_BL<3>_XI0/XI24/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM6 N_XI0/XI24/XI12/NET35_XI0/XI24/XI12/MM6_d
+ N_XI0/XI24/XI12/NET36_XI0/XI24/XI12/MM6_g N_VSS_XI0/XI24/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM7 N_XI0/XI24/XI12/NET36_XI0/XI24/XI12/MM7_d
+ N_XI0/XI24/XI12/NET35_XI0/XI24/XI12/MM7_g N_VSS_XI0/XI24/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM8 N_XI0/XI24/XI12/NET35_XI0/XI24/XI12/MM8_d
+ N_WL<45>_XI0/XI24/XI12/MM8_g N_BLN<3>_XI0/XI24/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI12/MM5 N_XI0/XI24/XI12/NET34_XI0/XI24/XI12/MM5_d
+ N_XI0/XI24/XI12/NET33_XI0/XI24/XI12/MM5_g N_VDD_XI0/XI24/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI12/MM4 N_XI0/XI24/XI12/NET33_XI0/XI24/XI12/MM4_d
+ N_XI0/XI24/XI12/NET34_XI0/XI24/XI12/MM4_g N_VDD_XI0/XI24/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI12/MM10 N_XI0/XI24/XI12/NET35_XI0/XI24/XI12/MM10_d
+ N_XI0/XI24/XI12/NET36_XI0/XI24/XI12/MM10_g N_VDD_XI0/XI24/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI12/MM11 N_XI0/XI24/XI12/NET36_XI0/XI24/XI12/MM11_d
+ N_XI0/XI24/XI12/NET35_XI0/XI24/XI12/MM11_g N_VDD_XI0/XI24/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI13/MM2 N_XI0/XI24/XI13/NET34_XI0/XI24/XI13/MM2_d
+ N_XI0/XI24/XI13/NET33_XI0/XI24/XI13/MM2_g N_VSS_XI0/XI24/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM3 N_XI0/XI24/XI13/NET33_XI0/XI24/XI13/MM3_d
+ N_WL<44>_XI0/XI24/XI13/MM3_g N_BLN<2>_XI0/XI24/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM0 N_XI0/XI24/XI13/NET34_XI0/XI24/XI13/MM0_d
+ N_WL<44>_XI0/XI24/XI13/MM0_g N_BL<2>_XI0/XI24/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM1 N_XI0/XI24/XI13/NET33_XI0/XI24/XI13/MM1_d
+ N_XI0/XI24/XI13/NET34_XI0/XI24/XI13/MM1_g N_VSS_XI0/XI24/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM9 N_XI0/XI24/XI13/NET36_XI0/XI24/XI13/MM9_d
+ N_WL<45>_XI0/XI24/XI13/MM9_g N_BL<2>_XI0/XI24/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM6 N_XI0/XI24/XI13/NET35_XI0/XI24/XI13/MM6_d
+ N_XI0/XI24/XI13/NET36_XI0/XI24/XI13/MM6_g N_VSS_XI0/XI24/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM7 N_XI0/XI24/XI13/NET36_XI0/XI24/XI13/MM7_d
+ N_XI0/XI24/XI13/NET35_XI0/XI24/XI13/MM7_g N_VSS_XI0/XI24/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM8 N_XI0/XI24/XI13/NET35_XI0/XI24/XI13/MM8_d
+ N_WL<45>_XI0/XI24/XI13/MM8_g N_BLN<2>_XI0/XI24/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI13/MM5 N_XI0/XI24/XI13/NET34_XI0/XI24/XI13/MM5_d
+ N_XI0/XI24/XI13/NET33_XI0/XI24/XI13/MM5_g N_VDD_XI0/XI24/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI13/MM4 N_XI0/XI24/XI13/NET33_XI0/XI24/XI13/MM4_d
+ N_XI0/XI24/XI13/NET34_XI0/XI24/XI13/MM4_g N_VDD_XI0/XI24/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI13/MM10 N_XI0/XI24/XI13/NET35_XI0/XI24/XI13/MM10_d
+ N_XI0/XI24/XI13/NET36_XI0/XI24/XI13/MM10_g N_VDD_XI0/XI24/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI13/MM11 N_XI0/XI24/XI13/NET36_XI0/XI24/XI13/MM11_d
+ N_XI0/XI24/XI13/NET35_XI0/XI24/XI13/MM11_g N_VDD_XI0/XI24/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI14/MM2 N_XI0/XI24/XI14/NET34_XI0/XI24/XI14/MM2_d
+ N_XI0/XI24/XI14/NET33_XI0/XI24/XI14/MM2_g N_VSS_XI0/XI24/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM3 N_XI0/XI24/XI14/NET33_XI0/XI24/XI14/MM3_d
+ N_WL<44>_XI0/XI24/XI14/MM3_g N_BLN<1>_XI0/XI24/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM0 N_XI0/XI24/XI14/NET34_XI0/XI24/XI14/MM0_d
+ N_WL<44>_XI0/XI24/XI14/MM0_g N_BL<1>_XI0/XI24/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM1 N_XI0/XI24/XI14/NET33_XI0/XI24/XI14/MM1_d
+ N_XI0/XI24/XI14/NET34_XI0/XI24/XI14/MM1_g N_VSS_XI0/XI24/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM9 N_XI0/XI24/XI14/NET36_XI0/XI24/XI14/MM9_d
+ N_WL<45>_XI0/XI24/XI14/MM9_g N_BL<1>_XI0/XI24/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM6 N_XI0/XI24/XI14/NET35_XI0/XI24/XI14/MM6_d
+ N_XI0/XI24/XI14/NET36_XI0/XI24/XI14/MM6_g N_VSS_XI0/XI24/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM7 N_XI0/XI24/XI14/NET36_XI0/XI24/XI14/MM7_d
+ N_XI0/XI24/XI14/NET35_XI0/XI24/XI14/MM7_g N_VSS_XI0/XI24/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM8 N_XI0/XI24/XI14/NET35_XI0/XI24/XI14/MM8_d
+ N_WL<45>_XI0/XI24/XI14/MM8_g N_BLN<1>_XI0/XI24/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI14/MM5 N_XI0/XI24/XI14/NET34_XI0/XI24/XI14/MM5_d
+ N_XI0/XI24/XI14/NET33_XI0/XI24/XI14/MM5_g N_VDD_XI0/XI24/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI14/MM4 N_XI0/XI24/XI14/NET33_XI0/XI24/XI14/MM4_d
+ N_XI0/XI24/XI14/NET34_XI0/XI24/XI14/MM4_g N_VDD_XI0/XI24/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI14/MM10 N_XI0/XI24/XI14/NET35_XI0/XI24/XI14/MM10_d
+ N_XI0/XI24/XI14/NET36_XI0/XI24/XI14/MM10_g N_VDD_XI0/XI24/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI14/MM11 N_XI0/XI24/XI14/NET36_XI0/XI24/XI14/MM11_d
+ N_XI0/XI24/XI14/NET35_XI0/XI24/XI14/MM11_g N_VDD_XI0/XI24/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI15/MM2 N_XI0/XI24/XI15/NET34_XI0/XI24/XI15/MM2_d
+ N_XI0/XI24/XI15/NET33_XI0/XI24/XI15/MM2_g N_VSS_XI0/XI24/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM3 N_XI0/XI24/XI15/NET33_XI0/XI24/XI15/MM3_d
+ N_WL<44>_XI0/XI24/XI15/MM3_g N_BLN<0>_XI0/XI24/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM0 N_XI0/XI24/XI15/NET34_XI0/XI24/XI15/MM0_d
+ N_WL<44>_XI0/XI24/XI15/MM0_g N_BL<0>_XI0/XI24/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM1 N_XI0/XI24/XI15/NET33_XI0/XI24/XI15/MM1_d
+ N_XI0/XI24/XI15/NET34_XI0/XI24/XI15/MM1_g N_VSS_XI0/XI24/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM9 N_XI0/XI24/XI15/NET36_XI0/XI24/XI15/MM9_d
+ N_WL<45>_XI0/XI24/XI15/MM9_g N_BL<0>_XI0/XI24/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM6 N_XI0/XI24/XI15/NET35_XI0/XI24/XI15/MM6_d
+ N_XI0/XI24/XI15/NET36_XI0/XI24/XI15/MM6_g N_VSS_XI0/XI24/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM7 N_XI0/XI24/XI15/NET36_XI0/XI24/XI15/MM7_d
+ N_XI0/XI24/XI15/NET35_XI0/XI24/XI15/MM7_g N_VSS_XI0/XI24/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM8 N_XI0/XI24/XI15/NET35_XI0/XI24/XI15/MM8_d
+ N_WL<45>_XI0/XI24/XI15/MM8_g N_BLN<0>_XI0/XI24/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI24/XI15/MM5 N_XI0/XI24/XI15/NET34_XI0/XI24/XI15/MM5_d
+ N_XI0/XI24/XI15/NET33_XI0/XI24/XI15/MM5_g N_VDD_XI0/XI24/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI15/MM4 N_XI0/XI24/XI15/NET33_XI0/XI24/XI15/MM4_d
+ N_XI0/XI24/XI15/NET34_XI0/XI24/XI15/MM4_g N_VDD_XI0/XI24/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI15/MM10 N_XI0/XI24/XI15/NET35_XI0/XI24/XI15/MM10_d
+ N_XI0/XI24/XI15/NET36_XI0/XI24/XI15/MM10_g N_VDD_XI0/XI24/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI24/XI15/MM11 N_XI0/XI24/XI15/NET36_XI0/XI24/XI15/MM11_d
+ N_XI0/XI24/XI15/NET35_XI0/XI24/XI15/MM11_g N_VDD_XI0/XI24/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI0/MM2 N_XI0/XI25/XI0/NET34_XI0/XI25/XI0/MM2_d
+ N_XI0/XI25/XI0/NET33_XI0/XI25/XI0/MM2_g N_VSS_XI0/XI25/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM3 N_XI0/XI25/XI0/NET33_XI0/XI25/XI0/MM3_d
+ N_WL<46>_XI0/XI25/XI0/MM3_g N_BLN<15>_XI0/XI25/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM0 N_XI0/XI25/XI0/NET34_XI0/XI25/XI0/MM0_d
+ N_WL<46>_XI0/XI25/XI0/MM0_g N_BL<15>_XI0/XI25/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM1 N_XI0/XI25/XI0/NET33_XI0/XI25/XI0/MM1_d
+ N_XI0/XI25/XI0/NET34_XI0/XI25/XI0/MM1_g N_VSS_XI0/XI25/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM9 N_XI0/XI25/XI0/NET36_XI0/XI25/XI0/MM9_d
+ N_WL<47>_XI0/XI25/XI0/MM9_g N_BL<15>_XI0/XI25/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM6 N_XI0/XI25/XI0/NET35_XI0/XI25/XI0/MM6_d
+ N_XI0/XI25/XI0/NET36_XI0/XI25/XI0/MM6_g N_VSS_XI0/XI25/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM7 N_XI0/XI25/XI0/NET36_XI0/XI25/XI0/MM7_d
+ N_XI0/XI25/XI0/NET35_XI0/XI25/XI0/MM7_g N_VSS_XI0/XI25/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM8 N_XI0/XI25/XI0/NET35_XI0/XI25/XI0/MM8_d
+ N_WL<47>_XI0/XI25/XI0/MM8_g N_BLN<15>_XI0/XI25/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI0/MM5 N_XI0/XI25/XI0/NET34_XI0/XI25/XI0/MM5_d
+ N_XI0/XI25/XI0/NET33_XI0/XI25/XI0/MM5_g N_VDD_XI0/XI25/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI0/MM4 N_XI0/XI25/XI0/NET33_XI0/XI25/XI0/MM4_d
+ N_XI0/XI25/XI0/NET34_XI0/XI25/XI0/MM4_g N_VDD_XI0/XI25/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI0/MM10 N_XI0/XI25/XI0/NET35_XI0/XI25/XI0/MM10_d
+ N_XI0/XI25/XI0/NET36_XI0/XI25/XI0/MM10_g N_VDD_XI0/XI25/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI0/MM11 N_XI0/XI25/XI0/NET36_XI0/XI25/XI0/MM11_d
+ N_XI0/XI25/XI0/NET35_XI0/XI25/XI0/MM11_g N_VDD_XI0/XI25/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI1/MM2 N_XI0/XI25/XI1/NET34_XI0/XI25/XI1/MM2_d
+ N_XI0/XI25/XI1/NET33_XI0/XI25/XI1/MM2_g N_VSS_XI0/XI25/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM3 N_XI0/XI25/XI1/NET33_XI0/XI25/XI1/MM3_d
+ N_WL<46>_XI0/XI25/XI1/MM3_g N_BLN<14>_XI0/XI25/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM0 N_XI0/XI25/XI1/NET34_XI0/XI25/XI1/MM0_d
+ N_WL<46>_XI0/XI25/XI1/MM0_g N_BL<14>_XI0/XI25/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM1 N_XI0/XI25/XI1/NET33_XI0/XI25/XI1/MM1_d
+ N_XI0/XI25/XI1/NET34_XI0/XI25/XI1/MM1_g N_VSS_XI0/XI25/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM9 N_XI0/XI25/XI1/NET36_XI0/XI25/XI1/MM9_d
+ N_WL<47>_XI0/XI25/XI1/MM9_g N_BL<14>_XI0/XI25/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM6 N_XI0/XI25/XI1/NET35_XI0/XI25/XI1/MM6_d
+ N_XI0/XI25/XI1/NET36_XI0/XI25/XI1/MM6_g N_VSS_XI0/XI25/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM7 N_XI0/XI25/XI1/NET36_XI0/XI25/XI1/MM7_d
+ N_XI0/XI25/XI1/NET35_XI0/XI25/XI1/MM7_g N_VSS_XI0/XI25/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM8 N_XI0/XI25/XI1/NET35_XI0/XI25/XI1/MM8_d
+ N_WL<47>_XI0/XI25/XI1/MM8_g N_BLN<14>_XI0/XI25/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI1/MM5 N_XI0/XI25/XI1/NET34_XI0/XI25/XI1/MM5_d
+ N_XI0/XI25/XI1/NET33_XI0/XI25/XI1/MM5_g N_VDD_XI0/XI25/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI1/MM4 N_XI0/XI25/XI1/NET33_XI0/XI25/XI1/MM4_d
+ N_XI0/XI25/XI1/NET34_XI0/XI25/XI1/MM4_g N_VDD_XI0/XI25/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI1/MM10 N_XI0/XI25/XI1/NET35_XI0/XI25/XI1/MM10_d
+ N_XI0/XI25/XI1/NET36_XI0/XI25/XI1/MM10_g N_VDD_XI0/XI25/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI1/MM11 N_XI0/XI25/XI1/NET36_XI0/XI25/XI1/MM11_d
+ N_XI0/XI25/XI1/NET35_XI0/XI25/XI1/MM11_g N_VDD_XI0/XI25/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI2/MM2 N_XI0/XI25/XI2/NET34_XI0/XI25/XI2/MM2_d
+ N_XI0/XI25/XI2/NET33_XI0/XI25/XI2/MM2_g N_VSS_XI0/XI25/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM3 N_XI0/XI25/XI2/NET33_XI0/XI25/XI2/MM3_d
+ N_WL<46>_XI0/XI25/XI2/MM3_g N_BLN<13>_XI0/XI25/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM0 N_XI0/XI25/XI2/NET34_XI0/XI25/XI2/MM0_d
+ N_WL<46>_XI0/XI25/XI2/MM0_g N_BL<13>_XI0/XI25/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM1 N_XI0/XI25/XI2/NET33_XI0/XI25/XI2/MM1_d
+ N_XI0/XI25/XI2/NET34_XI0/XI25/XI2/MM1_g N_VSS_XI0/XI25/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM9 N_XI0/XI25/XI2/NET36_XI0/XI25/XI2/MM9_d
+ N_WL<47>_XI0/XI25/XI2/MM9_g N_BL<13>_XI0/XI25/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM6 N_XI0/XI25/XI2/NET35_XI0/XI25/XI2/MM6_d
+ N_XI0/XI25/XI2/NET36_XI0/XI25/XI2/MM6_g N_VSS_XI0/XI25/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM7 N_XI0/XI25/XI2/NET36_XI0/XI25/XI2/MM7_d
+ N_XI0/XI25/XI2/NET35_XI0/XI25/XI2/MM7_g N_VSS_XI0/XI25/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM8 N_XI0/XI25/XI2/NET35_XI0/XI25/XI2/MM8_d
+ N_WL<47>_XI0/XI25/XI2/MM8_g N_BLN<13>_XI0/XI25/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI2/MM5 N_XI0/XI25/XI2/NET34_XI0/XI25/XI2/MM5_d
+ N_XI0/XI25/XI2/NET33_XI0/XI25/XI2/MM5_g N_VDD_XI0/XI25/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI2/MM4 N_XI0/XI25/XI2/NET33_XI0/XI25/XI2/MM4_d
+ N_XI0/XI25/XI2/NET34_XI0/XI25/XI2/MM4_g N_VDD_XI0/XI25/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI2/MM10 N_XI0/XI25/XI2/NET35_XI0/XI25/XI2/MM10_d
+ N_XI0/XI25/XI2/NET36_XI0/XI25/XI2/MM10_g N_VDD_XI0/XI25/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI2/MM11 N_XI0/XI25/XI2/NET36_XI0/XI25/XI2/MM11_d
+ N_XI0/XI25/XI2/NET35_XI0/XI25/XI2/MM11_g N_VDD_XI0/XI25/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI3/MM2 N_XI0/XI25/XI3/NET34_XI0/XI25/XI3/MM2_d
+ N_XI0/XI25/XI3/NET33_XI0/XI25/XI3/MM2_g N_VSS_XI0/XI25/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM3 N_XI0/XI25/XI3/NET33_XI0/XI25/XI3/MM3_d
+ N_WL<46>_XI0/XI25/XI3/MM3_g N_BLN<12>_XI0/XI25/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM0 N_XI0/XI25/XI3/NET34_XI0/XI25/XI3/MM0_d
+ N_WL<46>_XI0/XI25/XI3/MM0_g N_BL<12>_XI0/XI25/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM1 N_XI0/XI25/XI3/NET33_XI0/XI25/XI3/MM1_d
+ N_XI0/XI25/XI3/NET34_XI0/XI25/XI3/MM1_g N_VSS_XI0/XI25/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM9 N_XI0/XI25/XI3/NET36_XI0/XI25/XI3/MM9_d
+ N_WL<47>_XI0/XI25/XI3/MM9_g N_BL<12>_XI0/XI25/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM6 N_XI0/XI25/XI3/NET35_XI0/XI25/XI3/MM6_d
+ N_XI0/XI25/XI3/NET36_XI0/XI25/XI3/MM6_g N_VSS_XI0/XI25/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM7 N_XI0/XI25/XI3/NET36_XI0/XI25/XI3/MM7_d
+ N_XI0/XI25/XI3/NET35_XI0/XI25/XI3/MM7_g N_VSS_XI0/XI25/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM8 N_XI0/XI25/XI3/NET35_XI0/XI25/XI3/MM8_d
+ N_WL<47>_XI0/XI25/XI3/MM8_g N_BLN<12>_XI0/XI25/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI3/MM5 N_XI0/XI25/XI3/NET34_XI0/XI25/XI3/MM5_d
+ N_XI0/XI25/XI3/NET33_XI0/XI25/XI3/MM5_g N_VDD_XI0/XI25/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI3/MM4 N_XI0/XI25/XI3/NET33_XI0/XI25/XI3/MM4_d
+ N_XI0/XI25/XI3/NET34_XI0/XI25/XI3/MM4_g N_VDD_XI0/XI25/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI3/MM10 N_XI0/XI25/XI3/NET35_XI0/XI25/XI3/MM10_d
+ N_XI0/XI25/XI3/NET36_XI0/XI25/XI3/MM10_g N_VDD_XI0/XI25/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI3/MM11 N_XI0/XI25/XI3/NET36_XI0/XI25/XI3/MM11_d
+ N_XI0/XI25/XI3/NET35_XI0/XI25/XI3/MM11_g N_VDD_XI0/XI25/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI4/MM2 N_XI0/XI25/XI4/NET34_XI0/XI25/XI4/MM2_d
+ N_XI0/XI25/XI4/NET33_XI0/XI25/XI4/MM2_g N_VSS_XI0/XI25/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM3 N_XI0/XI25/XI4/NET33_XI0/XI25/XI4/MM3_d
+ N_WL<46>_XI0/XI25/XI4/MM3_g N_BLN<11>_XI0/XI25/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM0 N_XI0/XI25/XI4/NET34_XI0/XI25/XI4/MM0_d
+ N_WL<46>_XI0/XI25/XI4/MM0_g N_BL<11>_XI0/XI25/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM1 N_XI0/XI25/XI4/NET33_XI0/XI25/XI4/MM1_d
+ N_XI0/XI25/XI4/NET34_XI0/XI25/XI4/MM1_g N_VSS_XI0/XI25/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM9 N_XI0/XI25/XI4/NET36_XI0/XI25/XI4/MM9_d
+ N_WL<47>_XI0/XI25/XI4/MM9_g N_BL<11>_XI0/XI25/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM6 N_XI0/XI25/XI4/NET35_XI0/XI25/XI4/MM6_d
+ N_XI0/XI25/XI4/NET36_XI0/XI25/XI4/MM6_g N_VSS_XI0/XI25/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM7 N_XI0/XI25/XI4/NET36_XI0/XI25/XI4/MM7_d
+ N_XI0/XI25/XI4/NET35_XI0/XI25/XI4/MM7_g N_VSS_XI0/XI25/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM8 N_XI0/XI25/XI4/NET35_XI0/XI25/XI4/MM8_d
+ N_WL<47>_XI0/XI25/XI4/MM8_g N_BLN<11>_XI0/XI25/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI4/MM5 N_XI0/XI25/XI4/NET34_XI0/XI25/XI4/MM5_d
+ N_XI0/XI25/XI4/NET33_XI0/XI25/XI4/MM5_g N_VDD_XI0/XI25/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI4/MM4 N_XI0/XI25/XI4/NET33_XI0/XI25/XI4/MM4_d
+ N_XI0/XI25/XI4/NET34_XI0/XI25/XI4/MM4_g N_VDD_XI0/XI25/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI4/MM10 N_XI0/XI25/XI4/NET35_XI0/XI25/XI4/MM10_d
+ N_XI0/XI25/XI4/NET36_XI0/XI25/XI4/MM10_g N_VDD_XI0/XI25/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI4/MM11 N_XI0/XI25/XI4/NET36_XI0/XI25/XI4/MM11_d
+ N_XI0/XI25/XI4/NET35_XI0/XI25/XI4/MM11_g N_VDD_XI0/XI25/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI5/MM2 N_XI0/XI25/XI5/NET34_XI0/XI25/XI5/MM2_d
+ N_XI0/XI25/XI5/NET33_XI0/XI25/XI5/MM2_g N_VSS_XI0/XI25/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM3 N_XI0/XI25/XI5/NET33_XI0/XI25/XI5/MM3_d
+ N_WL<46>_XI0/XI25/XI5/MM3_g N_BLN<10>_XI0/XI25/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM0 N_XI0/XI25/XI5/NET34_XI0/XI25/XI5/MM0_d
+ N_WL<46>_XI0/XI25/XI5/MM0_g N_BL<10>_XI0/XI25/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM1 N_XI0/XI25/XI5/NET33_XI0/XI25/XI5/MM1_d
+ N_XI0/XI25/XI5/NET34_XI0/XI25/XI5/MM1_g N_VSS_XI0/XI25/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM9 N_XI0/XI25/XI5/NET36_XI0/XI25/XI5/MM9_d
+ N_WL<47>_XI0/XI25/XI5/MM9_g N_BL<10>_XI0/XI25/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM6 N_XI0/XI25/XI5/NET35_XI0/XI25/XI5/MM6_d
+ N_XI0/XI25/XI5/NET36_XI0/XI25/XI5/MM6_g N_VSS_XI0/XI25/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM7 N_XI0/XI25/XI5/NET36_XI0/XI25/XI5/MM7_d
+ N_XI0/XI25/XI5/NET35_XI0/XI25/XI5/MM7_g N_VSS_XI0/XI25/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM8 N_XI0/XI25/XI5/NET35_XI0/XI25/XI5/MM8_d
+ N_WL<47>_XI0/XI25/XI5/MM8_g N_BLN<10>_XI0/XI25/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI5/MM5 N_XI0/XI25/XI5/NET34_XI0/XI25/XI5/MM5_d
+ N_XI0/XI25/XI5/NET33_XI0/XI25/XI5/MM5_g N_VDD_XI0/XI25/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI5/MM4 N_XI0/XI25/XI5/NET33_XI0/XI25/XI5/MM4_d
+ N_XI0/XI25/XI5/NET34_XI0/XI25/XI5/MM4_g N_VDD_XI0/XI25/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI5/MM10 N_XI0/XI25/XI5/NET35_XI0/XI25/XI5/MM10_d
+ N_XI0/XI25/XI5/NET36_XI0/XI25/XI5/MM10_g N_VDD_XI0/XI25/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI5/MM11 N_XI0/XI25/XI5/NET36_XI0/XI25/XI5/MM11_d
+ N_XI0/XI25/XI5/NET35_XI0/XI25/XI5/MM11_g N_VDD_XI0/XI25/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI6/MM2 N_XI0/XI25/XI6/NET34_XI0/XI25/XI6/MM2_d
+ N_XI0/XI25/XI6/NET33_XI0/XI25/XI6/MM2_g N_VSS_XI0/XI25/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM3 N_XI0/XI25/XI6/NET33_XI0/XI25/XI6/MM3_d
+ N_WL<46>_XI0/XI25/XI6/MM3_g N_BLN<9>_XI0/XI25/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM0 N_XI0/XI25/XI6/NET34_XI0/XI25/XI6/MM0_d
+ N_WL<46>_XI0/XI25/XI6/MM0_g N_BL<9>_XI0/XI25/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM1 N_XI0/XI25/XI6/NET33_XI0/XI25/XI6/MM1_d
+ N_XI0/XI25/XI6/NET34_XI0/XI25/XI6/MM1_g N_VSS_XI0/XI25/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM9 N_XI0/XI25/XI6/NET36_XI0/XI25/XI6/MM9_d
+ N_WL<47>_XI0/XI25/XI6/MM9_g N_BL<9>_XI0/XI25/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM6 N_XI0/XI25/XI6/NET35_XI0/XI25/XI6/MM6_d
+ N_XI0/XI25/XI6/NET36_XI0/XI25/XI6/MM6_g N_VSS_XI0/XI25/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM7 N_XI0/XI25/XI6/NET36_XI0/XI25/XI6/MM7_d
+ N_XI0/XI25/XI6/NET35_XI0/XI25/XI6/MM7_g N_VSS_XI0/XI25/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM8 N_XI0/XI25/XI6/NET35_XI0/XI25/XI6/MM8_d
+ N_WL<47>_XI0/XI25/XI6/MM8_g N_BLN<9>_XI0/XI25/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI6/MM5 N_XI0/XI25/XI6/NET34_XI0/XI25/XI6/MM5_d
+ N_XI0/XI25/XI6/NET33_XI0/XI25/XI6/MM5_g N_VDD_XI0/XI25/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI6/MM4 N_XI0/XI25/XI6/NET33_XI0/XI25/XI6/MM4_d
+ N_XI0/XI25/XI6/NET34_XI0/XI25/XI6/MM4_g N_VDD_XI0/XI25/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI6/MM10 N_XI0/XI25/XI6/NET35_XI0/XI25/XI6/MM10_d
+ N_XI0/XI25/XI6/NET36_XI0/XI25/XI6/MM10_g N_VDD_XI0/XI25/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI6/MM11 N_XI0/XI25/XI6/NET36_XI0/XI25/XI6/MM11_d
+ N_XI0/XI25/XI6/NET35_XI0/XI25/XI6/MM11_g N_VDD_XI0/XI25/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI7/MM2 N_XI0/XI25/XI7/NET34_XI0/XI25/XI7/MM2_d
+ N_XI0/XI25/XI7/NET33_XI0/XI25/XI7/MM2_g N_VSS_XI0/XI25/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM3 N_XI0/XI25/XI7/NET33_XI0/XI25/XI7/MM3_d
+ N_WL<46>_XI0/XI25/XI7/MM3_g N_BLN<8>_XI0/XI25/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM0 N_XI0/XI25/XI7/NET34_XI0/XI25/XI7/MM0_d
+ N_WL<46>_XI0/XI25/XI7/MM0_g N_BL<8>_XI0/XI25/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM1 N_XI0/XI25/XI7/NET33_XI0/XI25/XI7/MM1_d
+ N_XI0/XI25/XI7/NET34_XI0/XI25/XI7/MM1_g N_VSS_XI0/XI25/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM9 N_XI0/XI25/XI7/NET36_XI0/XI25/XI7/MM9_d
+ N_WL<47>_XI0/XI25/XI7/MM9_g N_BL<8>_XI0/XI25/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM6 N_XI0/XI25/XI7/NET35_XI0/XI25/XI7/MM6_d
+ N_XI0/XI25/XI7/NET36_XI0/XI25/XI7/MM6_g N_VSS_XI0/XI25/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM7 N_XI0/XI25/XI7/NET36_XI0/XI25/XI7/MM7_d
+ N_XI0/XI25/XI7/NET35_XI0/XI25/XI7/MM7_g N_VSS_XI0/XI25/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM8 N_XI0/XI25/XI7/NET35_XI0/XI25/XI7/MM8_d
+ N_WL<47>_XI0/XI25/XI7/MM8_g N_BLN<8>_XI0/XI25/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI7/MM5 N_XI0/XI25/XI7/NET34_XI0/XI25/XI7/MM5_d
+ N_XI0/XI25/XI7/NET33_XI0/XI25/XI7/MM5_g N_VDD_XI0/XI25/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI7/MM4 N_XI0/XI25/XI7/NET33_XI0/XI25/XI7/MM4_d
+ N_XI0/XI25/XI7/NET34_XI0/XI25/XI7/MM4_g N_VDD_XI0/XI25/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI7/MM10 N_XI0/XI25/XI7/NET35_XI0/XI25/XI7/MM10_d
+ N_XI0/XI25/XI7/NET36_XI0/XI25/XI7/MM10_g N_VDD_XI0/XI25/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI7/MM11 N_XI0/XI25/XI7/NET36_XI0/XI25/XI7/MM11_d
+ N_XI0/XI25/XI7/NET35_XI0/XI25/XI7/MM11_g N_VDD_XI0/XI25/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI8/MM2 N_XI0/XI25/XI8/NET34_XI0/XI25/XI8/MM2_d
+ N_XI0/XI25/XI8/NET33_XI0/XI25/XI8/MM2_g N_VSS_XI0/XI25/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM3 N_XI0/XI25/XI8/NET33_XI0/XI25/XI8/MM3_d
+ N_WL<46>_XI0/XI25/XI8/MM3_g N_BLN<7>_XI0/XI25/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM0 N_XI0/XI25/XI8/NET34_XI0/XI25/XI8/MM0_d
+ N_WL<46>_XI0/XI25/XI8/MM0_g N_BL<7>_XI0/XI25/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM1 N_XI0/XI25/XI8/NET33_XI0/XI25/XI8/MM1_d
+ N_XI0/XI25/XI8/NET34_XI0/XI25/XI8/MM1_g N_VSS_XI0/XI25/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM9 N_XI0/XI25/XI8/NET36_XI0/XI25/XI8/MM9_d
+ N_WL<47>_XI0/XI25/XI8/MM9_g N_BL<7>_XI0/XI25/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM6 N_XI0/XI25/XI8/NET35_XI0/XI25/XI8/MM6_d
+ N_XI0/XI25/XI8/NET36_XI0/XI25/XI8/MM6_g N_VSS_XI0/XI25/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM7 N_XI0/XI25/XI8/NET36_XI0/XI25/XI8/MM7_d
+ N_XI0/XI25/XI8/NET35_XI0/XI25/XI8/MM7_g N_VSS_XI0/XI25/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM8 N_XI0/XI25/XI8/NET35_XI0/XI25/XI8/MM8_d
+ N_WL<47>_XI0/XI25/XI8/MM8_g N_BLN<7>_XI0/XI25/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI8/MM5 N_XI0/XI25/XI8/NET34_XI0/XI25/XI8/MM5_d
+ N_XI0/XI25/XI8/NET33_XI0/XI25/XI8/MM5_g N_VDD_XI0/XI25/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI8/MM4 N_XI0/XI25/XI8/NET33_XI0/XI25/XI8/MM4_d
+ N_XI0/XI25/XI8/NET34_XI0/XI25/XI8/MM4_g N_VDD_XI0/XI25/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI8/MM10 N_XI0/XI25/XI8/NET35_XI0/XI25/XI8/MM10_d
+ N_XI0/XI25/XI8/NET36_XI0/XI25/XI8/MM10_g N_VDD_XI0/XI25/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI8/MM11 N_XI0/XI25/XI8/NET36_XI0/XI25/XI8/MM11_d
+ N_XI0/XI25/XI8/NET35_XI0/XI25/XI8/MM11_g N_VDD_XI0/XI25/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI9/MM2 N_XI0/XI25/XI9/NET34_XI0/XI25/XI9/MM2_d
+ N_XI0/XI25/XI9/NET33_XI0/XI25/XI9/MM2_g N_VSS_XI0/XI25/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM3 N_XI0/XI25/XI9/NET33_XI0/XI25/XI9/MM3_d
+ N_WL<46>_XI0/XI25/XI9/MM3_g N_BLN<6>_XI0/XI25/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM0 N_XI0/XI25/XI9/NET34_XI0/XI25/XI9/MM0_d
+ N_WL<46>_XI0/XI25/XI9/MM0_g N_BL<6>_XI0/XI25/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM1 N_XI0/XI25/XI9/NET33_XI0/XI25/XI9/MM1_d
+ N_XI0/XI25/XI9/NET34_XI0/XI25/XI9/MM1_g N_VSS_XI0/XI25/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM9 N_XI0/XI25/XI9/NET36_XI0/XI25/XI9/MM9_d
+ N_WL<47>_XI0/XI25/XI9/MM9_g N_BL<6>_XI0/XI25/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM6 N_XI0/XI25/XI9/NET35_XI0/XI25/XI9/MM6_d
+ N_XI0/XI25/XI9/NET36_XI0/XI25/XI9/MM6_g N_VSS_XI0/XI25/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM7 N_XI0/XI25/XI9/NET36_XI0/XI25/XI9/MM7_d
+ N_XI0/XI25/XI9/NET35_XI0/XI25/XI9/MM7_g N_VSS_XI0/XI25/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM8 N_XI0/XI25/XI9/NET35_XI0/XI25/XI9/MM8_d
+ N_WL<47>_XI0/XI25/XI9/MM8_g N_BLN<6>_XI0/XI25/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI9/MM5 N_XI0/XI25/XI9/NET34_XI0/XI25/XI9/MM5_d
+ N_XI0/XI25/XI9/NET33_XI0/XI25/XI9/MM5_g N_VDD_XI0/XI25/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI9/MM4 N_XI0/XI25/XI9/NET33_XI0/XI25/XI9/MM4_d
+ N_XI0/XI25/XI9/NET34_XI0/XI25/XI9/MM4_g N_VDD_XI0/XI25/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI9/MM10 N_XI0/XI25/XI9/NET35_XI0/XI25/XI9/MM10_d
+ N_XI0/XI25/XI9/NET36_XI0/XI25/XI9/MM10_g N_VDD_XI0/XI25/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI9/MM11 N_XI0/XI25/XI9/NET36_XI0/XI25/XI9/MM11_d
+ N_XI0/XI25/XI9/NET35_XI0/XI25/XI9/MM11_g N_VDD_XI0/XI25/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI10/MM2 N_XI0/XI25/XI10/NET34_XI0/XI25/XI10/MM2_d
+ N_XI0/XI25/XI10/NET33_XI0/XI25/XI10/MM2_g N_VSS_XI0/XI25/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM3 N_XI0/XI25/XI10/NET33_XI0/XI25/XI10/MM3_d
+ N_WL<46>_XI0/XI25/XI10/MM3_g N_BLN<5>_XI0/XI25/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM0 N_XI0/XI25/XI10/NET34_XI0/XI25/XI10/MM0_d
+ N_WL<46>_XI0/XI25/XI10/MM0_g N_BL<5>_XI0/XI25/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM1 N_XI0/XI25/XI10/NET33_XI0/XI25/XI10/MM1_d
+ N_XI0/XI25/XI10/NET34_XI0/XI25/XI10/MM1_g N_VSS_XI0/XI25/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM9 N_XI0/XI25/XI10/NET36_XI0/XI25/XI10/MM9_d
+ N_WL<47>_XI0/XI25/XI10/MM9_g N_BL<5>_XI0/XI25/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM6 N_XI0/XI25/XI10/NET35_XI0/XI25/XI10/MM6_d
+ N_XI0/XI25/XI10/NET36_XI0/XI25/XI10/MM6_g N_VSS_XI0/XI25/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM7 N_XI0/XI25/XI10/NET36_XI0/XI25/XI10/MM7_d
+ N_XI0/XI25/XI10/NET35_XI0/XI25/XI10/MM7_g N_VSS_XI0/XI25/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM8 N_XI0/XI25/XI10/NET35_XI0/XI25/XI10/MM8_d
+ N_WL<47>_XI0/XI25/XI10/MM8_g N_BLN<5>_XI0/XI25/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI10/MM5 N_XI0/XI25/XI10/NET34_XI0/XI25/XI10/MM5_d
+ N_XI0/XI25/XI10/NET33_XI0/XI25/XI10/MM5_g N_VDD_XI0/XI25/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI10/MM4 N_XI0/XI25/XI10/NET33_XI0/XI25/XI10/MM4_d
+ N_XI0/XI25/XI10/NET34_XI0/XI25/XI10/MM4_g N_VDD_XI0/XI25/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI10/MM10 N_XI0/XI25/XI10/NET35_XI0/XI25/XI10/MM10_d
+ N_XI0/XI25/XI10/NET36_XI0/XI25/XI10/MM10_g N_VDD_XI0/XI25/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI10/MM11 N_XI0/XI25/XI10/NET36_XI0/XI25/XI10/MM11_d
+ N_XI0/XI25/XI10/NET35_XI0/XI25/XI10/MM11_g N_VDD_XI0/XI25/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI11/MM2 N_XI0/XI25/XI11/NET34_XI0/XI25/XI11/MM2_d
+ N_XI0/XI25/XI11/NET33_XI0/XI25/XI11/MM2_g N_VSS_XI0/XI25/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM3 N_XI0/XI25/XI11/NET33_XI0/XI25/XI11/MM3_d
+ N_WL<46>_XI0/XI25/XI11/MM3_g N_BLN<4>_XI0/XI25/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM0 N_XI0/XI25/XI11/NET34_XI0/XI25/XI11/MM0_d
+ N_WL<46>_XI0/XI25/XI11/MM0_g N_BL<4>_XI0/XI25/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM1 N_XI0/XI25/XI11/NET33_XI0/XI25/XI11/MM1_d
+ N_XI0/XI25/XI11/NET34_XI0/XI25/XI11/MM1_g N_VSS_XI0/XI25/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM9 N_XI0/XI25/XI11/NET36_XI0/XI25/XI11/MM9_d
+ N_WL<47>_XI0/XI25/XI11/MM9_g N_BL<4>_XI0/XI25/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM6 N_XI0/XI25/XI11/NET35_XI0/XI25/XI11/MM6_d
+ N_XI0/XI25/XI11/NET36_XI0/XI25/XI11/MM6_g N_VSS_XI0/XI25/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM7 N_XI0/XI25/XI11/NET36_XI0/XI25/XI11/MM7_d
+ N_XI0/XI25/XI11/NET35_XI0/XI25/XI11/MM7_g N_VSS_XI0/XI25/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM8 N_XI0/XI25/XI11/NET35_XI0/XI25/XI11/MM8_d
+ N_WL<47>_XI0/XI25/XI11/MM8_g N_BLN<4>_XI0/XI25/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI11/MM5 N_XI0/XI25/XI11/NET34_XI0/XI25/XI11/MM5_d
+ N_XI0/XI25/XI11/NET33_XI0/XI25/XI11/MM5_g N_VDD_XI0/XI25/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI11/MM4 N_XI0/XI25/XI11/NET33_XI0/XI25/XI11/MM4_d
+ N_XI0/XI25/XI11/NET34_XI0/XI25/XI11/MM4_g N_VDD_XI0/XI25/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI11/MM10 N_XI0/XI25/XI11/NET35_XI0/XI25/XI11/MM10_d
+ N_XI0/XI25/XI11/NET36_XI0/XI25/XI11/MM10_g N_VDD_XI0/XI25/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI11/MM11 N_XI0/XI25/XI11/NET36_XI0/XI25/XI11/MM11_d
+ N_XI0/XI25/XI11/NET35_XI0/XI25/XI11/MM11_g N_VDD_XI0/XI25/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI12/MM2 N_XI0/XI25/XI12/NET34_XI0/XI25/XI12/MM2_d
+ N_XI0/XI25/XI12/NET33_XI0/XI25/XI12/MM2_g N_VSS_XI0/XI25/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM3 N_XI0/XI25/XI12/NET33_XI0/XI25/XI12/MM3_d
+ N_WL<46>_XI0/XI25/XI12/MM3_g N_BLN<3>_XI0/XI25/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM0 N_XI0/XI25/XI12/NET34_XI0/XI25/XI12/MM0_d
+ N_WL<46>_XI0/XI25/XI12/MM0_g N_BL<3>_XI0/XI25/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM1 N_XI0/XI25/XI12/NET33_XI0/XI25/XI12/MM1_d
+ N_XI0/XI25/XI12/NET34_XI0/XI25/XI12/MM1_g N_VSS_XI0/XI25/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM9 N_XI0/XI25/XI12/NET36_XI0/XI25/XI12/MM9_d
+ N_WL<47>_XI0/XI25/XI12/MM9_g N_BL<3>_XI0/XI25/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM6 N_XI0/XI25/XI12/NET35_XI0/XI25/XI12/MM6_d
+ N_XI0/XI25/XI12/NET36_XI0/XI25/XI12/MM6_g N_VSS_XI0/XI25/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM7 N_XI0/XI25/XI12/NET36_XI0/XI25/XI12/MM7_d
+ N_XI0/XI25/XI12/NET35_XI0/XI25/XI12/MM7_g N_VSS_XI0/XI25/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM8 N_XI0/XI25/XI12/NET35_XI0/XI25/XI12/MM8_d
+ N_WL<47>_XI0/XI25/XI12/MM8_g N_BLN<3>_XI0/XI25/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI12/MM5 N_XI0/XI25/XI12/NET34_XI0/XI25/XI12/MM5_d
+ N_XI0/XI25/XI12/NET33_XI0/XI25/XI12/MM5_g N_VDD_XI0/XI25/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI12/MM4 N_XI0/XI25/XI12/NET33_XI0/XI25/XI12/MM4_d
+ N_XI0/XI25/XI12/NET34_XI0/XI25/XI12/MM4_g N_VDD_XI0/XI25/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI12/MM10 N_XI0/XI25/XI12/NET35_XI0/XI25/XI12/MM10_d
+ N_XI0/XI25/XI12/NET36_XI0/XI25/XI12/MM10_g N_VDD_XI0/XI25/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI12/MM11 N_XI0/XI25/XI12/NET36_XI0/XI25/XI12/MM11_d
+ N_XI0/XI25/XI12/NET35_XI0/XI25/XI12/MM11_g N_VDD_XI0/XI25/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI13/MM2 N_XI0/XI25/XI13/NET34_XI0/XI25/XI13/MM2_d
+ N_XI0/XI25/XI13/NET33_XI0/XI25/XI13/MM2_g N_VSS_XI0/XI25/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM3 N_XI0/XI25/XI13/NET33_XI0/XI25/XI13/MM3_d
+ N_WL<46>_XI0/XI25/XI13/MM3_g N_BLN<2>_XI0/XI25/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM0 N_XI0/XI25/XI13/NET34_XI0/XI25/XI13/MM0_d
+ N_WL<46>_XI0/XI25/XI13/MM0_g N_BL<2>_XI0/XI25/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM1 N_XI0/XI25/XI13/NET33_XI0/XI25/XI13/MM1_d
+ N_XI0/XI25/XI13/NET34_XI0/XI25/XI13/MM1_g N_VSS_XI0/XI25/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM9 N_XI0/XI25/XI13/NET36_XI0/XI25/XI13/MM9_d
+ N_WL<47>_XI0/XI25/XI13/MM9_g N_BL<2>_XI0/XI25/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM6 N_XI0/XI25/XI13/NET35_XI0/XI25/XI13/MM6_d
+ N_XI0/XI25/XI13/NET36_XI0/XI25/XI13/MM6_g N_VSS_XI0/XI25/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM7 N_XI0/XI25/XI13/NET36_XI0/XI25/XI13/MM7_d
+ N_XI0/XI25/XI13/NET35_XI0/XI25/XI13/MM7_g N_VSS_XI0/XI25/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM8 N_XI0/XI25/XI13/NET35_XI0/XI25/XI13/MM8_d
+ N_WL<47>_XI0/XI25/XI13/MM8_g N_BLN<2>_XI0/XI25/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI13/MM5 N_XI0/XI25/XI13/NET34_XI0/XI25/XI13/MM5_d
+ N_XI0/XI25/XI13/NET33_XI0/XI25/XI13/MM5_g N_VDD_XI0/XI25/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI13/MM4 N_XI0/XI25/XI13/NET33_XI0/XI25/XI13/MM4_d
+ N_XI0/XI25/XI13/NET34_XI0/XI25/XI13/MM4_g N_VDD_XI0/XI25/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI13/MM10 N_XI0/XI25/XI13/NET35_XI0/XI25/XI13/MM10_d
+ N_XI0/XI25/XI13/NET36_XI0/XI25/XI13/MM10_g N_VDD_XI0/XI25/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI13/MM11 N_XI0/XI25/XI13/NET36_XI0/XI25/XI13/MM11_d
+ N_XI0/XI25/XI13/NET35_XI0/XI25/XI13/MM11_g N_VDD_XI0/XI25/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI14/MM2 N_XI0/XI25/XI14/NET34_XI0/XI25/XI14/MM2_d
+ N_XI0/XI25/XI14/NET33_XI0/XI25/XI14/MM2_g N_VSS_XI0/XI25/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM3 N_XI0/XI25/XI14/NET33_XI0/XI25/XI14/MM3_d
+ N_WL<46>_XI0/XI25/XI14/MM3_g N_BLN<1>_XI0/XI25/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM0 N_XI0/XI25/XI14/NET34_XI0/XI25/XI14/MM0_d
+ N_WL<46>_XI0/XI25/XI14/MM0_g N_BL<1>_XI0/XI25/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM1 N_XI0/XI25/XI14/NET33_XI0/XI25/XI14/MM1_d
+ N_XI0/XI25/XI14/NET34_XI0/XI25/XI14/MM1_g N_VSS_XI0/XI25/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM9 N_XI0/XI25/XI14/NET36_XI0/XI25/XI14/MM9_d
+ N_WL<47>_XI0/XI25/XI14/MM9_g N_BL<1>_XI0/XI25/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM6 N_XI0/XI25/XI14/NET35_XI0/XI25/XI14/MM6_d
+ N_XI0/XI25/XI14/NET36_XI0/XI25/XI14/MM6_g N_VSS_XI0/XI25/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM7 N_XI0/XI25/XI14/NET36_XI0/XI25/XI14/MM7_d
+ N_XI0/XI25/XI14/NET35_XI0/XI25/XI14/MM7_g N_VSS_XI0/XI25/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM8 N_XI0/XI25/XI14/NET35_XI0/XI25/XI14/MM8_d
+ N_WL<47>_XI0/XI25/XI14/MM8_g N_BLN<1>_XI0/XI25/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI14/MM5 N_XI0/XI25/XI14/NET34_XI0/XI25/XI14/MM5_d
+ N_XI0/XI25/XI14/NET33_XI0/XI25/XI14/MM5_g N_VDD_XI0/XI25/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI14/MM4 N_XI0/XI25/XI14/NET33_XI0/XI25/XI14/MM4_d
+ N_XI0/XI25/XI14/NET34_XI0/XI25/XI14/MM4_g N_VDD_XI0/XI25/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI14/MM10 N_XI0/XI25/XI14/NET35_XI0/XI25/XI14/MM10_d
+ N_XI0/XI25/XI14/NET36_XI0/XI25/XI14/MM10_g N_VDD_XI0/XI25/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI14/MM11 N_XI0/XI25/XI14/NET36_XI0/XI25/XI14/MM11_d
+ N_XI0/XI25/XI14/NET35_XI0/XI25/XI14/MM11_g N_VDD_XI0/XI25/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI15/MM2 N_XI0/XI25/XI15/NET34_XI0/XI25/XI15/MM2_d
+ N_XI0/XI25/XI15/NET33_XI0/XI25/XI15/MM2_g N_VSS_XI0/XI25/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM3 N_XI0/XI25/XI15/NET33_XI0/XI25/XI15/MM3_d
+ N_WL<46>_XI0/XI25/XI15/MM3_g N_BLN<0>_XI0/XI25/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM0 N_XI0/XI25/XI15/NET34_XI0/XI25/XI15/MM0_d
+ N_WL<46>_XI0/XI25/XI15/MM0_g N_BL<0>_XI0/XI25/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM1 N_XI0/XI25/XI15/NET33_XI0/XI25/XI15/MM1_d
+ N_XI0/XI25/XI15/NET34_XI0/XI25/XI15/MM1_g N_VSS_XI0/XI25/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM9 N_XI0/XI25/XI15/NET36_XI0/XI25/XI15/MM9_d
+ N_WL<47>_XI0/XI25/XI15/MM9_g N_BL<0>_XI0/XI25/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM6 N_XI0/XI25/XI15/NET35_XI0/XI25/XI15/MM6_d
+ N_XI0/XI25/XI15/NET36_XI0/XI25/XI15/MM6_g N_VSS_XI0/XI25/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM7 N_XI0/XI25/XI15/NET36_XI0/XI25/XI15/MM7_d
+ N_XI0/XI25/XI15/NET35_XI0/XI25/XI15/MM7_g N_VSS_XI0/XI25/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM8 N_XI0/XI25/XI15/NET35_XI0/XI25/XI15/MM8_d
+ N_WL<47>_XI0/XI25/XI15/MM8_g N_BLN<0>_XI0/XI25/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI25/XI15/MM5 N_XI0/XI25/XI15/NET34_XI0/XI25/XI15/MM5_d
+ N_XI0/XI25/XI15/NET33_XI0/XI25/XI15/MM5_g N_VDD_XI0/XI25/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI15/MM4 N_XI0/XI25/XI15/NET33_XI0/XI25/XI15/MM4_d
+ N_XI0/XI25/XI15/NET34_XI0/XI25/XI15/MM4_g N_VDD_XI0/XI25/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI15/MM10 N_XI0/XI25/XI15/NET35_XI0/XI25/XI15/MM10_d
+ N_XI0/XI25/XI15/NET36_XI0/XI25/XI15/MM10_g N_VDD_XI0/XI25/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI25/XI15/MM11 N_XI0/XI25/XI15/NET36_XI0/XI25/XI15/MM11_d
+ N_XI0/XI25/XI15/NET35_XI0/XI25/XI15/MM11_g N_VDD_XI0/XI25/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI0/MM2 N_XI0/XI26/XI0/NET34_XI0/XI26/XI0/MM2_d
+ N_XI0/XI26/XI0/NET33_XI0/XI26/XI0/MM2_g N_VSS_XI0/XI26/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM3 N_XI0/XI26/XI0/NET33_XI0/XI26/XI0/MM3_d
+ N_WL<48>_XI0/XI26/XI0/MM3_g N_BLN<15>_XI0/XI26/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM0 N_XI0/XI26/XI0/NET34_XI0/XI26/XI0/MM0_d
+ N_WL<48>_XI0/XI26/XI0/MM0_g N_BL<15>_XI0/XI26/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM1 N_XI0/XI26/XI0/NET33_XI0/XI26/XI0/MM1_d
+ N_XI0/XI26/XI0/NET34_XI0/XI26/XI0/MM1_g N_VSS_XI0/XI26/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM9 N_XI0/XI26/XI0/NET36_XI0/XI26/XI0/MM9_d
+ N_WL<49>_XI0/XI26/XI0/MM9_g N_BL<15>_XI0/XI26/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM6 N_XI0/XI26/XI0/NET35_XI0/XI26/XI0/MM6_d
+ N_XI0/XI26/XI0/NET36_XI0/XI26/XI0/MM6_g N_VSS_XI0/XI26/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM7 N_XI0/XI26/XI0/NET36_XI0/XI26/XI0/MM7_d
+ N_XI0/XI26/XI0/NET35_XI0/XI26/XI0/MM7_g N_VSS_XI0/XI26/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM8 N_XI0/XI26/XI0/NET35_XI0/XI26/XI0/MM8_d
+ N_WL<49>_XI0/XI26/XI0/MM8_g N_BLN<15>_XI0/XI26/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI0/MM5 N_XI0/XI26/XI0/NET34_XI0/XI26/XI0/MM5_d
+ N_XI0/XI26/XI0/NET33_XI0/XI26/XI0/MM5_g N_VDD_XI0/XI26/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI0/MM4 N_XI0/XI26/XI0/NET33_XI0/XI26/XI0/MM4_d
+ N_XI0/XI26/XI0/NET34_XI0/XI26/XI0/MM4_g N_VDD_XI0/XI26/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI0/MM10 N_XI0/XI26/XI0/NET35_XI0/XI26/XI0/MM10_d
+ N_XI0/XI26/XI0/NET36_XI0/XI26/XI0/MM10_g N_VDD_XI0/XI26/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI0/MM11 N_XI0/XI26/XI0/NET36_XI0/XI26/XI0/MM11_d
+ N_XI0/XI26/XI0/NET35_XI0/XI26/XI0/MM11_g N_VDD_XI0/XI26/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI1/MM2 N_XI0/XI26/XI1/NET34_XI0/XI26/XI1/MM2_d
+ N_XI0/XI26/XI1/NET33_XI0/XI26/XI1/MM2_g N_VSS_XI0/XI26/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM3 N_XI0/XI26/XI1/NET33_XI0/XI26/XI1/MM3_d
+ N_WL<48>_XI0/XI26/XI1/MM3_g N_BLN<14>_XI0/XI26/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM0 N_XI0/XI26/XI1/NET34_XI0/XI26/XI1/MM0_d
+ N_WL<48>_XI0/XI26/XI1/MM0_g N_BL<14>_XI0/XI26/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM1 N_XI0/XI26/XI1/NET33_XI0/XI26/XI1/MM1_d
+ N_XI0/XI26/XI1/NET34_XI0/XI26/XI1/MM1_g N_VSS_XI0/XI26/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM9 N_XI0/XI26/XI1/NET36_XI0/XI26/XI1/MM9_d
+ N_WL<49>_XI0/XI26/XI1/MM9_g N_BL<14>_XI0/XI26/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM6 N_XI0/XI26/XI1/NET35_XI0/XI26/XI1/MM6_d
+ N_XI0/XI26/XI1/NET36_XI0/XI26/XI1/MM6_g N_VSS_XI0/XI26/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM7 N_XI0/XI26/XI1/NET36_XI0/XI26/XI1/MM7_d
+ N_XI0/XI26/XI1/NET35_XI0/XI26/XI1/MM7_g N_VSS_XI0/XI26/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM8 N_XI0/XI26/XI1/NET35_XI0/XI26/XI1/MM8_d
+ N_WL<49>_XI0/XI26/XI1/MM8_g N_BLN<14>_XI0/XI26/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI1/MM5 N_XI0/XI26/XI1/NET34_XI0/XI26/XI1/MM5_d
+ N_XI0/XI26/XI1/NET33_XI0/XI26/XI1/MM5_g N_VDD_XI0/XI26/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI1/MM4 N_XI0/XI26/XI1/NET33_XI0/XI26/XI1/MM4_d
+ N_XI0/XI26/XI1/NET34_XI0/XI26/XI1/MM4_g N_VDD_XI0/XI26/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI1/MM10 N_XI0/XI26/XI1/NET35_XI0/XI26/XI1/MM10_d
+ N_XI0/XI26/XI1/NET36_XI0/XI26/XI1/MM10_g N_VDD_XI0/XI26/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI1/MM11 N_XI0/XI26/XI1/NET36_XI0/XI26/XI1/MM11_d
+ N_XI0/XI26/XI1/NET35_XI0/XI26/XI1/MM11_g N_VDD_XI0/XI26/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI2/MM2 N_XI0/XI26/XI2/NET34_XI0/XI26/XI2/MM2_d
+ N_XI0/XI26/XI2/NET33_XI0/XI26/XI2/MM2_g N_VSS_XI0/XI26/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM3 N_XI0/XI26/XI2/NET33_XI0/XI26/XI2/MM3_d
+ N_WL<48>_XI0/XI26/XI2/MM3_g N_BLN<13>_XI0/XI26/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM0 N_XI0/XI26/XI2/NET34_XI0/XI26/XI2/MM0_d
+ N_WL<48>_XI0/XI26/XI2/MM0_g N_BL<13>_XI0/XI26/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM1 N_XI0/XI26/XI2/NET33_XI0/XI26/XI2/MM1_d
+ N_XI0/XI26/XI2/NET34_XI0/XI26/XI2/MM1_g N_VSS_XI0/XI26/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM9 N_XI0/XI26/XI2/NET36_XI0/XI26/XI2/MM9_d
+ N_WL<49>_XI0/XI26/XI2/MM9_g N_BL<13>_XI0/XI26/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM6 N_XI0/XI26/XI2/NET35_XI0/XI26/XI2/MM6_d
+ N_XI0/XI26/XI2/NET36_XI0/XI26/XI2/MM6_g N_VSS_XI0/XI26/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM7 N_XI0/XI26/XI2/NET36_XI0/XI26/XI2/MM7_d
+ N_XI0/XI26/XI2/NET35_XI0/XI26/XI2/MM7_g N_VSS_XI0/XI26/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM8 N_XI0/XI26/XI2/NET35_XI0/XI26/XI2/MM8_d
+ N_WL<49>_XI0/XI26/XI2/MM8_g N_BLN<13>_XI0/XI26/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI2/MM5 N_XI0/XI26/XI2/NET34_XI0/XI26/XI2/MM5_d
+ N_XI0/XI26/XI2/NET33_XI0/XI26/XI2/MM5_g N_VDD_XI0/XI26/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI2/MM4 N_XI0/XI26/XI2/NET33_XI0/XI26/XI2/MM4_d
+ N_XI0/XI26/XI2/NET34_XI0/XI26/XI2/MM4_g N_VDD_XI0/XI26/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI2/MM10 N_XI0/XI26/XI2/NET35_XI0/XI26/XI2/MM10_d
+ N_XI0/XI26/XI2/NET36_XI0/XI26/XI2/MM10_g N_VDD_XI0/XI26/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI2/MM11 N_XI0/XI26/XI2/NET36_XI0/XI26/XI2/MM11_d
+ N_XI0/XI26/XI2/NET35_XI0/XI26/XI2/MM11_g N_VDD_XI0/XI26/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI3/MM2 N_XI0/XI26/XI3/NET34_XI0/XI26/XI3/MM2_d
+ N_XI0/XI26/XI3/NET33_XI0/XI26/XI3/MM2_g N_VSS_XI0/XI26/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM3 N_XI0/XI26/XI3/NET33_XI0/XI26/XI3/MM3_d
+ N_WL<48>_XI0/XI26/XI3/MM3_g N_BLN<12>_XI0/XI26/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM0 N_XI0/XI26/XI3/NET34_XI0/XI26/XI3/MM0_d
+ N_WL<48>_XI0/XI26/XI3/MM0_g N_BL<12>_XI0/XI26/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM1 N_XI0/XI26/XI3/NET33_XI0/XI26/XI3/MM1_d
+ N_XI0/XI26/XI3/NET34_XI0/XI26/XI3/MM1_g N_VSS_XI0/XI26/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM9 N_XI0/XI26/XI3/NET36_XI0/XI26/XI3/MM9_d
+ N_WL<49>_XI0/XI26/XI3/MM9_g N_BL<12>_XI0/XI26/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM6 N_XI0/XI26/XI3/NET35_XI0/XI26/XI3/MM6_d
+ N_XI0/XI26/XI3/NET36_XI0/XI26/XI3/MM6_g N_VSS_XI0/XI26/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM7 N_XI0/XI26/XI3/NET36_XI0/XI26/XI3/MM7_d
+ N_XI0/XI26/XI3/NET35_XI0/XI26/XI3/MM7_g N_VSS_XI0/XI26/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM8 N_XI0/XI26/XI3/NET35_XI0/XI26/XI3/MM8_d
+ N_WL<49>_XI0/XI26/XI3/MM8_g N_BLN<12>_XI0/XI26/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI3/MM5 N_XI0/XI26/XI3/NET34_XI0/XI26/XI3/MM5_d
+ N_XI0/XI26/XI3/NET33_XI0/XI26/XI3/MM5_g N_VDD_XI0/XI26/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI3/MM4 N_XI0/XI26/XI3/NET33_XI0/XI26/XI3/MM4_d
+ N_XI0/XI26/XI3/NET34_XI0/XI26/XI3/MM4_g N_VDD_XI0/XI26/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI3/MM10 N_XI0/XI26/XI3/NET35_XI0/XI26/XI3/MM10_d
+ N_XI0/XI26/XI3/NET36_XI0/XI26/XI3/MM10_g N_VDD_XI0/XI26/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI3/MM11 N_XI0/XI26/XI3/NET36_XI0/XI26/XI3/MM11_d
+ N_XI0/XI26/XI3/NET35_XI0/XI26/XI3/MM11_g N_VDD_XI0/XI26/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI4/MM2 N_XI0/XI26/XI4/NET34_XI0/XI26/XI4/MM2_d
+ N_XI0/XI26/XI4/NET33_XI0/XI26/XI4/MM2_g N_VSS_XI0/XI26/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM3 N_XI0/XI26/XI4/NET33_XI0/XI26/XI4/MM3_d
+ N_WL<48>_XI0/XI26/XI4/MM3_g N_BLN<11>_XI0/XI26/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM0 N_XI0/XI26/XI4/NET34_XI0/XI26/XI4/MM0_d
+ N_WL<48>_XI0/XI26/XI4/MM0_g N_BL<11>_XI0/XI26/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM1 N_XI0/XI26/XI4/NET33_XI0/XI26/XI4/MM1_d
+ N_XI0/XI26/XI4/NET34_XI0/XI26/XI4/MM1_g N_VSS_XI0/XI26/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM9 N_XI0/XI26/XI4/NET36_XI0/XI26/XI4/MM9_d
+ N_WL<49>_XI0/XI26/XI4/MM9_g N_BL<11>_XI0/XI26/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM6 N_XI0/XI26/XI4/NET35_XI0/XI26/XI4/MM6_d
+ N_XI0/XI26/XI4/NET36_XI0/XI26/XI4/MM6_g N_VSS_XI0/XI26/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM7 N_XI0/XI26/XI4/NET36_XI0/XI26/XI4/MM7_d
+ N_XI0/XI26/XI4/NET35_XI0/XI26/XI4/MM7_g N_VSS_XI0/XI26/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM8 N_XI0/XI26/XI4/NET35_XI0/XI26/XI4/MM8_d
+ N_WL<49>_XI0/XI26/XI4/MM8_g N_BLN<11>_XI0/XI26/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI4/MM5 N_XI0/XI26/XI4/NET34_XI0/XI26/XI4/MM5_d
+ N_XI0/XI26/XI4/NET33_XI0/XI26/XI4/MM5_g N_VDD_XI0/XI26/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI4/MM4 N_XI0/XI26/XI4/NET33_XI0/XI26/XI4/MM4_d
+ N_XI0/XI26/XI4/NET34_XI0/XI26/XI4/MM4_g N_VDD_XI0/XI26/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI4/MM10 N_XI0/XI26/XI4/NET35_XI0/XI26/XI4/MM10_d
+ N_XI0/XI26/XI4/NET36_XI0/XI26/XI4/MM10_g N_VDD_XI0/XI26/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI4/MM11 N_XI0/XI26/XI4/NET36_XI0/XI26/XI4/MM11_d
+ N_XI0/XI26/XI4/NET35_XI0/XI26/XI4/MM11_g N_VDD_XI0/XI26/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI5/MM2 N_XI0/XI26/XI5/NET34_XI0/XI26/XI5/MM2_d
+ N_XI0/XI26/XI5/NET33_XI0/XI26/XI5/MM2_g N_VSS_XI0/XI26/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM3 N_XI0/XI26/XI5/NET33_XI0/XI26/XI5/MM3_d
+ N_WL<48>_XI0/XI26/XI5/MM3_g N_BLN<10>_XI0/XI26/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM0 N_XI0/XI26/XI5/NET34_XI0/XI26/XI5/MM0_d
+ N_WL<48>_XI0/XI26/XI5/MM0_g N_BL<10>_XI0/XI26/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM1 N_XI0/XI26/XI5/NET33_XI0/XI26/XI5/MM1_d
+ N_XI0/XI26/XI5/NET34_XI0/XI26/XI5/MM1_g N_VSS_XI0/XI26/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM9 N_XI0/XI26/XI5/NET36_XI0/XI26/XI5/MM9_d
+ N_WL<49>_XI0/XI26/XI5/MM9_g N_BL<10>_XI0/XI26/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM6 N_XI0/XI26/XI5/NET35_XI0/XI26/XI5/MM6_d
+ N_XI0/XI26/XI5/NET36_XI0/XI26/XI5/MM6_g N_VSS_XI0/XI26/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM7 N_XI0/XI26/XI5/NET36_XI0/XI26/XI5/MM7_d
+ N_XI0/XI26/XI5/NET35_XI0/XI26/XI5/MM7_g N_VSS_XI0/XI26/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM8 N_XI0/XI26/XI5/NET35_XI0/XI26/XI5/MM8_d
+ N_WL<49>_XI0/XI26/XI5/MM8_g N_BLN<10>_XI0/XI26/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI5/MM5 N_XI0/XI26/XI5/NET34_XI0/XI26/XI5/MM5_d
+ N_XI0/XI26/XI5/NET33_XI0/XI26/XI5/MM5_g N_VDD_XI0/XI26/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI5/MM4 N_XI0/XI26/XI5/NET33_XI0/XI26/XI5/MM4_d
+ N_XI0/XI26/XI5/NET34_XI0/XI26/XI5/MM4_g N_VDD_XI0/XI26/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI5/MM10 N_XI0/XI26/XI5/NET35_XI0/XI26/XI5/MM10_d
+ N_XI0/XI26/XI5/NET36_XI0/XI26/XI5/MM10_g N_VDD_XI0/XI26/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI5/MM11 N_XI0/XI26/XI5/NET36_XI0/XI26/XI5/MM11_d
+ N_XI0/XI26/XI5/NET35_XI0/XI26/XI5/MM11_g N_VDD_XI0/XI26/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI6/MM2 N_XI0/XI26/XI6/NET34_XI0/XI26/XI6/MM2_d
+ N_XI0/XI26/XI6/NET33_XI0/XI26/XI6/MM2_g N_VSS_XI0/XI26/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM3 N_XI0/XI26/XI6/NET33_XI0/XI26/XI6/MM3_d
+ N_WL<48>_XI0/XI26/XI6/MM3_g N_BLN<9>_XI0/XI26/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM0 N_XI0/XI26/XI6/NET34_XI0/XI26/XI6/MM0_d
+ N_WL<48>_XI0/XI26/XI6/MM0_g N_BL<9>_XI0/XI26/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM1 N_XI0/XI26/XI6/NET33_XI0/XI26/XI6/MM1_d
+ N_XI0/XI26/XI6/NET34_XI0/XI26/XI6/MM1_g N_VSS_XI0/XI26/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM9 N_XI0/XI26/XI6/NET36_XI0/XI26/XI6/MM9_d
+ N_WL<49>_XI0/XI26/XI6/MM9_g N_BL<9>_XI0/XI26/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM6 N_XI0/XI26/XI6/NET35_XI0/XI26/XI6/MM6_d
+ N_XI0/XI26/XI6/NET36_XI0/XI26/XI6/MM6_g N_VSS_XI0/XI26/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM7 N_XI0/XI26/XI6/NET36_XI0/XI26/XI6/MM7_d
+ N_XI0/XI26/XI6/NET35_XI0/XI26/XI6/MM7_g N_VSS_XI0/XI26/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM8 N_XI0/XI26/XI6/NET35_XI0/XI26/XI6/MM8_d
+ N_WL<49>_XI0/XI26/XI6/MM8_g N_BLN<9>_XI0/XI26/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI6/MM5 N_XI0/XI26/XI6/NET34_XI0/XI26/XI6/MM5_d
+ N_XI0/XI26/XI6/NET33_XI0/XI26/XI6/MM5_g N_VDD_XI0/XI26/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI6/MM4 N_XI0/XI26/XI6/NET33_XI0/XI26/XI6/MM4_d
+ N_XI0/XI26/XI6/NET34_XI0/XI26/XI6/MM4_g N_VDD_XI0/XI26/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI6/MM10 N_XI0/XI26/XI6/NET35_XI0/XI26/XI6/MM10_d
+ N_XI0/XI26/XI6/NET36_XI0/XI26/XI6/MM10_g N_VDD_XI0/XI26/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI6/MM11 N_XI0/XI26/XI6/NET36_XI0/XI26/XI6/MM11_d
+ N_XI0/XI26/XI6/NET35_XI0/XI26/XI6/MM11_g N_VDD_XI0/XI26/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI7/MM2 N_XI0/XI26/XI7/NET34_XI0/XI26/XI7/MM2_d
+ N_XI0/XI26/XI7/NET33_XI0/XI26/XI7/MM2_g N_VSS_XI0/XI26/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM3 N_XI0/XI26/XI7/NET33_XI0/XI26/XI7/MM3_d
+ N_WL<48>_XI0/XI26/XI7/MM3_g N_BLN<8>_XI0/XI26/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM0 N_XI0/XI26/XI7/NET34_XI0/XI26/XI7/MM0_d
+ N_WL<48>_XI0/XI26/XI7/MM0_g N_BL<8>_XI0/XI26/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM1 N_XI0/XI26/XI7/NET33_XI0/XI26/XI7/MM1_d
+ N_XI0/XI26/XI7/NET34_XI0/XI26/XI7/MM1_g N_VSS_XI0/XI26/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM9 N_XI0/XI26/XI7/NET36_XI0/XI26/XI7/MM9_d
+ N_WL<49>_XI0/XI26/XI7/MM9_g N_BL<8>_XI0/XI26/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM6 N_XI0/XI26/XI7/NET35_XI0/XI26/XI7/MM6_d
+ N_XI0/XI26/XI7/NET36_XI0/XI26/XI7/MM6_g N_VSS_XI0/XI26/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM7 N_XI0/XI26/XI7/NET36_XI0/XI26/XI7/MM7_d
+ N_XI0/XI26/XI7/NET35_XI0/XI26/XI7/MM7_g N_VSS_XI0/XI26/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM8 N_XI0/XI26/XI7/NET35_XI0/XI26/XI7/MM8_d
+ N_WL<49>_XI0/XI26/XI7/MM8_g N_BLN<8>_XI0/XI26/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI7/MM5 N_XI0/XI26/XI7/NET34_XI0/XI26/XI7/MM5_d
+ N_XI0/XI26/XI7/NET33_XI0/XI26/XI7/MM5_g N_VDD_XI0/XI26/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI7/MM4 N_XI0/XI26/XI7/NET33_XI0/XI26/XI7/MM4_d
+ N_XI0/XI26/XI7/NET34_XI0/XI26/XI7/MM4_g N_VDD_XI0/XI26/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI7/MM10 N_XI0/XI26/XI7/NET35_XI0/XI26/XI7/MM10_d
+ N_XI0/XI26/XI7/NET36_XI0/XI26/XI7/MM10_g N_VDD_XI0/XI26/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI7/MM11 N_XI0/XI26/XI7/NET36_XI0/XI26/XI7/MM11_d
+ N_XI0/XI26/XI7/NET35_XI0/XI26/XI7/MM11_g N_VDD_XI0/XI26/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI8/MM2 N_XI0/XI26/XI8/NET34_XI0/XI26/XI8/MM2_d
+ N_XI0/XI26/XI8/NET33_XI0/XI26/XI8/MM2_g N_VSS_XI0/XI26/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM3 N_XI0/XI26/XI8/NET33_XI0/XI26/XI8/MM3_d
+ N_WL<48>_XI0/XI26/XI8/MM3_g N_BLN<7>_XI0/XI26/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM0 N_XI0/XI26/XI8/NET34_XI0/XI26/XI8/MM0_d
+ N_WL<48>_XI0/XI26/XI8/MM0_g N_BL<7>_XI0/XI26/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM1 N_XI0/XI26/XI8/NET33_XI0/XI26/XI8/MM1_d
+ N_XI0/XI26/XI8/NET34_XI0/XI26/XI8/MM1_g N_VSS_XI0/XI26/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM9 N_XI0/XI26/XI8/NET36_XI0/XI26/XI8/MM9_d
+ N_WL<49>_XI0/XI26/XI8/MM9_g N_BL<7>_XI0/XI26/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM6 N_XI0/XI26/XI8/NET35_XI0/XI26/XI8/MM6_d
+ N_XI0/XI26/XI8/NET36_XI0/XI26/XI8/MM6_g N_VSS_XI0/XI26/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM7 N_XI0/XI26/XI8/NET36_XI0/XI26/XI8/MM7_d
+ N_XI0/XI26/XI8/NET35_XI0/XI26/XI8/MM7_g N_VSS_XI0/XI26/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM8 N_XI0/XI26/XI8/NET35_XI0/XI26/XI8/MM8_d
+ N_WL<49>_XI0/XI26/XI8/MM8_g N_BLN<7>_XI0/XI26/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI8/MM5 N_XI0/XI26/XI8/NET34_XI0/XI26/XI8/MM5_d
+ N_XI0/XI26/XI8/NET33_XI0/XI26/XI8/MM5_g N_VDD_XI0/XI26/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI8/MM4 N_XI0/XI26/XI8/NET33_XI0/XI26/XI8/MM4_d
+ N_XI0/XI26/XI8/NET34_XI0/XI26/XI8/MM4_g N_VDD_XI0/XI26/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI8/MM10 N_XI0/XI26/XI8/NET35_XI0/XI26/XI8/MM10_d
+ N_XI0/XI26/XI8/NET36_XI0/XI26/XI8/MM10_g N_VDD_XI0/XI26/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI8/MM11 N_XI0/XI26/XI8/NET36_XI0/XI26/XI8/MM11_d
+ N_XI0/XI26/XI8/NET35_XI0/XI26/XI8/MM11_g N_VDD_XI0/XI26/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI9/MM2 N_XI0/XI26/XI9/NET34_XI0/XI26/XI9/MM2_d
+ N_XI0/XI26/XI9/NET33_XI0/XI26/XI9/MM2_g N_VSS_XI0/XI26/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM3 N_XI0/XI26/XI9/NET33_XI0/XI26/XI9/MM3_d
+ N_WL<48>_XI0/XI26/XI9/MM3_g N_BLN<6>_XI0/XI26/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM0 N_XI0/XI26/XI9/NET34_XI0/XI26/XI9/MM0_d
+ N_WL<48>_XI0/XI26/XI9/MM0_g N_BL<6>_XI0/XI26/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM1 N_XI0/XI26/XI9/NET33_XI0/XI26/XI9/MM1_d
+ N_XI0/XI26/XI9/NET34_XI0/XI26/XI9/MM1_g N_VSS_XI0/XI26/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM9 N_XI0/XI26/XI9/NET36_XI0/XI26/XI9/MM9_d
+ N_WL<49>_XI0/XI26/XI9/MM9_g N_BL<6>_XI0/XI26/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM6 N_XI0/XI26/XI9/NET35_XI0/XI26/XI9/MM6_d
+ N_XI0/XI26/XI9/NET36_XI0/XI26/XI9/MM6_g N_VSS_XI0/XI26/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM7 N_XI0/XI26/XI9/NET36_XI0/XI26/XI9/MM7_d
+ N_XI0/XI26/XI9/NET35_XI0/XI26/XI9/MM7_g N_VSS_XI0/XI26/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM8 N_XI0/XI26/XI9/NET35_XI0/XI26/XI9/MM8_d
+ N_WL<49>_XI0/XI26/XI9/MM8_g N_BLN<6>_XI0/XI26/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI9/MM5 N_XI0/XI26/XI9/NET34_XI0/XI26/XI9/MM5_d
+ N_XI0/XI26/XI9/NET33_XI0/XI26/XI9/MM5_g N_VDD_XI0/XI26/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI9/MM4 N_XI0/XI26/XI9/NET33_XI0/XI26/XI9/MM4_d
+ N_XI0/XI26/XI9/NET34_XI0/XI26/XI9/MM4_g N_VDD_XI0/XI26/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI9/MM10 N_XI0/XI26/XI9/NET35_XI0/XI26/XI9/MM10_d
+ N_XI0/XI26/XI9/NET36_XI0/XI26/XI9/MM10_g N_VDD_XI0/XI26/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI9/MM11 N_XI0/XI26/XI9/NET36_XI0/XI26/XI9/MM11_d
+ N_XI0/XI26/XI9/NET35_XI0/XI26/XI9/MM11_g N_VDD_XI0/XI26/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI10/MM2 N_XI0/XI26/XI10/NET34_XI0/XI26/XI10/MM2_d
+ N_XI0/XI26/XI10/NET33_XI0/XI26/XI10/MM2_g N_VSS_XI0/XI26/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM3 N_XI0/XI26/XI10/NET33_XI0/XI26/XI10/MM3_d
+ N_WL<48>_XI0/XI26/XI10/MM3_g N_BLN<5>_XI0/XI26/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM0 N_XI0/XI26/XI10/NET34_XI0/XI26/XI10/MM0_d
+ N_WL<48>_XI0/XI26/XI10/MM0_g N_BL<5>_XI0/XI26/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM1 N_XI0/XI26/XI10/NET33_XI0/XI26/XI10/MM1_d
+ N_XI0/XI26/XI10/NET34_XI0/XI26/XI10/MM1_g N_VSS_XI0/XI26/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM9 N_XI0/XI26/XI10/NET36_XI0/XI26/XI10/MM9_d
+ N_WL<49>_XI0/XI26/XI10/MM9_g N_BL<5>_XI0/XI26/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM6 N_XI0/XI26/XI10/NET35_XI0/XI26/XI10/MM6_d
+ N_XI0/XI26/XI10/NET36_XI0/XI26/XI10/MM6_g N_VSS_XI0/XI26/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM7 N_XI0/XI26/XI10/NET36_XI0/XI26/XI10/MM7_d
+ N_XI0/XI26/XI10/NET35_XI0/XI26/XI10/MM7_g N_VSS_XI0/XI26/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM8 N_XI0/XI26/XI10/NET35_XI0/XI26/XI10/MM8_d
+ N_WL<49>_XI0/XI26/XI10/MM8_g N_BLN<5>_XI0/XI26/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI10/MM5 N_XI0/XI26/XI10/NET34_XI0/XI26/XI10/MM5_d
+ N_XI0/XI26/XI10/NET33_XI0/XI26/XI10/MM5_g N_VDD_XI0/XI26/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI10/MM4 N_XI0/XI26/XI10/NET33_XI0/XI26/XI10/MM4_d
+ N_XI0/XI26/XI10/NET34_XI0/XI26/XI10/MM4_g N_VDD_XI0/XI26/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI10/MM10 N_XI0/XI26/XI10/NET35_XI0/XI26/XI10/MM10_d
+ N_XI0/XI26/XI10/NET36_XI0/XI26/XI10/MM10_g N_VDD_XI0/XI26/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI10/MM11 N_XI0/XI26/XI10/NET36_XI0/XI26/XI10/MM11_d
+ N_XI0/XI26/XI10/NET35_XI0/XI26/XI10/MM11_g N_VDD_XI0/XI26/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI11/MM2 N_XI0/XI26/XI11/NET34_XI0/XI26/XI11/MM2_d
+ N_XI0/XI26/XI11/NET33_XI0/XI26/XI11/MM2_g N_VSS_XI0/XI26/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM3 N_XI0/XI26/XI11/NET33_XI0/XI26/XI11/MM3_d
+ N_WL<48>_XI0/XI26/XI11/MM3_g N_BLN<4>_XI0/XI26/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM0 N_XI0/XI26/XI11/NET34_XI0/XI26/XI11/MM0_d
+ N_WL<48>_XI0/XI26/XI11/MM0_g N_BL<4>_XI0/XI26/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM1 N_XI0/XI26/XI11/NET33_XI0/XI26/XI11/MM1_d
+ N_XI0/XI26/XI11/NET34_XI0/XI26/XI11/MM1_g N_VSS_XI0/XI26/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM9 N_XI0/XI26/XI11/NET36_XI0/XI26/XI11/MM9_d
+ N_WL<49>_XI0/XI26/XI11/MM9_g N_BL<4>_XI0/XI26/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM6 N_XI0/XI26/XI11/NET35_XI0/XI26/XI11/MM6_d
+ N_XI0/XI26/XI11/NET36_XI0/XI26/XI11/MM6_g N_VSS_XI0/XI26/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM7 N_XI0/XI26/XI11/NET36_XI0/XI26/XI11/MM7_d
+ N_XI0/XI26/XI11/NET35_XI0/XI26/XI11/MM7_g N_VSS_XI0/XI26/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM8 N_XI0/XI26/XI11/NET35_XI0/XI26/XI11/MM8_d
+ N_WL<49>_XI0/XI26/XI11/MM8_g N_BLN<4>_XI0/XI26/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI11/MM5 N_XI0/XI26/XI11/NET34_XI0/XI26/XI11/MM5_d
+ N_XI0/XI26/XI11/NET33_XI0/XI26/XI11/MM5_g N_VDD_XI0/XI26/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI11/MM4 N_XI0/XI26/XI11/NET33_XI0/XI26/XI11/MM4_d
+ N_XI0/XI26/XI11/NET34_XI0/XI26/XI11/MM4_g N_VDD_XI0/XI26/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI11/MM10 N_XI0/XI26/XI11/NET35_XI0/XI26/XI11/MM10_d
+ N_XI0/XI26/XI11/NET36_XI0/XI26/XI11/MM10_g N_VDD_XI0/XI26/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI11/MM11 N_XI0/XI26/XI11/NET36_XI0/XI26/XI11/MM11_d
+ N_XI0/XI26/XI11/NET35_XI0/XI26/XI11/MM11_g N_VDD_XI0/XI26/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI12/MM2 N_XI0/XI26/XI12/NET34_XI0/XI26/XI12/MM2_d
+ N_XI0/XI26/XI12/NET33_XI0/XI26/XI12/MM2_g N_VSS_XI0/XI26/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM3 N_XI0/XI26/XI12/NET33_XI0/XI26/XI12/MM3_d
+ N_WL<48>_XI0/XI26/XI12/MM3_g N_BLN<3>_XI0/XI26/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM0 N_XI0/XI26/XI12/NET34_XI0/XI26/XI12/MM0_d
+ N_WL<48>_XI0/XI26/XI12/MM0_g N_BL<3>_XI0/XI26/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM1 N_XI0/XI26/XI12/NET33_XI0/XI26/XI12/MM1_d
+ N_XI0/XI26/XI12/NET34_XI0/XI26/XI12/MM1_g N_VSS_XI0/XI26/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM9 N_XI0/XI26/XI12/NET36_XI0/XI26/XI12/MM9_d
+ N_WL<49>_XI0/XI26/XI12/MM9_g N_BL<3>_XI0/XI26/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM6 N_XI0/XI26/XI12/NET35_XI0/XI26/XI12/MM6_d
+ N_XI0/XI26/XI12/NET36_XI0/XI26/XI12/MM6_g N_VSS_XI0/XI26/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM7 N_XI0/XI26/XI12/NET36_XI0/XI26/XI12/MM7_d
+ N_XI0/XI26/XI12/NET35_XI0/XI26/XI12/MM7_g N_VSS_XI0/XI26/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM8 N_XI0/XI26/XI12/NET35_XI0/XI26/XI12/MM8_d
+ N_WL<49>_XI0/XI26/XI12/MM8_g N_BLN<3>_XI0/XI26/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI12/MM5 N_XI0/XI26/XI12/NET34_XI0/XI26/XI12/MM5_d
+ N_XI0/XI26/XI12/NET33_XI0/XI26/XI12/MM5_g N_VDD_XI0/XI26/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI12/MM4 N_XI0/XI26/XI12/NET33_XI0/XI26/XI12/MM4_d
+ N_XI0/XI26/XI12/NET34_XI0/XI26/XI12/MM4_g N_VDD_XI0/XI26/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI12/MM10 N_XI0/XI26/XI12/NET35_XI0/XI26/XI12/MM10_d
+ N_XI0/XI26/XI12/NET36_XI0/XI26/XI12/MM10_g N_VDD_XI0/XI26/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI12/MM11 N_XI0/XI26/XI12/NET36_XI0/XI26/XI12/MM11_d
+ N_XI0/XI26/XI12/NET35_XI0/XI26/XI12/MM11_g N_VDD_XI0/XI26/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI13/MM2 N_XI0/XI26/XI13/NET34_XI0/XI26/XI13/MM2_d
+ N_XI0/XI26/XI13/NET33_XI0/XI26/XI13/MM2_g N_VSS_XI0/XI26/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM3 N_XI0/XI26/XI13/NET33_XI0/XI26/XI13/MM3_d
+ N_WL<48>_XI0/XI26/XI13/MM3_g N_BLN<2>_XI0/XI26/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM0 N_XI0/XI26/XI13/NET34_XI0/XI26/XI13/MM0_d
+ N_WL<48>_XI0/XI26/XI13/MM0_g N_BL<2>_XI0/XI26/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM1 N_XI0/XI26/XI13/NET33_XI0/XI26/XI13/MM1_d
+ N_XI0/XI26/XI13/NET34_XI0/XI26/XI13/MM1_g N_VSS_XI0/XI26/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM9 N_XI0/XI26/XI13/NET36_XI0/XI26/XI13/MM9_d
+ N_WL<49>_XI0/XI26/XI13/MM9_g N_BL<2>_XI0/XI26/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM6 N_XI0/XI26/XI13/NET35_XI0/XI26/XI13/MM6_d
+ N_XI0/XI26/XI13/NET36_XI0/XI26/XI13/MM6_g N_VSS_XI0/XI26/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM7 N_XI0/XI26/XI13/NET36_XI0/XI26/XI13/MM7_d
+ N_XI0/XI26/XI13/NET35_XI0/XI26/XI13/MM7_g N_VSS_XI0/XI26/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM8 N_XI0/XI26/XI13/NET35_XI0/XI26/XI13/MM8_d
+ N_WL<49>_XI0/XI26/XI13/MM8_g N_BLN<2>_XI0/XI26/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI13/MM5 N_XI0/XI26/XI13/NET34_XI0/XI26/XI13/MM5_d
+ N_XI0/XI26/XI13/NET33_XI0/XI26/XI13/MM5_g N_VDD_XI0/XI26/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI13/MM4 N_XI0/XI26/XI13/NET33_XI0/XI26/XI13/MM4_d
+ N_XI0/XI26/XI13/NET34_XI0/XI26/XI13/MM4_g N_VDD_XI0/XI26/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI13/MM10 N_XI0/XI26/XI13/NET35_XI0/XI26/XI13/MM10_d
+ N_XI0/XI26/XI13/NET36_XI0/XI26/XI13/MM10_g N_VDD_XI0/XI26/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI13/MM11 N_XI0/XI26/XI13/NET36_XI0/XI26/XI13/MM11_d
+ N_XI0/XI26/XI13/NET35_XI0/XI26/XI13/MM11_g N_VDD_XI0/XI26/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI14/MM2 N_XI0/XI26/XI14/NET34_XI0/XI26/XI14/MM2_d
+ N_XI0/XI26/XI14/NET33_XI0/XI26/XI14/MM2_g N_VSS_XI0/XI26/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM3 N_XI0/XI26/XI14/NET33_XI0/XI26/XI14/MM3_d
+ N_WL<48>_XI0/XI26/XI14/MM3_g N_BLN<1>_XI0/XI26/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM0 N_XI0/XI26/XI14/NET34_XI0/XI26/XI14/MM0_d
+ N_WL<48>_XI0/XI26/XI14/MM0_g N_BL<1>_XI0/XI26/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM1 N_XI0/XI26/XI14/NET33_XI0/XI26/XI14/MM1_d
+ N_XI0/XI26/XI14/NET34_XI0/XI26/XI14/MM1_g N_VSS_XI0/XI26/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM9 N_XI0/XI26/XI14/NET36_XI0/XI26/XI14/MM9_d
+ N_WL<49>_XI0/XI26/XI14/MM9_g N_BL<1>_XI0/XI26/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM6 N_XI0/XI26/XI14/NET35_XI0/XI26/XI14/MM6_d
+ N_XI0/XI26/XI14/NET36_XI0/XI26/XI14/MM6_g N_VSS_XI0/XI26/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM7 N_XI0/XI26/XI14/NET36_XI0/XI26/XI14/MM7_d
+ N_XI0/XI26/XI14/NET35_XI0/XI26/XI14/MM7_g N_VSS_XI0/XI26/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM8 N_XI0/XI26/XI14/NET35_XI0/XI26/XI14/MM8_d
+ N_WL<49>_XI0/XI26/XI14/MM8_g N_BLN<1>_XI0/XI26/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI14/MM5 N_XI0/XI26/XI14/NET34_XI0/XI26/XI14/MM5_d
+ N_XI0/XI26/XI14/NET33_XI0/XI26/XI14/MM5_g N_VDD_XI0/XI26/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI14/MM4 N_XI0/XI26/XI14/NET33_XI0/XI26/XI14/MM4_d
+ N_XI0/XI26/XI14/NET34_XI0/XI26/XI14/MM4_g N_VDD_XI0/XI26/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI14/MM10 N_XI0/XI26/XI14/NET35_XI0/XI26/XI14/MM10_d
+ N_XI0/XI26/XI14/NET36_XI0/XI26/XI14/MM10_g N_VDD_XI0/XI26/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI14/MM11 N_XI0/XI26/XI14/NET36_XI0/XI26/XI14/MM11_d
+ N_XI0/XI26/XI14/NET35_XI0/XI26/XI14/MM11_g N_VDD_XI0/XI26/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI15/MM2 N_XI0/XI26/XI15/NET34_XI0/XI26/XI15/MM2_d
+ N_XI0/XI26/XI15/NET33_XI0/XI26/XI15/MM2_g N_VSS_XI0/XI26/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM3 N_XI0/XI26/XI15/NET33_XI0/XI26/XI15/MM3_d
+ N_WL<48>_XI0/XI26/XI15/MM3_g N_BLN<0>_XI0/XI26/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM0 N_XI0/XI26/XI15/NET34_XI0/XI26/XI15/MM0_d
+ N_WL<48>_XI0/XI26/XI15/MM0_g N_BL<0>_XI0/XI26/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM1 N_XI0/XI26/XI15/NET33_XI0/XI26/XI15/MM1_d
+ N_XI0/XI26/XI15/NET34_XI0/XI26/XI15/MM1_g N_VSS_XI0/XI26/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM9 N_XI0/XI26/XI15/NET36_XI0/XI26/XI15/MM9_d
+ N_WL<49>_XI0/XI26/XI15/MM9_g N_BL<0>_XI0/XI26/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM6 N_XI0/XI26/XI15/NET35_XI0/XI26/XI15/MM6_d
+ N_XI0/XI26/XI15/NET36_XI0/XI26/XI15/MM6_g N_VSS_XI0/XI26/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM7 N_XI0/XI26/XI15/NET36_XI0/XI26/XI15/MM7_d
+ N_XI0/XI26/XI15/NET35_XI0/XI26/XI15/MM7_g N_VSS_XI0/XI26/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM8 N_XI0/XI26/XI15/NET35_XI0/XI26/XI15/MM8_d
+ N_WL<49>_XI0/XI26/XI15/MM8_g N_BLN<0>_XI0/XI26/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI26/XI15/MM5 N_XI0/XI26/XI15/NET34_XI0/XI26/XI15/MM5_d
+ N_XI0/XI26/XI15/NET33_XI0/XI26/XI15/MM5_g N_VDD_XI0/XI26/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI15/MM4 N_XI0/XI26/XI15/NET33_XI0/XI26/XI15/MM4_d
+ N_XI0/XI26/XI15/NET34_XI0/XI26/XI15/MM4_g N_VDD_XI0/XI26/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI15/MM10 N_XI0/XI26/XI15/NET35_XI0/XI26/XI15/MM10_d
+ N_XI0/XI26/XI15/NET36_XI0/XI26/XI15/MM10_g N_VDD_XI0/XI26/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI26/XI15/MM11 N_XI0/XI26/XI15/NET36_XI0/XI26/XI15/MM11_d
+ N_XI0/XI26/XI15/NET35_XI0/XI26/XI15/MM11_g N_VDD_XI0/XI26/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI0/MM2 N_XI0/XI27/XI0/NET34_XI0/XI27/XI0/MM2_d
+ N_XI0/XI27/XI0/NET33_XI0/XI27/XI0/MM2_g N_VSS_XI0/XI27/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM3 N_XI0/XI27/XI0/NET33_XI0/XI27/XI0/MM3_d
+ N_WL<50>_XI0/XI27/XI0/MM3_g N_BLN<15>_XI0/XI27/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM0 N_XI0/XI27/XI0/NET34_XI0/XI27/XI0/MM0_d
+ N_WL<50>_XI0/XI27/XI0/MM0_g N_BL<15>_XI0/XI27/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM1 N_XI0/XI27/XI0/NET33_XI0/XI27/XI0/MM1_d
+ N_XI0/XI27/XI0/NET34_XI0/XI27/XI0/MM1_g N_VSS_XI0/XI27/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM9 N_XI0/XI27/XI0/NET36_XI0/XI27/XI0/MM9_d
+ N_WL<51>_XI0/XI27/XI0/MM9_g N_BL<15>_XI0/XI27/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM6 N_XI0/XI27/XI0/NET35_XI0/XI27/XI0/MM6_d
+ N_XI0/XI27/XI0/NET36_XI0/XI27/XI0/MM6_g N_VSS_XI0/XI27/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM7 N_XI0/XI27/XI0/NET36_XI0/XI27/XI0/MM7_d
+ N_XI0/XI27/XI0/NET35_XI0/XI27/XI0/MM7_g N_VSS_XI0/XI27/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM8 N_XI0/XI27/XI0/NET35_XI0/XI27/XI0/MM8_d
+ N_WL<51>_XI0/XI27/XI0/MM8_g N_BLN<15>_XI0/XI27/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI0/MM5 N_XI0/XI27/XI0/NET34_XI0/XI27/XI0/MM5_d
+ N_XI0/XI27/XI0/NET33_XI0/XI27/XI0/MM5_g N_VDD_XI0/XI27/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI0/MM4 N_XI0/XI27/XI0/NET33_XI0/XI27/XI0/MM4_d
+ N_XI0/XI27/XI0/NET34_XI0/XI27/XI0/MM4_g N_VDD_XI0/XI27/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI0/MM10 N_XI0/XI27/XI0/NET35_XI0/XI27/XI0/MM10_d
+ N_XI0/XI27/XI0/NET36_XI0/XI27/XI0/MM10_g N_VDD_XI0/XI27/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI0/MM11 N_XI0/XI27/XI0/NET36_XI0/XI27/XI0/MM11_d
+ N_XI0/XI27/XI0/NET35_XI0/XI27/XI0/MM11_g N_VDD_XI0/XI27/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI1/MM2 N_XI0/XI27/XI1/NET34_XI0/XI27/XI1/MM2_d
+ N_XI0/XI27/XI1/NET33_XI0/XI27/XI1/MM2_g N_VSS_XI0/XI27/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM3 N_XI0/XI27/XI1/NET33_XI0/XI27/XI1/MM3_d
+ N_WL<50>_XI0/XI27/XI1/MM3_g N_BLN<14>_XI0/XI27/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM0 N_XI0/XI27/XI1/NET34_XI0/XI27/XI1/MM0_d
+ N_WL<50>_XI0/XI27/XI1/MM0_g N_BL<14>_XI0/XI27/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM1 N_XI0/XI27/XI1/NET33_XI0/XI27/XI1/MM1_d
+ N_XI0/XI27/XI1/NET34_XI0/XI27/XI1/MM1_g N_VSS_XI0/XI27/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM9 N_XI0/XI27/XI1/NET36_XI0/XI27/XI1/MM9_d
+ N_WL<51>_XI0/XI27/XI1/MM9_g N_BL<14>_XI0/XI27/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM6 N_XI0/XI27/XI1/NET35_XI0/XI27/XI1/MM6_d
+ N_XI0/XI27/XI1/NET36_XI0/XI27/XI1/MM6_g N_VSS_XI0/XI27/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM7 N_XI0/XI27/XI1/NET36_XI0/XI27/XI1/MM7_d
+ N_XI0/XI27/XI1/NET35_XI0/XI27/XI1/MM7_g N_VSS_XI0/XI27/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM8 N_XI0/XI27/XI1/NET35_XI0/XI27/XI1/MM8_d
+ N_WL<51>_XI0/XI27/XI1/MM8_g N_BLN<14>_XI0/XI27/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI1/MM5 N_XI0/XI27/XI1/NET34_XI0/XI27/XI1/MM5_d
+ N_XI0/XI27/XI1/NET33_XI0/XI27/XI1/MM5_g N_VDD_XI0/XI27/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI1/MM4 N_XI0/XI27/XI1/NET33_XI0/XI27/XI1/MM4_d
+ N_XI0/XI27/XI1/NET34_XI0/XI27/XI1/MM4_g N_VDD_XI0/XI27/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI1/MM10 N_XI0/XI27/XI1/NET35_XI0/XI27/XI1/MM10_d
+ N_XI0/XI27/XI1/NET36_XI0/XI27/XI1/MM10_g N_VDD_XI0/XI27/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI1/MM11 N_XI0/XI27/XI1/NET36_XI0/XI27/XI1/MM11_d
+ N_XI0/XI27/XI1/NET35_XI0/XI27/XI1/MM11_g N_VDD_XI0/XI27/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI2/MM2 N_XI0/XI27/XI2/NET34_XI0/XI27/XI2/MM2_d
+ N_XI0/XI27/XI2/NET33_XI0/XI27/XI2/MM2_g N_VSS_XI0/XI27/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM3 N_XI0/XI27/XI2/NET33_XI0/XI27/XI2/MM3_d
+ N_WL<50>_XI0/XI27/XI2/MM3_g N_BLN<13>_XI0/XI27/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM0 N_XI0/XI27/XI2/NET34_XI0/XI27/XI2/MM0_d
+ N_WL<50>_XI0/XI27/XI2/MM0_g N_BL<13>_XI0/XI27/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM1 N_XI0/XI27/XI2/NET33_XI0/XI27/XI2/MM1_d
+ N_XI0/XI27/XI2/NET34_XI0/XI27/XI2/MM1_g N_VSS_XI0/XI27/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM9 N_XI0/XI27/XI2/NET36_XI0/XI27/XI2/MM9_d
+ N_WL<51>_XI0/XI27/XI2/MM9_g N_BL<13>_XI0/XI27/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM6 N_XI0/XI27/XI2/NET35_XI0/XI27/XI2/MM6_d
+ N_XI0/XI27/XI2/NET36_XI0/XI27/XI2/MM6_g N_VSS_XI0/XI27/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM7 N_XI0/XI27/XI2/NET36_XI0/XI27/XI2/MM7_d
+ N_XI0/XI27/XI2/NET35_XI0/XI27/XI2/MM7_g N_VSS_XI0/XI27/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM8 N_XI0/XI27/XI2/NET35_XI0/XI27/XI2/MM8_d
+ N_WL<51>_XI0/XI27/XI2/MM8_g N_BLN<13>_XI0/XI27/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI2/MM5 N_XI0/XI27/XI2/NET34_XI0/XI27/XI2/MM5_d
+ N_XI0/XI27/XI2/NET33_XI0/XI27/XI2/MM5_g N_VDD_XI0/XI27/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI2/MM4 N_XI0/XI27/XI2/NET33_XI0/XI27/XI2/MM4_d
+ N_XI0/XI27/XI2/NET34_XI0/XI27/XI2/MM4_g N_VDD_XI0/XI27/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI2/MM10 N_XI0/XI27/XI2/NET35_XI0/XI27/XI2/MM10_d
+ N_XI0/XI27/XI2/NET36_XI0/XI27/XI2/MM10_g N_VDD_XI0/XI27/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI2/MM11 N_XI0/XI27/XI2/NET36_XI0/XI27/XI2/MM11_d
+ N_XI0/XI27/XI2/NET35_XI0/XI27/XI2/MM11_g N_VDD_XI0/XI27/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI3/MM2 N_XI0/XI27/XI3/NET34_XI0/XI27/XI3/MM2_d
+ N_XI0/XI27/XI3/NET33_XI0/XI27/XI3/MM2_g N_VSS_XI0/XI27/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM3 N_XI0/XI27/XI3/NET33_XI0/XI27/XI3/MM3_d
+ N_WL<50>_XI0/XI27/XI3/MM3_g N_BLN<12>_XI0/XI27/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM0 N_XI0/XI27/XI3/NET34_XI0/XI27/XI3/MM0_d
+ N_WL<50>_XI0/XI27/XI3/MM0_g N_BL<12>_XI0/XI27/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM1 N_XI0/XI27/XI3/NET33_XI0/XI27/XI3/MM1_d
+ N_XI0/XI27/XI3/NET34_XI0/XI27/XI3/MM1_g N_VSS_XI0/XI27/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM9 N_XI0/XI27/XI3/NET36_XI0/XI27/XI3/MM9_d
+ N_WL<51>_XI0/XI27/XI3/MM9_g N_BL<12>_XI0/XI27/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM6 N_XI0/XI27/XI3/NET35_XI0/XI27/XI3/MM6_d
+ N_XI0/XI27/XI3/NET36_XI0/XI27/XI3/MM6_g N_VSS_XI0/XI27/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM7 N_XI0/XI27/XI3/NET36_XI0/XI27/XI3/MM7_d
+ N_XI0/XI27/XI3/NET35_XI0/XI27/XI3/MM7_g N_VSS_XI0/XI27/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM8 N_XI0/XI27/XI3/NET35_XI0/XI27/XI3/MM8_d
+ N_WL<51>_XI0/XI27/XI3/MM8_g N_BLN<12>_XI0/XI27/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI3/MM5 N_XI0/XI27/XI3/NET34_XI0/XI27/XI3/MM5_d
+ N_XI0/XI27/XI3/NET33_XI0/XI27/XI3/MM5_g N_VDD_XI0/XI27/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI3/MM4 N_XI0/XI27/XI3/NET33_XI0/XI27/XI3/MM4_d
+ N_XI0/XI27/XI3/NET34_XI0/XI27/XI3/MM4_g N_VDD_XI0/XI27/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI3/MM10 N_XI0/XI27/XI3/NET35_XI0/XI27/XI3/MM10_d
+ N_XI0/XI27/XI3/NET36_XI0/XI27/XI3/MM10_g N_VDD_XI0/XI27/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI3/MM11 N_XI0/XI27/XI3/NET36_XI0/XI27/XI3/MM11_d
+ N_XI0/XI27/XI3/NET35_XI0/XI27/XI3/MM11_g N_VDD_XI0/XI27/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI4/MM2 N_XI0/XI27/XI4/NET34_XI0/XI27/XI4/MM2_d
+ N_XI0/XI27/XI4/NET33_XI0/XI27/XI4/MM2_g N_VSS_XI0/XI27/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM3 N_XI0/XI27/XI4/NET33_XI0/XI27/XI4/MM3_d
+ N_WL<50>_XI0/XI27/XI4/MM3_g N_BLN<11>_XI0/XI27/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM0 N_XI0/XI27/XI4/NET34_XI0/XI27/XI4/MM0_d
+ N_WL<50>_XI0/XI27/XI4/MM0_g N_BL<11>_XI0/XI27/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM1 N_XI0/XI27/XI4/NET33_XI0/XI27/XI4/MM1_d
+ N_XI0/XI27/XI4/NET34_XI0/XI27/XI4/MM1_g N_VSS_XI0/XI27/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM9 N_XI0/XI27/XI4/NET36_XI0/XI27/XI4/MM9_d
+ N_WL<51>_XI0/XI27/XI4/MM9_g N_BL<11>_XI0/XI27/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM6 N_XI0/XI27/XI4/NET35_XI0/XI27/XI4/MM6_d
+ N_XI0/XI27/XI4/NET36_XI0/XI27/XI4/MM6_g N_VSS_XI0/XI27/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM7 N_XI0/XI27/XI4/NET36_XI0/XI27/XI4/MM7_d
+ N_XI0/XI27/XI4/NET35_XI0/XI27/XI4/MM7_g N_VSS_XI0/XI27/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM8 N_XI0/XI27/XI4/NET35_XI0/XI27/XI4/MM8_d
+ N_WL<51>_XI0/XI27/XI4/MM8_g N_BLN<11>_XI0/XI27/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI4/MM5 N_XI0/XI27/XI4/NET34_XI0/XI27/XI4/MM5_d
+ N_XI0/XI27/XI4/NET33_XI0/XI27/XI4/MM5_g N_VDD_XI0/XI27/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI4/MM4 N_XI0/XI27/XI4/NET33_XI0/XI27/XI4/MM4_d
+ N_XI0/XI27/XI4/NET34_XI0/XI27/XI4/MM4_g N_VDD_XI0/XI27/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI4/MM10 N_XI0/XI27/XI4/NET35_XI0/XI27/XI4/MM10_d
+ N_XI0/XI27/XI4/NET36_XI0/XI27/XI4/MM10_g N_VDD_XI0/XI27/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI4/MM11 N_XI0/XI27/XI4/NET36_XI0/XI27/XI4/MM11_d
+ N_XI0/XI27/XI4/NET35_XI0/XI27/XI4/MM11_g N_VDD_XI0/XI27/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI5/MM2 N_XI0/XI27/XI5/NET34_XI0/XI27/XI5/MM2_d
+ N_XI0/XI27/XI5/NET33_XI0/XI27/XI5/MM2_g N_VSS_XI0/XI27/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM3 N_XI0/XI27/XI5/NET33_XI0/XI27/XI5/MM3_d
+ N_WL<50>_XI0/XI27/XI5/MM3_g N_BLN<10>_XI0/XI27/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM0 N_XI0/XI27/XI5/NET34_XI0/XI27/XI5/MM0_d
+ N_WL<50>_XI0/XI27/XI5/MM0_g N_BL<10>_XI0/XI27/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM1 N_XI0/XI27/XI5/NET33_XI0/XI27/XI5/MM1_d
+ N_XI0/XI27/XI5/NET34_XI0/XI27/XI5/MM1_g N_VSS_XI0/XI27/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM9 N_XI0/XI27/XI5/NET36_XI0/XI27/XI5/MM9_d
+ N_WL<51>_XI0/XI27/XI5/MM9_g N_BL<10>_XI0/XI27/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM6 N_XI0/XI27/XI5/NET35_XI0/XI27/XI5/MM6_d
+ N_XI0/XI27/XI5/NET36_XI0/XI27/XI5/MM6_g N_VSS_XI0/XI27/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM7 N_XI0/XI27/XI5/NET36_XI0/XI27/XI5/MM7_d
+ N_XI0/XI27/XI5/NET35_XI0/XI27/XI5/MM7_g N_VSS_XI0/XI27/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM8 N_XI0/XI27/XI5/NET35_XI0/XI27/XI5/MM8_d
+ N_WL<51>_XI0/XI27/XI5/MM8_g N_BLN<10>_XI0/XI27/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI5/MM5 N_XI0/XI27/XI5/NET34_XI0/XI27/XI5/MM5_d
+ N_XI0/XI27/XI5/NET33_XI0/XI27/XI5/MM5_g N_VDD_XI0/XI27/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI5/MM4 N_XI0/XI27/XI5/NET33_XI0/XI27/XI5/MM4_d
+ N_XI0/XI27/XI5/NET34_XI0/XI27/XI5/MM4_g N_VDD_XI0/XI27/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI5/MM10 N_XI0/XI27/XI5/NET35_XI0/XI27/XI5/MM10_d
+ N_XI0/XI27/XI5/NET36_XI0/XI27/XI5/MM10_g N_VDD_XI0/XI27/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI5/MM11 N_XI0/XI27/XI5/NET36_XI0/XI27/XI5/MM11_d
+ N_XI0/XI27/XI5/NET35_XI0/XI27/XI5/MM11_g N_VDD_XI0/XI27/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI6/MM2 N_XI0/XI27/XI6/NET34_XI0/XI27/XI6/MM2_d
+ N_XI0/XI27/XI6/NET33_XI0/XI27/XI6/MM2_g N_VSS_XI0/XI27/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM3 N_XI0/XI27/XI6/NET33_XI0/XI27/XI6/MM3_d
+ N_WL<50>_XI0/XI27/XI6/MM3_g N_BLN<9>_XI0/XI27/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM0 N_XI0/XI27/XI6/NET34_XI0/XI27/XI6/MM0_d
+ N_WL<50>_XI0/XI27/XI6/MM0_g N_BL<9>_XI0/XI27/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM1 N_XI0/XI27/XI6/NET33_XI0/XI27/XI6/MM1_d
+ N_XI0/XI27/XI6/NET34_XI0/XI27/XI6/MM1_g N_VSS_XI0/XI27/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM9 N_XI0/XI27/XI6/NET36_XI0/XI27/XI6/MM9_d
+ N_WL<51>_XI0/XI27/XI6/MM9_g N_BL<9>_XI0/XI27/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM6 N_XI0/XI27/XI6/NET35_XI0/XI27/XI6/MM6_d
+ N_XI0/XI27/XI6/NET36_XI0/XI27/XI6/MM6_g N_VSS_XI0/XI27/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM7 N_XI0/XI27/XI6/NET36_XI0/XI27/XI6/MM7_d
+ N_XI0/XI27/XI6/NET35_XI0/XI27/XI6/MM7_g N_VSS_XI0/XI27/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM8 N_XI0/XI27/XI6/NET35_XI0/XI27/XI6/MM8_d
+ N_WL<51>_XI0/XI27/XI6/MM8_g N_BLN<9>_XI0/XI27/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI6/MM5 N_XI0/XI27/XI6/NET34_XI0/XI27/XI6/MM5_d
+ N_XI0/XI27/XI6/NET33_XI0/XI27/XI6/MM5_g N_VDD_XI0/XI27/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI6/MM4 N_XI0/XI27/XI6/NET33_XI0/XI27/XI6/MM4_d
+ N_XI0/XI27/XI6/NET34_XI0/XI27/XI6/MM4_g N_VDD_XI0/XI27/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI6/MM10 N_XI0/XI27/XI6/NET35_XI0/XI27/XI6/MM10_d
+ N_XI0/XI27/XI6/NET36_XI0/XI27/XI6/MM10_g N_VDD_XI0/XI27/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI6/MM11 N_XI0/XI27/XI6/NET36_XI0/XI27/XI6/MM11_d
+ N_XI0/XI27/XI6/NET35_XI0/XI27/XI6/MM11_g N_VDD_XI0/XI27/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI7/MM2 N_XI0/XI27/XI7/NET34_XI0/XI27/XI7/MM2_d
+ N_XI0/XI27/XI7/NET33_XI0/XI27/XI7/MM2_g N_VSS_XI0/XI27/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM3 N_XI0/XI27/XI7/NET33_XI0/XI27/XI7/MM3_d
+ N_WL<50>_XI0/XI27/XI7/MM3_g N_BLN<8>_XI0/XI27/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM0 N_XI0/XI27/XI7/NET34_XI0/XI27/XI7/MM0_d
+ N_WL<50>_XI0/XI27/XI7/MM0_g N_BL<8>_XI0/XI27/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM1 N_XI0/XI27/XI7/NET33_XI0/XI27/XI7/MM1_d
+ N_XI0/XI27/XI7/NET34_XI0/XI27/XI7/MM1_g N_VSS_XI0/XI27/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM9 N_XI0/XI27/XI7/NET36_XI0/XI27/XI7/MM9_d
+ N_WL<51>_XI0/XI27/XI7/MM9_g N_BL<8>_XI0/XI27/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM6 N_XI0/XI27/XI7/NET35_XI0/XI27/XI7/MM6_d
+ N_XI0/XI27/XI7/NET36_XI0/XI27/XI7/MM6_g N_VSS_XI0/XI27/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM7 N_XI0/XI27/XI7/NET36_XI0/XI27/XI7/MM7_d
+ N_XI0/XI27/XI7/NET35_XI0/XI27/XI7/MM7_g N_VSS_XI0/XI27/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM8 N_XI0/XI27/XI7/NET35_XI0/XI27/XI7/MM8_d
+ N_WL<51>_XI0/XI27/XI7/MM8_g N_BLN<8>_XI0/XI27/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI7/MM5 N_XI0/XI27/XI7/NET34_XI0/XI27/XI7/MM5_d
+ N_XI0/XI27/XI7/NET33_XI0/XI27/XI7/MM5_g N_VDD_XI0/XI27/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI7/MM4 N_XI0/XI27/XI7/NET33_XI0/XI27/XI7/MM4_d
+ N_XI0/XI27/XI7/NET34_XI0/XI27/XI7/MM4_g N_VDD_XI0/XI27/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI7/MM10 N_XI0/XI27/XI7/NET35_XI0/XI27/XI7/MM10_d
+ N_XI0/XI27/XI7/NET36_XI0/XI27/XI7/MM10_g N_VDD_XI0/XI27/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI7/MM11 N_XI0/XI27/XI7/NET36_XI0/XI27/XI7/MM11_d
+ N_XI0/XI27/XI7/NET35_XI0/XI27/XI7/MM11_g N_VDD_XI0/XI27/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI8/MM2 N_XI0/XI27/XI8/NET34_XI0/XI27/XI8/MM2_d
+ N_XI0/XI27/XI8/NET33_XI0/XI27/XI8/MM2_g N_VSS_XI0/XI27/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM3 N_XI0/XI27/XI8/NET33_XI0/XI27/XI8/MM3_d
+ N_WL<50>_XI0/XI27/XI8/MM3_g N_BLN<7>_XI0/XI27/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM0 N_XI0/XI27/XI8/NET34_XI0/XI27/XI8/MM0_d
+ N_WL<50>_XI0/XI27/XI8/MM0_g N_BL<7>_XI0/XI27/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM1 N_XI0/XI27/XI8/NET33_XI0/XI27/XI8/MM1_d
+ N_XI0/XI27/XI8/NET34_XI0/XI27/XI8/MM1_g N_VSS_XI0/XI27/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM9 N_XI0/XI27/XI8/NET36_XI0/XI27/XI8/MM9_d
+ N_WL<51>_XI0/XI27/XI8/MM9_g N_BL<7>_XI0/XI27/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM6 N_XI0/XI27/XI8/NET35_XI0/XI27/XI8/MM6_d
+ N_XI0/XI27/XI8/NET36_XI0/XI27/XI8/MM6_g N_VSS_XI0/XI27/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM7 N_XI0/XI27/XI8/NET36_XI0/XI27/XI8/MM7_d
+ N_XI0/XI27/XI8/NET35_XI0/XI27/XI8/MM7_g N_VSS_XI0/XI27/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM8 N_XI0/XI27/XI8/NET35_XI0/XI27/XI8/MM8_d
+ N_WL<51>_XI0/XI27/XI8/MM8_g N_BLN<7>_XI0/XI27/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI8/MM5 N_XI0/XI27/XI8/NET34_XI0/XI27/XI8/MM5_d
+ N_XI0/XI27/XI8/NET33_XI0/XI27/XI8/MM5_g N_VDD_XI0/XI27/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI8/MM4 N_XI0/XI27/XI8/NET33_XI0/XI27/XI8/MM4_d
+ N_XI0/XI27/XI8/NET34_XI0/XI27/XI8/MM4_g N_VDD_XI0/XI27/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI8/MM10 N_XI0/XI27/XI8/NET35_XI0/XI27/XI8/MM10_d
+ N_XI0/XI27/XI8/NET36_XI0/XI27/XI8/MM10_g N_VDD_XI0/XI27/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI8/MM11 N_XI0/XI27/XI8/NET36_XI0/XI27/XI8/MM11_d
+ N_XI0/XI27/XI8/NET35_XI0/XI27/XI8/MM11_g N_VDD_XI0/XI27/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI9/MM2 N_XI0/XI27/XI9/NET34_XI0/XI27/XI9/MM2_d
+ N_XI0/XI27/XI9/NET33_XI0/XI27/XI9/MM2_g N_VSS_XI0/XI27/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM3 N_XI0/XI27/XI9/NET33_XI0/XI27/XI9/MM3_d
+ N_WL<50>_XI0/XI27/XI9/MM3_g N_BLN<6>_XI0/XI27/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM0 N_XI0/XI27/XI9/NET34_XI0/XI27/XI9/MM0_d
+ N_WL<50>_XI0/XI27/XI9/MM0_g N_BL<6>_XI0/XI27/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM1 N_XI0/XI27/XI9/NET33_XI0/XI27/XI9/MM1_d
+ N_XI0/XI27/XI9/NET34_XI0/XI27/XI9/MM1_g N_VSS_XI0/XI27/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM9 N_XI0/XI27/XI9/NET36_XI0/XI27/XI9/MM9_d
+ N_WL<51>_XI0/XI27/XI9/MM9_g N_BL<6>_XI0/XI27/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM6 N_XI0/XI27/XI9/NET35_XI0/XI27/XI9/MM6_d
+ N_XI0/XI27/XI9/NET36_XI0/XI27/XI9/MM6_g N_VSS_XI0/XI27/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM7 N_XI0/XI27/XI9/NET36_XI0/XI27/XI9/MM7_d
+ N_XI0/XI27/XI9/NET35_XI0/XI27/XI9/MM7_g N_VSS_XI0/XI27/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM8 N_XI0/XI27/XI9/NET35_XI0/XI27/XI9/MM8_d
+ N_WL<51>_XI0/XI27/XI9/MM8_g N_BLN<6>_XI0/XI27/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI9/MM5 N_XI0/XI27/XI9/NET34_XI0/XI27/XI9/MM5_d
+ N_XI0/XI27/XI9/NET33_XI0/XI27/XI9/MM5_g N_VDD_XI0/XI27/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI9/MM4 N_XI0/XI27/XI9/NET33_XI0/XI27/XI9/MM4_d
+ N_XI0/XI27/XI9/NET34_XI0/XI27/XI9/MM4_g N_VDD_XI0/XI27/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI9/MM10 N_XI0/XI27/XI9/NET35_XI0/XI27/XI9/MM10_d
+ N_XI0/XI27/XI9/NET36_XI0/XI27/XI9/MM10_g N_VDD_XI0/XI27/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI9/MM11 N_XI0/XI27/XI9/NET36_XI0/XI27/XI9/MM11_d
+ N_XI0/XI27/XI9/NET35_XI0/XI27/XI9/MM11_g N_VDD_XI0/XI27/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI10/MM2 N_XI0/XI27/XI10/NET34_XI0/XI27/XI10/MM2_d
+ N_XI0/XI27/XI10/NET33_XI0/XI27/XI10/MM2_g N_VSS_XI0/XI27/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM3 N_XI0/XI27/XI10/NET33_XI0/XI27/XI10/MM3_d
+ N_WL<50>_XI0/XI27/XI10/MM3_g N_BLN<5>_XI0/XI27/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM0 N_XI0/XI27/XI10/NET34_XI0/XI27/XI10/MM0_d
+ N_WL<50>_XI0/XI27/XI10/MM0_g N_BL<5>_XI0/XI27/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM1 N_XI0/XI27/XI10/NET33_XI0/XI27/XI10/MM1_d
+ N_XI0/XI27/XI10/NET34_XI0/XI27/XI10/MM1_g N_VSS_XI0/XI27/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM9 N_XI0/XI27/XI10/NET36_XI0/XI27/XI10/MM9_d
+ N_WL<51>_XI0/XI27/XI10/MM9_g N_BL<5>_XI0/XI27/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM6 N_XI0/XI27/XI10/NET35_XI0/XI27/XI10/MM6_d
+ N_XI0/XI27/XI10/NET36_XI0/XI27/XI10/MM6_g N_VSS_XI0/XI27/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM7 N_XI0/XI27/XI10/NET36_XI0/XI27/XI10/MM7_d
+ N_XI0/XI27/XI10/NET35_XI0/XI27/XI10/MM7_g N_VSS_XI0/XI27/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM8 N_XI0/XI27/XI10/NET35_XI0/XI27/XI10/MM8_d
+ N_WL<51>_XI0/XI27/XI10/MM8_g N_BLN<5>_XI0/XI27/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI10/MM5 N_XI0/XI27/XI10/NET34_XI0/XI27/XI10/MM5_d
+ N_XI0/XI27/XI10/NET33_XI0/XI27/XI10/MM5_g N_VDD_XI0/XI27/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI10/MM4 N_XI0/XI27/XI10/NET33_XI0/XI27/XI10/MM4_d
+ N_XI0/XI27/XI10/NET34_XI0/XI27/XI10/MM4_g N_VDD_XI0/XI27/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI10/MM10 N_XI0/XI27/XI10/NET35_XI0/XI27/XI10/MM10_d
+ N_XI0/XI27/XI10/NET36_XI0/XI27/XI10/MM10_g N_VDD_XI0/XI27/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI10/MM11 N_XI0/XI27/XI10/NET36_XI0/XI27/XI10/MM11_d
+ N_XI0/XI27/XI10/NET35_XI0/XI27/XI10/MM11_g N_VDD_XI0/XI27/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI11/MM2 N_XI0/XI27/XI11/NET34_XI0/XI27/XI11/MM2_d
+ N_XI0/XI27/XI11/NET33_XI0/XI27/XI11/MM2_g N_VSS_XI0/XI27/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM3 N_XI0/XI27/XI11/NET33_XI0/XI27/XI11/MM3_d
+ N_WL<50>_XI0/XI27/XI11/MM3_g N_BLN<4>_XI0/XI27/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM0 N_XI0/XI27/XI11/NET34_XI0/XI27/XI11/MM0_d
+ N_WL<50>_XI0/XI27/XI11/MM0_g N_BL<4>_XI0/XI27/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM1 N_XI0/XI27/XI11/NET33_XI0/XI27/XI11/MM1_d
+ N_XI0/XI27/XI11/NET34_XI0/XI27/XI11/MM1_g N_VSS_XI0/XI27/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM9 N_XI0/XI27/XI11/NET36_XI0/XI27/XI11/MM9_d
+ N_WL<51>_XI0/XI27/XI11/MM9_g N_BL<4>_XI0/XI27/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM6 N_XI0/XI27/XI11/NET35_XI0/XI27/XI11/MM6_d
+ N_XI0/XI27/XI11/NET36_XI0/XI27/XI11/MM6_g N_VSS_XI0/XI27/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM7 N_XI0/XI27/XI11/NET36_XI0/XI27/XI11/MM7_d
+ N_XI0/XI27/XI11/NET35_XI0/XI27/XI11/MM7_g N_VSS_XI0/XI27/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM8 N_XI0/XI27/XI11/NET35_XI0/XI27/XI11/MM8_d
+ N_WL<51>_XI0/XI27/XI11/MM8_g N_BLN<4>_XI0/XI27/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI11/MM5 N_XI0/XI27/XI11/NET34_XI0/XI27/XI11/MM5_d
+ N_XI0/XI27/XI11/NET33_XI0/XI27/XI11/MM5_g N_VDD_XI0/XI27/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI11/MM4 N_XI0/XI27/XI11/NET33_XI0/XI27/XI11/MM4_d
+ N_XI0/XI27/XI11/NET34_XI0/XI27/XI11/MM4_g N_VDD_XI0/XI27/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI11/MM10 N_XI0/XI27/XI11/NET35_XI0/XI27/XI11/MM10_d
+ N_XI0/XI27/XI11/NET36_XI0/XI27/XI11/MM10_g N_VDD_XI0/XI27/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI11/MM11 N_XI0/XI27/XI11/NET36_XI0/XI27/XI11/MM11_d
+ N_XI0/XI27/XI11/NET35_XI0/XI27/XI11/MM11_g N_VDD_XI0/XI27/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI12/MM2 N_XI0/XI27/XI12/NET34_XI0/XI27/XI12/MM2_d
+ N_XI0/XI27/XI12/NET33_XI0/XI27/XI12/MM2_g N_VSS_XI0/XI27/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM3 N_XI0/XI27/XI12/NET33_XI0/XI27/XI12/MM3_d
+ N_WL<50>_XI0/XI27/XI12/MM3_g N_BLN<3>_XI0/XI27/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM0 N_XI0/XI27/XI12/NET34_XI0/XI27/XI12/MM0_d
+ N_WL<50>_XI0/XI27/XI12/MM0_g N_BL<3>_XI0/XI27/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM1 N_XI0/XI27/XI12/NET33_XI0/XI27/XI12/MM1_d
+ N_XI0/XI27/XI12/NET34_XI0/XI27/XI12/MM1_g N_VSS_XI0/XI27/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM9 N_XI0/XI27/XI12/NET36_XI0/XI27/XI12/MM9_d
+ N_WL<51>_XI0/XI27/XI12/MM9_g N_BL<3>_XI0/XI27/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM6 N_XI0/XI27/XI12/NET35_XI0/XI27/XI12/MM6_d
+ N_XI0/XI27/XI12/NET36_XI0/XI27/XI12/MM6_g N_VSS_XI0/XI27/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM7 N_XI0/XI27/XI12/NET36_XI0/XI27/XI12/MM7_d
+ N_XI0/XI27/XI12/NET35_XI0/XI27/XI12/MM7_g N_VSS_XI0/XI27/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM8 N_XI0/XI27/XI12/NET35_XI0/XI27/XI12/MM8_d
+ N_WL<51>_XI0/XI27/XI12/MM8_g N_BLN<3>_XI0/XI27/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI12/MM5 N_XI0/XI27/XI12/NET34_XI0/XI27/XI12/MM5_d
+ N_XI0/XI27/XI12/NET33_XI0/XI27/XI12/MM5_g N_VDD_XI0/XI27/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI12/MM4 N_XI0/XI27/XI12/NET33_XI0/XI27/XI12/MM4_d
+ N_XI0/XI27/XI12/NET34_XI0/XI27/XI12/MM4_g N_VDD_XI0/XI27/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI12/MM10 N_XI0/XI27/XI12/NET35_XI0/XI27/XI12/MM10_d
+ N_XI0/XI27/XI12/NET36_XI0/XI27/XI12/MM10_g N_VDD_XI0/XI27/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI12/MM11 N_XI0/XI27/XI12/NET36_XI0/XI27/XI12/MM11_d
+ N_XI0/XI27/XI12/NET35_XI0/XI27/XI12/MM11_g N_VDD_XI0/XI27/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI13/MM2 N_XI0/XI27/XI13/NET34_XI0/XI27/XI13/MM2_d
+ N_XI0/XI27/XI13/NET33_XI0/XI27/XI13/MM2_g N_VSS_XI0/XI27/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM3 N_XI0/XI27/XI13/NET33_XI0/XI27/XI13/MM3_d
+ N_WL<50>_XI0/XI27/XI13/MM3_g N_BLN<2>_XI0/XI27/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM0 N_XI0/XI27/XI13/NET34_XI0/XI27/XI13/MM0_d
+ N_WL<50>_XI0/XI27/XI13/MM0_g N_BL<2>_XI0/XI27/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM1 N_XI0/XI27/XI13/NET33_XI0/XI27/XI13/MM1_d
+ N_XI0/XI27/XI13/NET34_XI0/XI27/XI13/MM1_g N_VSS_XI0/XI27/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM9 N_XI0/XI27/XI13/NET36_XI0/XI27/XI13/MM9_d
+ N_WL<51>_XI0/XI27/XI13/MM9_g N_BL<2>_XI0/XI27/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM6 N_XI0/XI27/XI13/NET35_XI0/XI27/XI13/MM6_d
+ N_XI0/XI27/XI13/NET36_XI0/XI27/XI13/MM6_g N_VSS_XI0/XI27/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM7 N_XI0/XI27/XI13/NET36_XI0/XI27/XI13/MM7_d
+ N_XI0/XI27/XI13/NET35_XI0/XI27/XI13/MM7_g N_VSS_XI0/XI27/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM8 N_XI0/XI27/XI13/NET35_XI0/XI27/XI13/MM8_d
+ N_WL<51>_XI0/XI27/XI13/MM8_g N_BLN<2>_XI0/XI27/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI13/MM5 N_XI0/XI27/XI13/NET34_XI0/XI27/XI13/MM5_d
+ N_XI0/XI27/XI13/NET33_XI0/XI27/XI13/MM5_g N_VDD_XI0/XI27/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI13/MM4 N_XI0/XI27/XI13/NET33_XI0/XI27/XI13/MM4_d
+ N_XI0/XI27/XI13/NET34_XI0/XI27/XI13/MM4_g N_VDD_XI0/XI27/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI13/MM10 N_XI0/XI27/XI13/NET35_XI0/XI27/XI13/MM10_d
+ N_XI0/XI27/XI13/NET36_XI0/XI27/XI13/MM10_g N_VDD_XI0/XI27/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI13/MM11 N_XI0/XI27/XI13/NET36_XI0/XI27/XI13/MM11_d
+ N_XI0/XI27/XI13/NET35_XI0/XI27/XI13/MM11_g N_VDD_XI0/XI27/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI14/MM2 N_XI0/XI27/XI14/NET34_XI0/XI27/XI14/MM2_d
+ N_XI0/XI27/XI14/NET33_XI0/XI27/XI14/MM2_g N_VSS_XI0/XI27/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM3 N_XI0/XI27/XI14/NET33_XI0/XI27/XI14/MM3_d
+ N_WL<50>_XI0/XI27/XI14/MM3_g N_BLN<1>_XI0/XI27/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM0 N_XI0/XI27/XI14/NET34_XI0/XI27/XI14/MM0_d
+ N_WL<50>_XI0/XI27/XI14/MM0_g N_BL<1>_XI0/XI27/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM1 N_XI0/XI27/XI14/NET33_XI0/XI27/XI14/MM1_d
+ N_XI0/XI27/XI14/NET34_XI0/XI27/XI14/MM1_g N_VSS_XI0/XI27/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM9 N_XI0/XI27/XI14/NET36_XI0/XI27/XI14/MM9_d
+ N_WL<51>_XI0/XI27/XI14/MM9_g N_BL<1>_XI0/XI27/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM6 N_XI0/XI27/XI14/NET35_XI0/XI27/XI14/MM6_d
+ N_XI0/XI27/XI14/NET36_XI0/XI27/XI14/MM6_g N_VSS_XI0/XI27/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM7 N_XI0/XI27/XI14/NET36_XI0/XI27/XI14/MM7_d
+ N_XI0/XI27/XI14/NET35_XI0/XI27/XI14/MM7_g N_VSS_XI0/XI27/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM8 N_XI0/XI27/XI14/NET35_XI0/XI27/XI14/MM8_d
+ N_WL<51>_XI0/XI27/XI14/MM8_g N_BLN<1>_XI0/XI27/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI14/MM5 N_XI0/XI27/XI14/NET34_XI0/XI27/XI14/MM5_d
+ N_XI0/XI27/XI14/NET33_XI0/XI27/XI14/MM5_g N_VDD_XI0/XI27/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI14/MM4 N_XI0/XI27/XI14/NET33_XI0/XI27/XI14/MM4_d
+ N_XI0/XI27/XI14/NET34_XI0/XI27/XI14/MM4_g N_VDD_XI0/XI27/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI14/MM10 N_XI0/XI27/XI14/NET35_XI0/XI27/XI14/MM10_d
+ N_XI0/XI27/XI14/NET36_XI0/XI27/XI14/MM10_g N_VDD_XI0/XI27/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI14/MM11 N_XI0/XI27/XI14/NET36_XI0/XI27/XI14/MM11_d
+ N_XI0/XI27/XI14/NET35_XI0/XI27/XI14/MM11_g N_VDD_XI0/XI27/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI15/MM2 N_XI0/XI27/XI15/NET34_XI0/XI27/XI15/MM2_d
+ N_XI0/XI27/XI15/NET33_XI0/XI27/XI15/MM2_g N_VSS_XI0/XI27/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM3 N_XI0/XI27/XI15/NET33_XI0/XI27/XI15/MM3_d
+ N_WL<50>_XI0/XI27/XI15/MM3_g N_BLN<0>_XI0/XI27/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM0 N_XI0/XI27/XI15/NET34_XI0/XI27/XI15/MM0_d
+ N_WL<50>_XI0/XI27/XI15/MM0_g N_BL<0>_XI0/XI27/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM1 N_XI0/XI27/XI15/NET33_XI0/XI27/XI15/MM1_d
+ N_XI0/XI27/XI15/NET34_XI0/XI27/XI15/MM1_g N_VSS_XI0/XI27/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM9 N_XI0/XI27/XI15/NET36_XI0/XI27/XI15/MM9_d
+ N_WL<51>_XI0/XI27/XI15/MM9_g N_BL<0>_XI0/XI27/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM6 N_XI0/XI27/XI15/NET35_XI0/XI27/XI15/MM6_d
+ N_XI0/XI27/XI15/NET36_XI0/XI27/XI15/MM6_g N_VSS_XI0/XI27/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM7 N_XI0/XI27/XI15/NET36_XI0/XI27/XI15/MM7_d
+ N_XI0/XI27/XI15/NET35_XI0/XI27/XI15/MM7_g N_VSS_XI0/XI27/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM8 N_XI0/XI27/XI15/NET35_XI0/XI27/XI15/MM8_d
+ N_WL<51>_XI0/XI27/XI15/MM8_g N_BLN<0>_XI0/XI27/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI27/XI15/MM5 N_XI0/XI27/XI15/NET34_XI0/XI27/XI15/MM5_d
+ N_XI0/XI27/XI15/NET33_XI0/XI27/XI15/MM5_g N_VDD_XI0/XI27/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI15/MM4 N_XI0/XI27/XI15/NET33_XI0/XI27/XI15/MM4_d
+ N_XI0/XI27/XI15/NET34_XI0/XI27/XI15/MM4_g N_VDD_XI0/XI27/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI15/MM10 N_XI0/XI27/XI15/NET35_XI0/XI27/XI15/MM10_d
+ N_XI0/XI27/XI15/NET36_XI0/XI27/XI15/MM10_g N_VDD_XI0/XI27/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI27/XI15/MM11 N_XI0/XI27/XI15/NET36_XI0/XI27/XI15/MM11_d
+ N_XI0/XI27/XI15/NET35_XI0/XI27/XI15/MM11_g N_VDD_XI0/XI27/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI0/MM2 N_XI0/XI28/XI0/NET34_XI0/XI28/XI0/MM2_d
+ N_XI0/XI28/XI0/NET33_XI0/XI28/XI0/MM2_g N_VSS_XI0/XI28/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM3 N_XI0/XI28/XI0/NET33_XI0/XI28/XI0/MM3_d
+ N_WL<52>_XI0/XI28/XI0/MM3_g N_BLN<15>_XI0/XI28/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM0 N_XI0/XI28/XI0/NET34_XI0/XI28/XI0/MM0_d
+ N_WL<52>_XI0/XI28/XI0/MM0_g N_BL<15>_XI0/XI28/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM1 N_XI0/XI28/XI0/NET33_XI0/XI28/XI0/MM1_d
+ N_XI0/XI28/XI0/NET34_XI0/XI28/XI0/MM1_g N_VSS_XI0/XI28/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM9 N_XI0/XI28/XI0/NET36_XI0/XI28/XI0/MM9_d
+ N_WL<53>_XI0/XI28/XI0/MM9_g N_BL<15>_XI0/XI28/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM6 N_XI0/XI28/XI0/NET35_XI0/XI28/XI0/MM6_d
+ N_XI0/XI28/XI0/NET36_XI0/XI28/XI0/MM6_g N_VSS_XI0/XI28/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM7 N_XI0/XI28/XI0/NET36_XI0/XI28/XI0/MM7_d
+ N_XI0/XI28/XI0/NET35_XI0/XI28/XI0/MM7_g N_VSS_XI0/XI28/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM8 N_XI0/XI28/XI0/NET35_XI0/XI28/XI0/MM8_d
+ N_WL<53>_XI0/XI28/XI0/MM8_g N_BLN<15>_XI0/XI28/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI0/MM5 N_XI0/XI28/XI0/NET34_XI0/XI28/XI0/MM5_d
+ N_XI0/XI28/XI0/NET33_XI0/XI28/XI0/MM5_g N_VDD_XI0/XI28/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI0/MM4 N_XI0/XI28/XI0/NET33_XI0/XI28/XI0/MM4_d
+ N_XI0/XI28/XI0/NET34_XI0/XI28/XI0/MM4_g N_VDD_XI0/XI28/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI0/MM10 N_XI0/XI28/XI0/NET35_XI0/XI28/XI0/MM10_d
+ N_XI0/XI28/XI0/NET36_XI0/XI28/XI0/MM10_g N_VDD_XI0/XI28/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI0/MM11 N_XI0/XI28/XI0/NET36_XI0/XI28/XI0/MM11_d
+ N_XI0/XI28/XI0/NET35_XI0/XI28/XI0/MM11_g N_VDD_XI0/XI28/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI1/MM2 N_XI0/XI28/XI1/NET34_XI0/XI28/XI1/MM2_d
+ N_XI0/XI28/XI1/NET33_XI0/XI28/XI1/MM2_g N_VSS_XI0/XI28/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM3 N_XI0/XI28/XI1/NET33_XI0/XI28/XI1/MM3_d
+ N_WL<52>_XI0/XI28/XI1/MM3_g N_BLN<14>_XI0/XI28/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM0 N_XI0/XI28/XI1/NET34_XI0/XI28/XI1/MM0_d
+ N_WL<52>_XI0/XI28/XI1/MM0_g N_BL<14>_XI0/XI28/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM1 N_XI0/XI28/XI1/NET33_XI0/XI28/XI1/MM1_d
+ N_XI0/XI28/XI1/NET34_XI0/XI28/XI1/MM1_g N_VSS_XI0/XI28/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM9 N_XI0/XI28/XI1/NET36_XI0/XI28/XI1/MM9_d
+ N_WL<53>_XI0/XI28/XI1/MM9_g N_BL<14>_XI0/XI28/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM6 N_XI0/XI28/XI1/NET35_XI0/XI28/XI1/MM6_d
+ N_XI0/XI28/XI1/NET36_XI0/XI28/XI1/MM6_g N_VSS_XI0/XI28/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM7 N_XI0/XI28/XI1/NET36_XI0/XI28/XI1/MM7_d
+ N_XI0/XI28/XI1/NET35_XI0/XI28/XI1/MM7_g N_VSS_XI0/XI28/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM8 N_XI0/XI28/XI1/NET35_XI0/XI28/XI1/MM8_d
+ N_WL<53>_XI0/XI28/XI1/MM8_g N_BLN<14>_XI0/XI28/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI1/MM5 N_XI0/XI28/XI1/NET34_XI0/XI28/XI1/MM5_d
+ N_XI0/XI28/XI1/NET33_XI0/XI28/XI1/MM5_g N_VDD_XI0/XI28/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI1/MM4 N_XI0/XI28/XI1/NET33_XI0/XI28/XI1/MM4_d
+ N_XI0/XI28/XI1/NET34_XI0/XI28/XI1/MM4_g N_VDD_XI0/XI28/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI1/MM10 N_XI0/XI28/XI1/NET35_XI0/XI28/XI1/MM10_d
+ N_XI0/XI28/XI1/NET36_XI0/XI28/XI1/MM10_g N_VDD_XI0/XI28/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI1/MM11 N_XI0/XI28/XI1/NET36_XI0/XI28/XI1/MM11_d
+ N_XI0/XI28/XI1/NET35_XI0/XI28/XI1/MM11_g N_VDD_XI0/XI28/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI2/MM2 N_XI0/XI28/XI2/NET34_XI0/XI28/XI2/MM2_d
+ N_XI0/XI28/XI2/NET33_XI0/XI28/XI2/MM2_g N_VSS_XI0/XI28/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM3 N_XI0/XI28/XI2/NET33_XI0/XI28/XI2/MM3_d
+ N_WL<52>_XI0/XI28/XI2/MM3_g N_BLN<13>_XI0/XI28/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM0 N_XI0/XI28/XI2/NET34_XI0/XI28/XI2/MM0_d
+ N_WL<52>_XI0/XI28/XI2/MM0_g N_BL<13>_XI0/XI28/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM1 N_XI0/XI28/XI2/NET33_XI0/XI28/XI2/MM1_d
+ N_XI0/XI28/XI2/NET34_XI0/XI28/XI2/MM1_g N_VSS_XI0/XI28/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM9 N_XI0/XI28/XI2/NET36_XI0/XI28/XI2/MM9_d
+ N_WL<53>_XI0/XI28/XI2/MM9_g N_BL<13>_XI0/XI28/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM6 N_XI0/XI28/XI2/NET35_XI0/XI28/XI2/MM6_d
+ N_XI0/XI28/XI2/NET36_XI0/XI28/XI2/MM6_g N_VSS_XI0/XI28/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM7 N_XI0/XI28/XI2/NET36_XI0/XI28/XI2/MM7_d
+ N_XI0/XI28/XI2/NET35_XI0/XI28/XI2/MM7_g N_VSS_XI0/XI28/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM8 N_XI0/XI28/XI2/NET35_XI0/XI28/XI2/MM8_d
+ N_WL<53>_XI0/XI28/XI2/MM8_g N_BLN<13>_XI0/XI28/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI2/MM5 N_XI0/XI28/XI2/NET34_XI0/XI28/XI2/MM5_d
+ N_XI0/XI28/XI2/NET33_XI0/XI28/XI2/MM5_g N_VDD_XI0/XI28/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI2/MM4 N_XI0/XI28/XI2/NET33_XI0/XI28/XI2/MM4_d
+ N_XI0/XI28/XI2/NET34_XI0/XI28/XI2/MM4_g N_VDD_XI0/XI28/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI2/MM10 N_XI0/XI28/XI2/NET35_XI0/XI28/XI2/MM10_d
+ N_XI0/XI28/XI2/NET36_XI0/XI28/XI2/MM10_g N_VDD_XI0/XI28/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI2/MM11 N_XI0/XI28/XI2/NET36_XI0/XI28/XI2/MM11_d
+ N_XI0/XI28/XI2/NET35_XI0/XI28/XI2/MM11_g N_VDD_XI0/XI28/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI3/MM2 N_XI0/XI28/XI3/NET34_XI0/XI28/XI3/MM2_d
+ N_XI0/XI28/XI3/NET33_XI0/XI28/XI3/MM2_g N_VSS_XI0/XI28/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM3 N_XI0/XI28/XI3/NET33_XI0/XI28/XI3/MM3_d
+ N_WL<52>_XI0/XI28/XI3/MM3_g N_BLN<12>_XI0/XI28/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM0 N_XI0/XI28/XI3/NET34_XI0/XI28/XI3/MM0_d
+ N_WL<52>_XI0/XI28/XI3/MM0_g N_BL<12>_XI0/XI28/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM1 N_XI0/XI28/XI3/NET33_XI0/XI28/XI3/MM1_d
+ N_XI0/XI28/XI3/NET34_XI0/XI28/XI3/MM1_g N_VSS_XI0/XI28/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM9 N_XI0/XI28/XI3/NET36_XI0/XI28/XI3/MM9_d
+ N_WL<53>_XI0/XI28/XI3/MM9_g N_BL<12>_XI0/XI28/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM6 N_XI0/XI28/XI3/NET35_XI0/XI28/XI3/MM6_d
+ N_XI0/XI28/XI3/NET36_XI0/XI28/XI3/MM6_g N_VSS_XI0/XI28/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM7 N_XI0/XI28/XI3/NET36_XI0/XI28/XI3/MM7_d
+ N_XI0/XI28/XI3/NET35_XI0/XI28/XI3/MM7_g N_VSS_XI0/XI28/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM8 N_XI0/XI28/XI3/NET35_XI0/XI28/XI3/MM8_d
+ N_WL<53>_XI0/XI28/XI3/MM8_g N_BLN<12>_XI0/XI28/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI3/MM5 N_XI0/XI28/XI3/NET34_XI0/XI28/XI3/MM5_d
+ N_XI0/XI28/XI3/NET33_XI0/XI28/XI3/MM5_g N_VDD_XI0/XI28/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI3/MM4 N_XI0/XI28/XI3/NET33_XI0/XI28/XI3/MM4_d
+ N_XI0/XI28/XI3/NET34_XI0/XI28/XI3/MM4_g N_VDD_XI0/XI28/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI3/MM10 N_XI0/XI28/XI3/NET35_XI0/XI28/XI3/MM10_d
+ N_XI0/XI28/XI3/NET36_XI0/XI28/XI3/MM10_g N_VDD_XI0/XI28/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI3/MM11 N_XI0/XI28/XI3/NET36_XI0/XI28/XI3/MM11_d
+ N_XI0/XI28/XI3/NET35_XI0/XI28/XI3/MM11_g N_VDD_XI0/XI28/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI4/MM2 N_XI0/XI28/XI4/NET34_XI0/XI28/XI4/MM2_d
+ N_XI0/XI28/XI4/NET33_XI0/XI28/XI4/MM2_g N_VSS_XI0/XI28/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM3 N_XI0/XI28/XI4/NET33_XI0/XI28/XI4/MM3_d
+ N_WL<52>_XI0/XI28/XI4/MM3_g N_BLN<11>_XI0/XI28/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM0 N_XI0/XI28/XI4/NET34_XI0/XI28/XI4/MM0_d
+ N_WL<52>_XI0/XI28/XI4/MM0_g N_BL<11>_XI0/XI28/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM1 N_XI0/XI28/XI4/NET33_XI0/XI28/XI4/MM1_d
+ N_XI0/XI28/XI4/NET34_XI0/XI28/XI4/MM1_g N_VSS_XI0/XI28/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM9 N_XI0/XI28/XI4/NET36_XI0/XI28/XI4/MM9_d
+ N_WL<53>_XI0/XI28/XI4/MM9_g N_BL<11>_XI0/XI28/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM6 N_XI0/XI28/XI4/NET35_XI0/XI28/XI4/MM6_d
+ N_XI0/XI28/XI4/NET36_XI0/XI28/XI4/MM6_g N_VSS_XI0/XI28/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM7 N_XI0/XI28/XI4/NET36_XI0/XI28/XI4/MM7_d
+ N_XI0/XI28/XI4/NET35_XI0/XI28/XI4/MM7_g N_VSS_XI0/XI28/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM8 N_XI0/XI28/XI4/NET35_XI0/XI28/XI4/MM8_d
+ N_WL<53>_XI0/XI28/XI4/MM8_g N_BLN<11>_XI0/XI28/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI4/MM5 N_XI0/XI28/XI4/NET34_XI0/XI28/XI4/MM5_d
+ N_XI0/XI28/XI4/NET33_XI0/XI28/XI4/MM5_g N_VDD_XI0/XI28/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI4/MM4 N_XI0/XI28/XI4/NET33_XI0/XI28/XI4/MM4_d
+ N_XI0/XI28/XI4/NET34_XI0/XI28/XI4/MM4_g N_VDD_XI0/XI28/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI4/MM10 N_XI0/XI28/XI4/NET35_XI0/XI28/XI4/MM10_d
+ N_XI0/XI28/XI4/NET36_XI0/XI28/XI4/MM10_g N_VDD_XI0/XI28/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI4/MM11 N_XI0/XI28/XI4/NET36_XI0/XI28/XI4/MM11_d
+ N_XI0/XI28/XI4/NET35_XI0/XI28/XI4/MM11_g N_VDD_XI0/XI28/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI5/MM2 N_XI0/XI28/XI5/NET34_XI0/XI28/XI5/MM2_d
+ N_XI0/XI28/XI5/NET33_XI0/XI28/XI5/MM2_g N_VSS_XI0/XI28/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM3 N_XI0/XI28/XI5/NET33_XI0/XI28/XI5/MM3_d
+ N_WL<52>_XI0/XI28/XI5/MM3_g N_BLN<10>_XI0/XI28/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM0 N_XI0/XI28/XI5/NET34_XI0/XI28/XI5/MM0_d
+ N_WL<52>_XI0/XI28/XI5/MM0_g N_BL<10>_XI0/XI28/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM1 N_XI0/XI28/XI5/NET33_XI0/XI28/XI5/MM1_d
+ N_XI0/XI28/XI5/NET34_XI0/XI28/XI5/MM1_g N_VSS_XI0/XI28/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM9 N_XI0/XI28/XI5/NET36_XI0/XI28/XI5/MM9_d
+ N_WL<53>_XI0/XI28/XI5/MM9_g N_BL<10>_XI0/XI28/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM6 N_XI0/XI28/XI5/NET35_XI0/XI28/XI5/MM6_d
+ N_XI0/XI28/XI5/NET36_XI0/XI28/XI5/MM6_g N_VSS_XI0/XI28/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM7 N_XI0/XI28/XI5/NET36_XI0/XI28/XI5/MM7_d
+ N_XI0/XI28/XI5/NET35_XI0/XI28/XI5/MM7_g N_VSS_XI0/XI28/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM8 N_XI0/XI28/XI5/NET35_XI0/XI28/XI5/MM8_d
+ N_WL<53>_XI0/XI28/XI5/MM8_g N_BLN<10>_XI0/XI28/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI5/MM5 N_XI0/XI28/XI5/NET34_XI0/XI28/XI5/MM5_d
+ N_XI0/XI28/XI5/NET33_XI0/XI28/XI5/MM5_g N_VDD_XI0/XI28/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI5/MM4 N_XI0/XI28/XI5/NET33_XI0/XI28/XI5/MM4_d
+ N_XI0/XI28/XI5/NET34_XI0/XI28/XI5/MM4_g N_VDD_XI0/XI28/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI5/MM10 N_XI0/XI28/XI5/NET35_XI0/XI28/XI5/MM10_d
+ N_XI0/XI28/XI5/NET36_XI0/XI28/XI5/MM10_g N_VDD_XI0/XI28/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI5/MM11 N_XI0/XI28/XI5/NET36_XI0/XI28/XI5/MM11_d
+ N_XI0/XI28/XI5/NET35_XI0/XI28/XI5/MM11_g N_VDD_XI0/XI28/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI6/MM2 N_XI0/XI28/XI6/NET34_XI0/XI28/XI6/MM2_d
+ N_XI0/XI28/XI6/NET33_XI0/XI28/XI6/MM2_g N_VSS_XI0/XI28/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM3 N_XI0/XI28/XI6/NET33_XI0/XI28/XI6/MM3_d
+ N_WL<52>_XI0/XI28/XI6/MM3_g N_BLN<9>_XI0/XI28/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM0 N_XI0/XI28/XI6/NET34_XI0/XI28/XI6/MM0_d
+ N_WL<52>_XI0/XI28/XI6/MM0_g N_BL<9>_XI0/XI28/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM1 N_XI0/XI28/XI6/NET33_XI0/XI28/XI6/MM1_d
+ N_XI0/XI28/XI6/NET34_XI0/XI28/XI6/MM1_g N_VSS_XI0/XI28/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM9 N_XI0/XI28/XI6/NET36_XI0/XI28/XI6/MM9_d
+ N_WL<53>_XI0/XI28/XI6/MM9_g N_BL<9>_XI0/XI28/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM6 N_XI0/XI28/XI6/NET35_XI0/XI28/XI6/MM6_d
+ N_XI0/XI28/XI6/NET36_XI0/XI28/XI6/MM6_g N_VSS_XI0/XI28/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM7 N_XI0/XI28/XI6/NET36_XI0/XI28/XI6/MM7_d
+ N_XI0/XI28/XI6/NET35_XI0/XI28/XI6/MM7_g N_VSS_XI0/XI28/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM8 N_XI0/XI28/XI6/NET35_XI0/XI28/XI6/MM8_d
+ N_WL<53>_XI0/XI28/XI6/MM8_g N_BLN<9>_XI0/XI28/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI6/MM5 N_XI0/XI28/XI6/NET34_XI0/XI28/XI6/MM5_d
+ N_XI0/XI28/XI6/NET33_XI0/XI28/XI6/MM5_g N_VDD_XI0/XI28/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI6/MM4 N_XI0/XI28/XI6/NET33_XI0/XI28/XI6/MM4_d
+ N_XI0/XI28/XI6/NET34_XI0/XI28/XI6/MM4_g N_VDD_XI0/XI28/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI6/MM10 N_XI0/XI28/XI6/NET35_XI0/XI28/XI6/MM10_d
+ N_XI0/XI28/XI6/NET36_XI0/XI28/XI6/MM10_g N_VDD_XI0/XI28/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI6/MM11 N_XI0/XI28/XI6/NET36_XI0/XI28/XI6/MM11_d
+ N_XI0/XI28/XI6/NET35_XI0/XI28/XI6/MM11_g N_VDD_XI0/XI28/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI7/MM2 N_XI0/XI28/XI7/NET34_XI0/XI28/XI7/MM2_d
+ N_XI0/XI28/XI7/NET33_XI0/XI28/XI7/MM2_g N_VSS_XI0/XI28/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM3 N_XI0/XI28/XI7/NET33_XI0/XI28/XI7/MM3_d
+ N_WL<52>_XI0/XI28/XI7/MM3_g N_BLN<8>_XI0/XI28/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM0 N_XI0/XI28/XI7/NET34_XI0/XI28/XI7/MM0_d
+ N_WL<52>_XI0/XI28/XI7/MM0_g N_BL<8>_XI0/XI28/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM1 N_XI0/XI28/XI7/NET33_XI0/XI28/XI7/MM1_d
+ N_XI0/XI28/XI7/NET34_XI0/XI28/XI7/MM1_g N_VSS_XI0/XI28/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM9 N_XI0/XI28/XI7/NET36_XI0/XI28/XI7/MM9_d
+ N_WL<53>_XI0/XI28/XI7/MM9_g N_BL<8>_XI0/XI28/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM6 N_XI0/XI28/XI7/NET35_XI0/XI28/XI7/MM6_d
+ N_XI0/XI28/XI7/NET36_XI0/XI28/XI7/MM6_g N_VSS_XI0/XI28/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM7 N_XI0/XI28/XI7/NET36_XI0/XI28/XI7/MM7_d
+ N_XI0/XI28/XI7/NET35_XI0/XI28/XI7/MM7_g N_VSS_XI0/XI28/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM8 N_XI0/XI28/XI7/NET35_XI0/XI28/XI7/MM8_d
+ N_WL<53>_XI0/XI28/XI7/MM8_g N_BLN<8>_XI0/XI28/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI7/MM5 N_XI0/XI28/XI7/NET34_XI0/XI28/XI7/MM5_d
+ N_XI0/XI28/XI7/NET33_XI0/XI28/XI7/MM5_g N_VDD_XI0/XI28/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI7/MM4 N_XI0/XI28/XI7/NET33_XI0/XI28/XI7/MM4_d
+ N_XI0/XI28/XI7/NET34_XI0/XI28/XI7/MM4_g N_VDD_XI0/XI28/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI7/MM10 N_XI0/XI28/XI7/NET35_XI0/XI28/XI7/MM10_d
+ N_XI0/XI28/XI7/NET36_XI0/XI28/XI7/MM10_g N_VDD_XI0/XI28/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI7/MM11 N_XI0/XI28/XI7/NET36_XI0/XI28/XI7/MM11_d
+ N_XI0/XI28/XI7/NET35_XI0/XI28/XI7/MM11_g N_VDD_XI0/XI28/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI8/MM2 N_XI0/XI28/XI8/NET34_XI0/XI28/XI8/MM2_d
+ N_XI0/XI28/XI8/NET33_XI0/XI28/XI8/MM2_g N_VSS_XI0/XI28/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM3 N_XI0/XI28/XI8/NET33_XI0/XI28/XI8/MM3_d
+ N_WL<52>_XI0/XI28/XI8/MM3_g N_BLN<7>_XI0/XI28/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM0 N_XI0/XI28/XI8/NET34_XI0/XI28/XI8/MM0_d
+ N_WL<52>_XI0/XI28/XI8/MM0_g N_BL<7>_XI0/XI28/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM1 N_XI0/XI28/XI8/NET33_XI0/XI28/XI8/MM1_d
+ N_XI0/XI28/XI8/NET34_XI0/XI28/XI8/MM1_g N_VSS_XI0/XI28/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM9 N_XI0/XI28/XI8/NET36_XI0/XI28/XI8/MM9_d
+ N_WL<53>_XI0/XI28/XI8/MM9_g N_BL<7>_XI0/XI28/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM6 N_XI0/XI28/XI8/NET35_XI0/XI28/XI8/MM6_d
+ N_XI0/XI28/XI8/NET36_XI0/XI28/XI8/MM6_g N_VSS_XI0/XI28/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM7 N_XI0/XI28/XI8/NET36_XI0/XI28/XI8/MM7_d
+ N_XI0/XI28/XI8/NET35_XI0/XI28/XI8/MM7_g N_VSS_XI0/XI28/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM8 N_XI0/XI28/XI8/NET35_XI0/XI28/XI8/MM8_d
+ N_WL<53>_XI0/XI28/XI8/MM8_g N_BLN<7>_XI0/XI28/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI8/MM5 N_XI0/XI28/XI8/NET34_XI0/XI28/XI8/MM5_d
+ N_XI0/XI28/XI8/NET33_XI0/XI28/XI8/MM5_g N_VDD_XI0/XI28/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI8/MM4 N_XI0/XI28/XI8/NET33_XI0/XI28/XI8/MM4_d
+ N_XI0/XI28/XI8/NET34_XI0/XI28/XI8/MM4_g N_VDD_XI0/XI28/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI8/MM10 N_XI0/XI28/XI8/NET35_XI0/XI28/XI8/MM10_d
+ N_XI0/XI28/XI8/NET36_XI0/XI28/XI8/MM10_g N_VDD_XI0/XI28/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI8/MM11 N_XI0/XI28/XI8/NET36_XI0/XI28/XI8/MM11_d
+ N_XI0/XI28/XI8/NET35_XI0/XI28/XI8/MM11_g N_VDD_XI0/XI28/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI9/MM2 N_XI0/XI28/XI9/NET34_XI0/XI28/XI9/MM2_d
+ N_XI0/XI28/XI9/NET33_XI0/XI28/XI9/MM2_g N_VSS_XI0/XI28/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM3 N_XI0/XI28/XI9/NET33_XI0/XI28/XI9/MM3_d
+ N_WL<52>_XI0/XI28/XI9/MM3_g N_BLN<6>_XI0/XI28/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM0 N_XI0/XI28/XI9/NET34_XI0/XI28/XI9/MM0_d
+ N_WL<52>_XI0/XI28/XI9/MM0_g N_BL<6>_XI0/XI28/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM1 N_XI0/XI28/XI9/NET33_XI0/XI28/XI9/MM1_d
+ N_XI0/XI28/XI9/NET34_XI0/XI28/XI9/MM1_g N_VSS_XI0/XI28/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM9 N_XI0/XI28/XI9/NET36_XI0/XI28/XI9/MM9_d
+ N_WL<53>_XI0/XI28/XI9/MM9_g N_BL<6>_XI0/XI28/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM6 N_XI0/XI28/XI9/NET35_XI0/XI28/XI9/MM6_d
+ N_XI0/XI28/XI9/NET36_XI0/XI28/XI9/MM6_g N_VSS_XI0/XI28/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM7 N_XI0/XI28/XI9/NET36_XI0/XI28/XI9/MM7_d
+ N_XI0/XI28/XI9/NET35_XI0/XI28/XI9/MM7_g N_VSS_XI0/XI28/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM8 N_XI0/XI28/XI9/NET35_XI0/XI28/XI9/MM8_d
+ N_WL<53>_XI0/XI28/XI9/MM8_g N_BLN<6>_XI0/XI28/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI9/MM5 N_XI0/XI28/XI9/NET34_XI0/XI28/XI9/MM5_d
+ N_XI0/XI28/XI9/NET33_XI0/XI28/XI9/MM5_g N_VDD_XI0/XI28/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI9/MM4 N_XI0/XI28/XI9/NET33_XI0/XI28/XI9/MM4_d
+ N_XI0/XI28/XI9/NET34_XI0/XI28/XI9/MM4_g N_VDD_XI0/XI28/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI9/MM10 N_XI0/XI28/XI9/NET35_XI0/XI28/XI9/MM10_d
+ N_XI0/XI28/XI9/NET36_XI0/XI28/XI9/MM10_g N_VDD_XI0/XI28/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI9/MM11 N_XI0/XI28/XI9/NET36_XI0/XI28/XI9/MM11_d
+ N_XI0/XI28/XI9/NET35_XI0/XI28/XI9/MM11_g N_VDD_XI0/XI28/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI10/MM2 N_XI0/XI28/XI10/NET34_XI0/XI28/XI10/MM2_d
+ N_XI0/XI28/XI10/NET33_XI0/XI28/XI10/MM2_g N_VSS_XI0/XI28/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM3 N_XI0/XI28/XI10/NET33_XI0/XI28/XI10/MM3_d
+ N_WL<52>_XI0/XI28/XI10/MM3_g N_BLN<5>_XI0/XI28/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM0 N_XI0/XI28/XI10/NET34_XI0/XI28/XI10/MM0_d
+ N_WL<52>_XI0/XI28/XI10/MM0_g N_BL<5>_XI0/XI28/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM1 N_XI0/XI28/XI10/NET33_XI0/XI28/XI10/MM1_d
+ N_XI0/XI28/XI10/NET34_XI0/XI28/XI10/MM1_g N_VSS_XI0/XI28/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM9 N_XI0/XI28/XI10/NET36_XI0/XI28/XI10/MM9_d
+ N_WL<53>_XI0/XI28/XI10/MM9_g N_BL<5>_XI0/XI28/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM6 N_XI0/XI28/XI10/NET35_XI0/XI28/XI10/MM6_d
+ N_XI0/XI28/XI10/NET36_XI0/XI28/XI10/MM6_g N_VSS_XI0/XI28/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM7 N_XI0/XI28/XI10/NET36_XI0/XI28/XI10/MM7_d
+ N_XI0/XI28/XI10/NET35_XI0/XI28/XI10/MM7_g N_VSS_XI0/XI28/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM8 N_XI0/XI28/XI10/NET35_XI0/XI28/XI10/MM8_d
+ N_WL<53>_XI0/XI28/XI10/MM8_g N_BLN<5>_XI0/XI28/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI10/MM5 N_XI0/XI28/XI10/NET34_XI0/XI28/XI10/MM5_d
+ N_XI0/XI28/XI10/NET33_XI0/XI28/XI10/MM5_g N_VDD_XI0/XI28/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI10/MM4 N_XI0/XI28/XI10/NET33_XI0/XI28/XI10/MM4_d
+ N_XI0/XI28/XI10/NET34_XI0/XI28/XI10/MM4_g N_VDD_XI0/XI28/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI10/MM10 N_XI0/XI28/XI10/NET35_XI0/XI28/XI10/MM10_d
+ N_XI0/XI28/XI10/NET36_XI0/XI28/XI10/MM10_g N_VDD_XI0/XI28/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI10/MM11 N_XI0/XI28/XI10/NET36_XI0/XI28/XI10/MM11_d
+ N_XI0/XI28/XI10/NET35_XI0/XI28/XI10/MM11_g N_VDD_XI0/XI28/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI11/MM2 N_XI0/XI28/XI11/NET34_XI0/XI28/XI11/MM2_d
+ N_XI0/XI28/XI11/NET33_XI0/XI28/XI11/MM2_g N_VSS_XI0/XI28/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM3 N_XI0/XI28/XI11/NET33_XI0/XI28/XI11/MM3_d
+ N_WL<52>_XI0/XI28/XI11/MM3_g N_BLN<4>_XI0/XI28/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM0 N_XI0/XI28/XI11/NET34_XI0/XI28/XI11/MM0_d
+ N_WL<52>_XI0/XI28/XI11/MM0_g N_BL<4>_XI0/XI28/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM1 N_XI0/XI28/XI11/NET33_XI0/XI28/XI11/MM1_d
+ N_XI0/XI28/XI11/NET34_XI0/XI28/XI11/MM1_g N_VSS_XI0/XI28/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM9 N_XI0/XI28/XI11/NET36_XI0/XI28/XI11/MM9_d
+ N_WL<53>_XI0/XI28/XI11/MM9_g N_BL<4>_XI0/XI28/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM6 N_XI0/XI28/XI11/NET35_XI0/XI28/XI11/MM6_d
+ N_XI0/XI28/XI11/NET36_XI0/XI28/XI11/MM6_g N_VSS_XI0/XI28/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM7 N_XI0/XI28/XI11/NET36_XI0/XI28/XI11/MM7_d
+ N_XI0/XI28/XI11/NET35_XI0/XI28/XI11/MM7_g N_VSS_XI0/XI28/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM8 N_XI0/XI28/XI11/NET35_XI0/XI28/XI11/MM8_d
+ N_WL<53>_XI0/XI28/XI11/MM8_g N_BLN<4>_XI0/XI28/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI11/MM5 N_XI0/XI28/XI11/NET34_XI0/XI28/XI11/MM5_d
+ N_XI0/XI28/XI11/NET33_XI0/XI28/XI11/MM5_g N_VDD_XI0/XI28/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI11/MM4 N_XI0/XI28/XI11/NET33_XI0/XI28/XI11/MM4_d
+ N_XI0/XI28/XI11/NET34_XI0/XI28/XI11/MM4_g N_VDD_XI0/XI28/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI11/MM10 N_XI0/XI28/XI11/NET35_XI0/XI28/XI11/MM10_d
+ N_XI0/XI28/XI11/NET36_XI0/XI28/XI11/MM10_g N_VDD_XI0/XI28/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI11/MM11 N_XI0/XI28/XI11/NET36_XI0/XI28/XI11/MM11_d
+ N_XI0/XI28/XI11/NET35_XI0/XI28/XI11/MM11_g N_VDD_XI0/XI28/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI12/MM2 N_XI0/XI28/XI12/NET34_XI0/XI28/XI12/MM2_d
+ N_XI0/XI28/XI12/NET33_XI0/XI28/XI12/MM2_g N_VSS_XI0/XI28/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM3 N_XI0/XI28/XI12/NET33_XI0/XI28/XI12/MM3_d
+ N_WL<52>_XI0/XI28/XI12/MM3_g N_BLN<3>_XI0/XI28/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM0 N_XI0/XI28/XI12/NET34_XI0/XI28/XI12/MM0_d
+ N_WL<52>_XI0/XI28/XI12/MM0_g N_BL<3>_XI0/XI28/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM1 N_XI0/XI28/XI12/NET33_XI0/XI28/XI12/MM1_d
+ N_XI0/XI28/XI12/NET34_XI0/XI28/XI12/MM1_g N_VSS_XI0/XI28/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM9 N_XI0/XI28/XI12/NET36_XI0/XI28/XI12/MM9_d
+ N_WL<53>_XI0/XI28/XI12/MM9_g N_BL<3>_XI0/XI28/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM6 N_XI0/XI28/XI12/NET35_XI0/XI28/XI12/MM6_d
+ N_XI0/XI28/XI12/NET36_XI0/XI28/XI12/MM6_g N_VSS_XI0/XI28/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM7 N_XI0/XI28/XI12/NET36_XI0/XI28/XI12/MM7_d
+ N_XI0/XI28/XI12/NET35_XI0/XI28/XI12/MM7_g N_VSS_XI0/XI28/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM8 N_XI0/XI28/XI12/NET35_XI0/XI28/XI12/MM8_d
+ N_WL<53>_XI0/XI28/XI12/MM8_g N_BLN<3>_XI0/XI28/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI12/MM5 N_XI0/XI28/XI12/NET34_XI0/XI28/XI12/MM5_d
+ N_XI0/XI28/XI12/NET33_XI0/XI28/XI12/MM5_g N_VDD_XI0/XI28/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI12/MM4 N_XI0/XI28/XI12/NET33_XI0/XI28/XI12/MM4_d
+ N_XI0/XI28/XI12/NET34_XI0/XI28/XI12/MM4_g N_VDD_XI0/XI28/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI12/MM10 N_XI0/XI28/XI12/NET35_XI0/XI28/XI12/MM10_d
+ N_XI0/XI28/XI12/NET36_XI0/XI28/XI12/MM10_g N_VDD_XI0/XI28/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI12/MM11 N_XI0/XI28/XI12/NET36_XI0/XI28/XI12/MM11_d
+ N_XI0/XI28/XI12/NET35_XI0/XI28/XI12/MM11_g N_VDD_XI0/XI28/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI13/MM2 N_XI0/XI28/XI13/NET34_XI0/XI28/XI13/MM2_d
+ N_XI0/XI28/XI13/NET33_XI0/XI28/XI13/MM2_g N_VSS_XI0/XI28/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM3 N_XI0/XI28/XI13/NET33_XI0/XI28/XI13/MM3_d
+ N_WL<52>_XI0/XI28/XI13/MM3_g N_BLN<2>_XI0/XI28/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM0 N_XI0/XI28/XI13/NET34_XI0/XI28/XI13/MM0_d
+ N_WL<52>_XI0/XI28/XI13/MM0_g N_BL<2>_XI0/XI28/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM1 N_XI0/XI28/XI13/NET33_XI0/XI28/XI13/MM1_d
+ N_XI0/XI28/XI13/NET34_XI0/XI28/XI13/MM1_g N_VSS_XI0/XI28/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM9 N_XI0/XI28/XI13/NET36_XI0/XI28/XI13/MM9_d
+ N_WL<53>_XI0/XI28/XI13/MM9_g N_BL<2>_XI0/XI28/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM6 N_XI0/XI28/XI13/NET35_XI0/XI28/XI13/MM6_d
+ N_XI0/XI28/XI13/NET36_XI0/XI28/XI13/MM6_g N_VSS_XI0/XI28/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM7 N_XI0/XI28/XI13/NET36_XI0/XI28/XI13/MM7_d
+ N_XI0/XI28/XI13/NET35_XI0/XI28/XI13/MM7_g N_VSS_XI0/XI28/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM8 N_XI0/XI28/XI13/NET35_XI0/XI28/XI13/MM8_d
+ N_WL<53>_XI0/XI28/XI13/MM8_g N_BLN<2>_XI0/XI28/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI13/MM5 N_XI0/XI28/XI13/NET34_XI0/XI28/XI13/MM5_d
+ N_XI0/XI28/XI13/NET33_XI0/XI28/XI13/MM5_g N_VDD_XI0/XI28/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI13/MM4 N_XI0/XI28/XI13/NET33_XI0/XI28/XI13/MM4_d
+ N_XI0/XI28/XI13/NET34_XI0/XI28/XI13/MM4_g N_VDD_XI0/XI28/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI13/MM10 N_XI0/XI28/XI13/NET35_XI0/XI28/XI13/MM10_d
+ N_XI0/XI28/XI13/NET36_XI0/XI28/XI13/MM10_g N_VDD_XI0/XI28/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI13/MM11 N_XI0/XI28/XI13/NET36_XI0/XI28/XI13/MM11_d
+ N_XI0/XI28/XI13/NET35_XI0/XI28/XI13/MM11_g N_VDD_XI0/XI28/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI14/MM2 N_XI0/XI28/XI14/NET34_XI0/XI28/XI14/MM2_d
+ N_XI0/XI28/XI14/NET33_XI0/XI28/XI14/MM2_g N_VSS_XI0/XI28/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM3 N_XI0/XI28/XI14/NET33_XI0/XI28/XI14/MM3_d
+ N_WL<52>_XI0/XI28/XI14/MM3_g N_BLN<1>_XI0/XI28/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM0 N_XI0/XI28/XI14/NET34_XI0/XI28/XI14/MM0_d
+ N_WL<52>_XI0/XI28/XI14/MM0_g N_BL<1>_XI0/XI28/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM1 N_XI0/XI28/XI14/NET33_XI0/XI28/XI14/MM1_d
+ N_XI0/XI28/XI14/NET34_XI0/XI28/XI14/MM1_g N_VSS_XI0/XI28/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM9 N_XI0/XI28/XI14/NET36_XI0/XI28/XI14/MM9_d
+ N_WL<53>_XI0/XI28/XI14/MM9_g N_BL<1>_XI0/XI28/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM6 N_XI0/XI28/XI14/NET35_XI0/XI28/XI14/MM6_d
+ N_XI0/XI28/XI14/NET36_XI0/XI28/XI14/MM6_g N_VSS_XI0/XI28/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM7 N_XI0/XI28/XI14/NET36_XI0/XI28/XI14/MM7_d
+ N_XI0/XI28/XI14/NET35_XI0/XI28/XI14/MM7_g N_VSS_XI0/XI28/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM8 N_XI0/XI28/XI14/NET35_XI0/XI28/XI14/MM8_d
+ N_WL<53>_XI0/XI28/XI14/MM8_g N_BLN<1>_XI0/XI28/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI14/MM5 N_XI0/XI28/XI14/NET34_XI0/XI28/XI14/MM5_d
+ N_XI0/XI28/XI14/NET33_XI0/XI28/XI14/MM5_g N_VDD_XI0/XI28/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI14/MM4 N_XI0/XI28/XI14/NET33_XI0/XI28/XI14/MM4_d
+ N_XI0/XI28/XI14/NET34_XI0/XI28/XI14/MM4_g N_VDD_XI0/XI28/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI14/MM10 N_XI0/XI28/XI14/NET35_XI0/XI28/XI14/MM10_d
+ N_XI0/XI28/XI14/NET36_XI0/XI28/XI14/MM10_g N_VDD_XI0/XI28/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI14/MM11 N_XI0/XI28/XI14/NET36_XI0/XI28/XI14/MM11_d
+ N_XI0/XI28/XI14/NET35_XI0/XI28/XI14/MM11_g N_VDD_XI0/XI28/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI15/MM2 N_XI0/XI28/XI15/NET34_XI0/XI28/XI15/MM2_d
+ N_XI0/XI28/XI15/NET33_XI0/XI28/XI15/MM2_g N_VSS_XI0/XI28/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM3 N_XI0/XI28/XI15/NET33_XI0/XI28/XI15/MM3_d
+ N_WL<52>_XI0/XI28/XI15/MM3_g N_BLN<0>_XI0/XI28/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM0 N_XI0/XI28/XI15/NET34_XI0/XI28/XI15/MM0_d
+ N_WL<52>_XI0/XI28/XI15/MM0_g N_BL<0>_XI0/XI28/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM1 N_XI0/XI28/XI15/NET33_XI0/XI28/XI15/MM1_d
+ N_XI0/XI28/XI15/NET34_XI0/XI28/XI15/MM1_g N_VSS_XI0/XI28/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM9 N_XI0/XI28/XI15/NET36_XI0/XI28/XI15/MM9_d
+ N_WL<53>_XI0/XI28/XI15/MM9_g N_BL<0>_XI0/XI28/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM6 N_XI0/XI28/XI15/NET35_XI0/XI28/XI15/MM6_d
+ N_XI0/XI28/XI15/NET36_XI0/XI28/XI15/MM6_g N_VSS_XI0/XI28/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM7 N_XI0/XI28/XI15/NET36_XI0/XI28/XI15/MM7_d
+ N_XI0/XI28/XI15/NET35_XI0/XI28/XI15/MM7_g N_VSS_XI0/XI28/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM8 N_XI0/XI28/XI15/NET35_XI0/XI28/XI15/MM8_d
+ N_WL<53>_XI0/XI28/XI15/MM8_g N_BLN<0>_XI0/XI28/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI28/XI15/MM5 N_XI0/XI28/XI15/NET34_XI0/XI28/XI15/MM5_d
+ N_XI0/XI28/XI15/NET33_XI0/XI28/XI15/MM5_g N_VDD_XI0/XI28/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI15/MM4 N_XI0/XI28/XI15/NET33_XI0/XI28/XI15/MM4_d
+ N_XI0/XI28/XI15/NET34_XI0/XI28/XI15/MM4_g N_VDD_XI0/XI28/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI15/MM10 N_XI0/XI28/XI15/NET35_XI0/XI28/XI15/MM10_d
+ N_XI0/XI28/XI15/NET36_XI0/XI28/XI15/MM10_g N_VDD_XI0/XI28/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI28/XI15/MM11 N_XI0/XI28/XI15/NET36_XI0/XI28/XI15/MM11_d
+ N_XI0/XI28/XI15/NET35_XI0/XI28/XI15/MM11_g N_VDD_XI0/XI28/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI0/MM2 N_XI0/XI29/XI0/NET34_XI0/XI29/XI0/MM2_d
+ N_XI0/XI29/XI0/NET33_XI0/XI29/XI0/MM2_g N_VSS_XI0/XI29/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM3 N_XI0/XI29/XI0/NET33_XI0/XI29/XI0/MM3_d
+ N_WL<54>_XI0/XI29/XI0/MM3_g N_BLN<15>_XI0/XI29/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM0 N_XI0/XI29/XI0/NET34_XI0/XI29/XI0/MM0_d
+ N_WL<54>_XI0/XI29/XI0/MM0_g N_BL<15>_XI0/XI29/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM1 N_XI0/XI29/XI0/NET33_XI0/XI29/XI0/MM1_d
+ N_XI0/XI29/XI0/NET34_XI0/XI29/XI0/MM1_g N_VSS_XI0/XI29/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM9 N_XI0/XI29/XI0/NET36_XI0/XI29/XI0/MM9_d
+ N_WL<55>_XI0/XI29/XI0/MM9_g N_BL<15>_XI0/XI29/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM6 N_XI0/XI29/XI0/NET35_XI0/XI29/XI0/MM6_d
+ N_XI0/XI29/XI0/NET36_XI0/XI29/XI0/MM6_g N_VSS_XI0/XI29/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM7 N_XI0/XI29/XI0/NET36_XI0/XI29/XI0/MM7_d
+ N_XI0/XI29/XI0/NET35_XI0/XI29/XI0/MM7_g N_VSS_XI0/XI29/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM8 N_XI0/XI29/XI0/NET35_XI0/XI29/XI0/MM8_d
+ N_WL<55>_XI0/XI29/XI0/MM8_g N_BLN<15>_XI0/XI29/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI0/MM5 N_XI0/XI29/XI0/NET34_XI0/XI29/XI0/MM5_d
+ N_XI0/XI29/XI0/NET33_XI0/XI29/XI0/MM5_g N_VDD_XI0/XI29/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI0/MM4 N_XI0/XI29/XI0/NET33_XI0/XI29/XI0/MM4_d
+ N_XI0/XI29/XI0/NET34_XI0/XI29/XI0/MM4_g N_VDD_XI0/XI29/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI0/MM10 N_XI0/XI29/XI0/NET35_XI0/XI29/XI0/MM10_d
+ N_XI0/XI29/XI0/NET36_XI0/XI29/XI0/MM10_g N_VDD_XI0/XI29/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI0/MM11 N_XI0/XI29/XI0/NET36_XI0/XI29/XI0/MM11_d
+ N_XI0/XI29/XI0/NET35_XI0/XI29/XI0/MM11_g N_VDD_XI0/XI29/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI1/MM2 N_XI0/XI29/XI1/NET34_XI0/XI29/XI1/MM2_d
+ N_XI0/XI29/XI1/NET33_XI0/XI29/XI1/MM2_g N_VSS_XI0/XI29/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM3 N_XI0/XI29/XI1/NET33_XI0/XI29/XI1/MM3_d
+ N_WL<54>_XI0/XI29/XI1/MM3_g N_BLN<14>_XI0/XI29/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM0 N_XI0/XI29/XI1/NET34_XI0/XI29/XI1/MM0_d
+ N_WL<54>_XI0/XI29/XI1/MM0_g N_BL<14>_XI0/XI29/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM1 N_XI0/XI29/XI1/NET33_XI0/XI29/XI1/MM1_d
+ N_XI0/XI29/XI1/NET34_XI0/XI29/XI1/MM1_g N_VSS_XI0/XI29/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM9 N_XI0/XI29/XI1/NET36_XI0/XI29/XI1/MM9_d
+ N_WL<55>_XI0/XI29/XI1/MM9_g N_BL<14>_XI0/XI29/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM6 N_XI0/XI29/XI1/NET35_XI0/XI29/XI1/MM6_d
+ N_XI0/XI29/XI1/NET36_XI0/XI29/XI1/MM6_g N_VSS_XI0/XI29/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM7 N_XI0/XI29/XI1/NET36_XI0/XI29/XI1/MM7_d
+ N_XI0/XI29/XI1/NET35_XI0/XI29/XI1/MM7_g N_VSS_XI0/XI29/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM8 N_XI0/XI29/XI1/NET35_XI0/XI29/XI1/MM8_d
+ N_WL<55>_XI0/XI29/XI1/MM8_g N_BLN<14>_XI0/XI29/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI1/MM5 N_XI0/XI29/XI1/NET34_XI0/XI29/XI1/MM5_d
+ N_XI0/XI29/XI1/NET33_XI0/XI29/XI1/MM5_g N_VDD_XI0/XI29/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI1/MM4 N_XI0/XI29/XI1/NET33_XI0/XI29/XI1/MM4_d
+ N_XI0/XI29/XI1/NET34_XI0/XI29/XI1/MM4_g N_VDD_XI0/XI29/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI1/MM10 N_XI0/XI29/XI1/NET35_XI0/XI29/XI1/MM10_d
+ N_XI0/XI29/XI1/NET36_XI0/XI29/XI1/MM10_g N_VDD_XI0/XI29/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI1/MM11 N_XI0/XI29/XI1/NET36_XI0/XI29/XI1/MM11_d
+ N_XI0/XI29/XI1/NET35_XI0/XI29/XI1/MM11_g N_VDD_XI0/XI29/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI2/MM2 N_XI0/XI29/XI2/NET34_XI0/XI29/XI2/MM2_d
+ N_XI0/XI29/XI2/NET33_XI0/XI29/XI2/MM2_g N_VSS_XI0/XI29/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM3 N_XI0/XI29/XI2/NET33_XI0/XI29/XI2/MM3_d
+ N_WL<54>_XI0/XI29/XI2/MM3_g N_BLN<13>_XI0/XI29/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM0 N_XI0/XI29/XI2/NET34_XI0/XI29/XI2/MM0_d
+ N_WL<54>_XI0/XI29/XI2/MM0_g N_BL<13>_XI0/XI29/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM1 N_XI0/XI29/XI2/NET33_XI0/XI29/XI2/MM1_d
+ N_XI0/XI29/XI2/NET34_XI0/XI29/XI2/MM1_g N_VSS_XI0/XI29/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM9 N_XI0/XI29/XI2/NET36_XI0/XI29/XI2/MM9_d
+ N_WL<55>_XI0/XI29/XI2/MM9_g N_BL<13>_XI0/XI29/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM6 N_XI0/XI29/XI2/NET35_XI0/XI29/XI2/MM6_d
+ N_XI0/XI29/XI2/NET36_XI0/XI29/XI2/MM6_g N_VSS_XI0/XI29/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM7 N_XI0/XI29/XI2/NET36_XI0/XI29/XI2/MM7_d
+ N_XI0/XI29/XI2/NET35_XI0/XI29/XI2/MM7_g N_VSS_XI0/XI29/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM8 N_XI0/XI29/XI2/NET35_XI0/XI29/XI2/MM8_d
+ N_WL<55>_XI0/XI29/XI2/MM8_g N_BLN<13>_XI0/XI29/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI2/MM5 N_XI0/XI29/XI2/NET34_XI0/XI29/XI2/MM5_d
+ N_XI0/XI29/XI2/NET33_XI0/XI29/XI2/MM5_g N_VDD_XI0/XI29/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI2/MM4 N_XI0/XI29/XI2/NET33_XI0/XI29/XI2/MM4_d
+ N_XI0/XI29/XI2/NET34_XI0/XI29/XI2/MM4_g N_VDD_XI0/XI29/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI2/MM10 N_XI0/XI29/XI2/NET35_XI0/XI29/XI2/MM10_d
+ N_XI0/XI29/XI2/NET36_XI0/XI29/XI2/MM10_g N_VDD_XI0/XI29/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI2/MM11 N_XI0/XI29/XI2/NET36_XI0/XI29/XI2/MM11_d
+ N_XI0/XI29/XI2/NET35_XI0/XI29/XI2/MM11_g N_VDD_XI0/XI29/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI3/MM2 N_XI0/XI29/XI3/NET34_XI0/XI29/XI3/MM2_d
+ N_XI0/XI29/XI3/NET33_XI0/XI29/XI3/MM2_g N_VSS_XI0/XI29/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM3 N_XI0/XI29/XI3/NET33_XI0/XI29/XI3/MM3_d
+ N_WL<54>_XI0/XI29/XI3/MM3_g N_BLN<12>_XI0/XI29/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM0 N_XI0/XI29/XI3/NET34_XI0/XI29/XI3/MM0_d
+ N_WL<54>_XI0/XI29/XI3/MM0_g N_BL<12>_XI0/XI29/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM1 N_XI0/XI29/XI3/NET33_XI0/XI29/XI3/MM1_d
+ N_XI0/XI29/XI3/NET34_XI0/XI29/XI3/MM1_g N_VSS_XI0/XI29/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM9 N_XI0/XI29/XI3/NET36_XI0/XI29/XI3/MM9_d
+ N_WL<55>_XI0/XI29/XI3/MM9_g N_BL<12>_XI0/XI29/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM6 N_XI0/XI29/XI3/NET35_XI0/XI29/XI3/MM6_d
+ N_XI0/XI29/XI3/NET36_XI0/XI29/XI3/MM6_g N_VSS_XI0/XI29/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM7 N_XI0/XI29/XI3/NET36_XI0/XI29/XI3/MM7_d
+ N_XI0/XI29/XI3/NET35_XI0/XI29/XI3/MM7_g N_VSS_XI0/XI29/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM8 N_XI0/XI29/XI3/NET35_XI0/XI29/XI3/MM8_d
+ N_WL<55>_XI0/XI29/XI3/MM8_g N_BLN<12>_XI0/XI29/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI3/MM5 N_XI0/XI29/XI3/NET34_XI0/XI29/XI3/MM5_d
+ N_XI0/XI29/XI3/NET33_XI0/XI29/XI3/MM5_g N_VDD_XI0/XI29/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI3/MM4 N_XI0/XI29/XI3/NET33_XI0/XI29/XI3/MM4_d
+ N_XI0/XI29/XI3/NET34_XI0/XI29/XI3/MM4_g N_VDD_XI0/XI29/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI3/MM10 N_XI0/XI29/XI3/NET35_XI0/XI29/XI3/MM10_d
+ N_XI0/XI29/XI3/NET36_XI0/XI29/XI3/MM10_g N_VDD_XI0/XI29/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI3/MM11 N_XI0/XI29/XI3/NET36_XI0/XI29/XI3/MM11_d
+ N_XI0/XI29/XI3/NET35_XI0/XI29/XI3/MM11_g N_VDD_XI0/XI29/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI4/MM2 N_XI0/XI29/XI4/NET34_XI0/XI29/XI4/MM2_d
+ N_XI0/XI29/XI4/NET33_XI0/XI29/XI4/MM2_g N_VSS_XI0/XI29/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM3 N_XI0/XI29/XI4/NET33_XI0/XI29/XI4/MM3_d
+ N_WL<54>_XI0/XI29/XI4/MM3_g N_BLN<11>_XI0/XI29/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM0 N_XI0/XI29/XI4/NET34_XI0/XI29/XI4/MM0_d
+ N_WL<54>_XI0/XI29/XI4/MM0_g N_BL<11>_XI0/XI29/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM1 N_XI0/XI29/XI4/NET33_XI0/XI29/XI4/MM1_d
+ N_XI0/XI29/XI4/NET34_XI0/XI29/XI4/MM1_g N_VSS_XI0/XI29/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM9 N_XI0/XI29/XI4/NET36_XI0/XI29/XI4/MM9_d
+ N_WL<55>_XI0/XI29/XI4/MM9_g N_BL<11>_XI0/XI29/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM6 N_XI0/XI29/XI4/NET35_XI0/XI29/XI4/MM6_d
+ N_XI0/XI29/XI4/NET36_XI0/XI29/XI4/MM6_g N_VSS_XI0/XI29/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM7 N_XI0/XI29/XI4/NET36_XI0/XI29/XI4/MM7_d
+ N_XI0/XI29/XI4/NET35_XI0/XI29/XI4/MM7_g N_VSS_XI0/XI29/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM8 N_XI0/XI29/XI4/NET35_XI0/XI29/XI4/MM8_d
+ N_WL<55>_XI0/XI29/XI4/MM8_g N_BLN<11>_XI0/XI29/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI4/MM5 N_XI0/XI29/XI4/NET34_XI0/XI29/XI4/MM5_d
+ N_XI0/XI29/XI4/NET33_XI0/XI29/XI4/MM5_g N_VDD_XI0/XI29/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI4/MM4 N_XI0/XI29/XI4/NET33_XI0/XI29/XI4/MM4_d
+ N_XI0/XI29/XI4/NET34_XI0/XI29/XI4/MM4_g N_VDD_XI0/XI29/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI4/MM10 N_XI0/XI29/XI4/NET35_XI0/XI29/XI4/MM10_d
+ N_XI0/XI29/XI4/NET36_XI0/XI29/XI4/MM10_g N_VDD_XI0/XI29/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI4/MM11 N_XI0/XI29/XI4/NET36_XI0/XI29/XI4/MM11_d
+ N_XI0/XI29/XI4/NET35_XI0/XI29/XI4/MM11_g N_VDD_XI0/XI29/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI5/MM2 N_XI0/XI29/XI5/NET34_XI0/XI29/XI5/MM2_d
+ N_XI0/XI29/XI5/NET33_XI0/XI29/XI5/MM2_g N_VSS_XI0/XI29/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM3 N_XI0/XI29/XI5/NET33_XI0/XI29/XI5/MM3_d
+ N_WL<54>_XI0/XI29/XI5/MM3_g N_BLN<10>_XI0/XI29/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM0 N_XI0/XI29/XI5/NET34_XI0/XI29/XI5/MM0_d
+ N_WL<54>_XI0/XI29/XI5/MM0_g N_BL<10>_XI0/XI29/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM1 N_XI0/XI29/XI5/NET33_XI0/XI29/XI5/MM1_d
+ N_XI0/XI29/XI5/NET34_XI0/XI29/XI5/MM1_g N_VSS_XI0/XI29/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM9 N_XI0/XI29/XI5/NET36_XI0/XI29/XI5/MM9_d
+ N_WL<55>_XI0/XI29/XI5/MM9_g N_BL<10>_XI0/XI29/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM6 N_XI0/XI29/XI5/NET35_XI0/XI29/XI5/MM6_d
+ N_XI0/XI29/XI5/NET36_XI0/XI29/XI5/MM6_g N_VSS_XI0/XI29/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM7 N_XI0/XI29/XI5/NET36_XI0/XI29/XI5/MM7_d
+ N_XI0/XI29/XI5/NET35_XI0/XI29/XI5/MM7_g N_VSS_XI0/XI29/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM8 N_XI0/XI29/XI5/NET35_XI0/XI29/XI5/MM8_d
+ N_WL<55>_XI0/XI29/XI5/MM8_g N_BLN<10>_XI0/XI29/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI5/MM5 N_XI0/XI29/XI5/NET34_XI0/XI29/XI5/MM5_d
+ N_XI0/XI29/XI5/NET33_XI0/XI29/XI5/MM5_g N_VDD_XI0/XI29/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI5/MM4 N_XI0/XI29/XI5/NET33_XI0/XI29/XI5/MM4_d
+ N_XI0/XI29/XI5/NET34_XI0/XI29/XI5/MM4_g N_VDD_XI0/XI29/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI5/MM10 N_XI0/XI29/XI5/NET35_XI0/XI29/XI5/MM10_d
+ N_XI0/XI29/XI5/NET36_XI0/XI29/XI5/MM10_g N_VDD_XI0/XI29/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI5/MM11 N_XI0/XI29/XI5/NET36_XI0/XI29/XI5/MM11_d
+ N_XI0/XI29/XI5/NET35_XI0/XI29/XI5/MM11_g N_VDD_XI0/XI29/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI6/MM2 N_XI0/XI29/XI6/NET34_XI0/XI29/XI6/MM2_d
+ N_XI0/XI29/XI6/NET33_XI0/XI29/XI6/MM2_g N_VSS_XI0/XI29/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM3 N_XI0/XI29/XI6/NET33_XI0/XI29/XI6/MM3_d
+ N_WL<54>_XI0/XI29/XI6/MM3_g N_BLN<9>_XI0/XI29/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM0 N_XI0/XI29/XI6/NET34_XI0/XI29/XI6/MM0_d
+ N_WL<54>_XI0/XI29/XI6/MM0_g N_BL<9>_XI0/XI29/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM1 N_XI0/XI29/XI6/NET33_XI0/XI29/XI6/MM1_d
+ N_XI0/XI29/XI6/NET34_XI0/XI29/XI6/MM1_g N_VSS_XI0/XI29/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM9 N_XI0/XI29/XI6/NET36_XI0/XI29/XI6/MM9_d
+ N_WL<55>_XI0/XI29/XI6/MM9_g N_BL<9>_XI0/XI29/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM6 N_XI0/XI29/XI6/NET35_XI0/XI29/XI6/MM6_d
+ N_XI0/XI29/XI6/NET36_XI0/XI29/XI6/MM6_g N_VSS_XI0/XI29/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM7 N_XI0/XI29/XI6/NET36_XI0/XI29/XI6/MM7_d
+ N_XI0/XI29/XI6/NET35_XI0/XI29/XI6/MM7_g N_VSS_XI0/XI29/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM8 N_XI0/XI29/XI6/NET35_XI0/XI29/XI6/MM8_d
+ N_WL<55>_XI0/XI29/XI6/MM8_g N_BLN<9>_XI0/XI29/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI6/MM5 N_XI0/XI29/XI6/NET34_XI0/XI29/XI6/MM5_d
+ N_XI0/XI29/XI6/NET33_XI0/XI29/XI6/MM5_g N_VDD_XI0/XI29/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI6/MM4 N_XI0/XI29/XI6/NET33_XI0/XI29/XI6/MM4_d
+ N_XI0/XI29/XI6/NET34_XI0/XI29/XI6/MM4_g N_VDD_XI0/XI29/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI6/MM10 N_XI0/XI29/XI6/NET35_XI0/XI29/XI6/MM10_d
+ N_XI0/XI29/XI6/NET36_XI0/XI29/XI6/MM10_g N_VDD_XI0/XI29/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI6/MM11 N_XI0/XI29/XI6/NET36_XI0/XI29/XI6/MM11_d
+ N_XI0/XI29/XI6/NET35_XI0/XI29/XI6/MM11_g N_VDD_XI0/XI29/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI7/MM2 N_XI0/XI29/XI7/NET34_XI0/XI29/XI7/MM2_d
+ N_XI0/XI29/XI7/NET33_XI0/XI29/XI7/MM2_g N_VSS_XI0/XI29/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM3 N_XI0/XI29/XI7/NET33_XI0/XI29/XI7/MM3_d
+ N_WL<54>_XI0/XI29/XI7/MM3_g N_BLN<8>_XI0/XI29/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM0 N_XI0/XI29/XI7/NET34_XI0/XI29/XI7/MM0_d
+ N_WL<54>_XI0/XI29/XI7/MM0_g N_BL<8>_XI0/XI29/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM1 N_XI0/XI29/XI7/NET33_XI0/XI29/XI7/MM1_d
+ N_XI0/XI29/XI7/NET34_XI0/XI29/XI7/MM1_g N_VSS_XI0/XI29/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM9 N_XI0/XI29/XI7/NET36_XI0/XI29/XI7/MM9_d
+ N_WL<55>_XI0/XI29/XI7/MM9_g N_BL<8>_XI0/XI29/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM6 N_XI0/XI29/XI7/NET35_XI0/XI29/XI7/MM6_d
+ N_XI0/XI29/XI7/NET36_XI0/XI29/XI7/MM6_g N_VSS_XI0/XI29/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM7 N_XI0/XI29/XI7/NET36_XI0/XI29/XI7/MM7_d
+ N_XI0/XI29/XI7/NET35_XI0/XI29/XI7/MM7_g N_VSS_XI0/XI29/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM8 N_XI0/XI29/XI7/NET35_XI0/XI29/XI7/MM8_d
+ N_WL<55>_XI0/XI29/XI7/MM8_g N_BLN<8>_XI0/XI29/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI7/MM5 N_XI0/XI29/XI7/NET34_XI0/XI29/XI7/MM5_d
+ N_XI0/XI29/XI7/NET33_XI0/XI29/XI7/MM5_g N_VDD_XI0/XI29/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI7/MM4 N_XI0/XI29/XI7/NET33_XI0/XI29/XI7/MM4_d
+ N_XI0/XI29/XI7/NET34_XI0/XI29/XI7/MM4_g N_VDD_XI0/XI29/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI7/MM10 N_XI0/XI29/XI7/NET35_XI0/XI29/XI7/MM10_d
+ N_XI0/XI29/XI7/NET36_XI0/XI29/XI7/MM10_g N_VDD_XI0/XI29/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI7/MM11 N_XI0/XI29/XI7/NET36_XI0/XI29/XI7/MM11_d
+ N_XI0/XI29/XI7/NET35_XI0/XI29/XI7/MM11_g N_VDD_XI0/XI29/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI8/MM2 N_XI0/XI29/XI8/NET34_XI0/XI29/XI8/MM2_d
+ N_XI0/XI29/XI8/NET33_XI0/XI29/XI8/MM2_g N_VSS_XI0/XI29/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM3 N_XI0/XI29/XI8/NET33_XI0/XI29/XI8/MM3_d
+ N_WL<54>_XI0/XI29/XI8/MM3_g N_BLN<7>_XI0/XI29/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM0 N_XI0/XI29/XI8/NET34_XI0/XI29/XI8/MM0_d
+ N_WL<54>_XI0/XI29/XI8/MM0_g N_BL<7>_XI0/XI29/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM1 N_XI0/XI29/XI8/NET33_XI0/XI29/XI8/MM1_d
+ N_XI0/XI29/XI8/NET34_XI0/XI29/XI8/MM1_g N_VSS_XI0/XI29/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM9 N_XI0/XI29/XI8/NET36_XI0/XI29/XI8/MM9_d
+ N_WL<55>_XI0/XI29/XI8/MM9_g N_BL<7>_XI0/XI29/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM6 N_XI0/XI29/XI8/NET35_XI0/XI29/XI8/MM6_d
+ N_XI0/XI29/XI8/NET36_XI0/XI29/XI8/MM6_g N_VSS_XI0/XI29/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM7 N_XI0/XI29/XI8/NET36_XI0/XI29/XI8/MM7_d
+ N_XI0/XI29/XI8/NET35_XI0/XI29/XI8/MM7_g N_VSS_XI0/XI29/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM8 N_XI0/XI29/XI8/NET35_XI0/XI29/XI8/MM8_d
+ N_WL<55>_XI0/XI29/XI8/MM8_g N_BLN<7>_XI0/XI29/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI8/MM5 N_XI0/XI29/XI8/NET34_XI0/XI29/XI8/MM5_d
+ N_XI0/XI29/XI8/NET33_XI0/XI29/XI8/MM5_g N_VDD_XI0/XI29/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI8/MM4 N_XI0/XI29/XI8/NET33_XI0/XI29/XI8/MM4_d
+ N_XI0/XI29/XI8/NET34_XI0/XI29/XI8/MM4_g N_VDD_XI0/XI29/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI8/MM10 N_XI0/XI29/XI8/NET35_XI0/XI29/XI8/MM10_d
+ N_XI0/XI29/XI8/NET36_XI0/XI29/XI8/MM10_g N_VDD_XI0/XI29/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI8/MM11 N_XI0/XI29/XI8/NET36_XI0/XI29/XI8/MM11_d
+ N_XI0/XI29/XI8/NET35_XI0/XI29/XI8/MM11_g N_VDD_XI0/XI29/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI9/MM2 N_XI0/XI29/XI9/NET34_XI0/XI29/XI9/MM2_d
+ N_XI0/XI29/XI9/NET33_XI0/XI29/XI9/MM2_g N_VSS_XI0/XI29/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM3 N_XI0/XI29/XI9/NET33_XI0/XI29/XI9/MM3_d
+ N_WL<54>_XI0/XI29/XI9/MM3_g N_BLN<6>_XI0/XI29/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM0 N_XI0/XI29/XI9/NET34_XI0/XI29/XI9/MM0_d
+ N_WL<54>_XI0/XI29/XI9/MM0_g N_BL<6>_XI0/XI29/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM1 N_XI0/XI29/XI9/NET33_XI0/XI29/XI9/MM1_d
+ N_XI0/XI29/XI9/NET34_XI0/XI29/XI9/MM1_g N_VSS_XI0/XI29/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM9 N_XI0/XI29/XI9/NET36_XI0/XI29/XI9/MM9_d
+ N_WL<55>_XI0/XI29/XI9/MM9_g N_BL<6>_XI0/XI29/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM6 N_XI0/XI29/XI9/NET35_XI0/XI29/XI9/MM6_d
+ N_XI0/XI29/XI9/NET36_XI0/XI29/XI9/MM6_g N_VSS_XI0/XI29/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM7 N_XI0/XI29/XI9/NET36_XI0/XI29/XI9/MM7_d
+ N_XI0/XI29/XI9/NET35_XI0/XI29/XI9/MM7_g N_VSS_XI0/XI29/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM8 N_XI0/XI29/XI9/NET35_XI0/XI29/XI9/MM8_d
+ N_WL<55>_XI0/XI29/XI9/MM8_g N_BLN<6>_XI0/XI29/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI9/MM5 N_XI0/XI29/XI9/NET34_XI0/XI29/XI9/MM5_d
+ N_XI0/XI29/XI9/NET33_XI0/XI29/XI9/MM5_g N_VDD_XI0/XI29/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI9/MM4 N_XI0/XI29/XI9/NET33_XI0/XI29/XI9/MM4_d
+ N_XI0/XI29/XI9/NET34_XI0/XI29/XI9/MM4_g N_VDD_XI0/XI29/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI9/MM10 N_XI0/XI29/XI9/NET35_XI0/XI29/XI9/MM10_d
+ N_XI0/XI29/XI9/NET36_XI0/XI29/XI9/MM10_g N_VDD_XI0/XI29/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI9/MM11 N_XI0/XI29/XI9/NET36_XI0/XI29/XI9/MM11_d
+ N_XI0/XI29/XI9/NET35_XI0/XI29/XI9/MM11_g N_VDD_XI0/XI29/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI10/MM2 N_XI0/XI29/XI10/NET34_XI0/XI29/XI10/MM2_d
+ N_XI0/XI29/XI10/NET33_XI0/XI29/XI10/MM2_g N_VSS_XI0/XI29/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM3 N_XI0/XI29/XI10/NET33_XI0/XI29/XI10/MM3_d
+ N_WL<54>_XI0/XI29/XI10/MM3_g N_BLN<5>_XI0/XI29/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM0 N_XI0/XI29/XI10/NET34_XI0/XI29/XI10/MM0_d
+ N_WL<54>_XI0/XI29/XI10/MM0_g N_BL<5>_XI0/XI29/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM1 N_XI0/XI29/XI10/NET33_XI0/XI29/XI10/MM1_d
+ N_XI0/XI29/XI10/NET34_XI0/XI29/XI10/MM1_g N_VSS_XI0/XI29/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM9 N_XI0/XI29/XI10/NET36_XI0/XI29/XI10/MM9_d
+ N_WL<55>_XI0/XI29/XI10/MM9_g N_BL<5>_XI0/XI29/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM6 N_XI0/XI29/XI10/NET35_XI0/XI29/XI10/MM6_d
+ N_XI0/XI29/XI10/NET36_XI0/XI29/XI10/MM6_g N_VSS_XI0/XI29/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM7 N_XI0/XI29/XI10/NET36_XI0/XI29/XI10/MM7_d
+ N_XI0/XI29/XI10/NET35_XI0/XI29/XI10/MM7_g N_VSS_XI0/XI29/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM8 N_XI0/XI29/XI10/NET35_XI0/XI29/XI10/MM8_d
+ N_WL<55>_XI0/XI29/XI10/MM8_g N_BLN<5>_XI0/XI29/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI10/MM5 N_XI0/XI29/XI10/NET34_XI0/XI29/XI10/MM5_d
+ N_XI0/XI29/XI10/NET33_XI0/XI29/XI10/MM5_g N_VDD_XI0/XI29/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI10/MM4 N_XI0/XI29/XI10/NET33_XI0/XI29/XI10/MM4_d
+ N_XI0/XI29/XI10/NET34_XI0/XI29/XI10/MM4_g N_VDD_XI0/XI29/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI10/MM10 N_XI0/XI29/XI10/NET35_XI0/XI29/XI10/MM10_d
+ N_XI0/XI29/XI10/NET36_XI0/XI29/XI10/MM10_g N_VDD_XI0/XI29/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI10/MM11 N_XI0/XI29/XI10/NET36_XI0/XI29/XI10/MM11_d
+ N_XI0/XI29/XI10/NET35_XI0/XI29/XI10/MM11_g N_VDD_XI0/XI29/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI11/MM2 N_XI0/XI29/XI11/NET34_XI0/XI29/XI11/MM2_d
+ N_XI0/XI29/XI11/NET33_XI0/XI29/XI11/MM2_g N_VSS_XI0/XI29/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM3 N_XI0/XI29/XI11/NET33_XI0/XI29/XI11/MM3_d
+ N_WL<54>_XI0/XI29/XI11/MM3_g N_BLN<4>_XI0/XI29/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM0 N_XI0/XI29/XI11/NET34_XI0/XI29/XI11/MM0_d
+ N_WL<54>_XI0/XI29/XI11/MM0_g N_BL<4>_XI0/XI29/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM1 N_XI0/XI29/XI11/NET33_XI0/XI29/XI11/MM1_d
+ N_XI0/XI29/XI11/NET34_XI0/XI29/XI11/MM1_g N_VSS_XI0/XI29/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM9 N_XI0/XI29/XI11/NET36_XI0/XI29/XI11/MM9_d
+ N_WL<55>_XI0/XI29/XI11/MM9_g N_BL<4>_XI0/XI29/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM6 N_XI0/XI29/XI11/NET35_XI0/XI29/XI11/MM6_d
+ N_XI0/XI29/XI11/NET36_XI0/XI29/XI11/MM6_g N_VSS_XI0/XI29/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM7 N_XI0/XI29/XI11/NET36_XI0/XI29/XI11/MM7_d
+ N_XI0/XI29/XI11/NET35_XI0/XI29/XI11/MM7_g N_VSS_XI0/XI29/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM8 N_XI0/XI29/XI11/NET35_XI0/XI29/XI11/MM8_d
+ N_WL<55>_XI0/XI29/XI11/MM8_g N_BLN<4>_XI0/XI29/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI11/MM5 N_XI0/XI29/XI11/NET34_XI0/XI29/XI11/MM5_d
+ N_XI0/XI29/XI11/NET33_XI0/XI29/XI11/MM5_g N_VDD_XI0/XI29/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI11/MM4 N_XI0/XI29/XI11/NET33_XI0/XI29/XI11/MM4_d
+ N_XI0/XI29/XI11/NET34_XI0/XI29/XI11/MM4_g N_VDD_XI0/XI29/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI11/MM10 N_XI0/XI29/XI11/NET35_XI0/XI29/XI11/MM10_d
+ N_XI0/XI29/XI11/NET36_XI0/XI29/XI11/MM10_g N_VDD_XI0/XI29/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI11/MM11 N_XI0/XI29/XI11/NET36_XI0/XI29/XI11/MM11_d
+ N_XI0/XI29/XI11/NET35_XI0/XI29/XI11/MM11_g N_VDD_XI0/XI29/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI12/MM2 N_XI0/XI29/XI12/NET34_XI0/XI29/XI12/MM2_d
+ N_XI0/XI29/XI12/NET33_XI0/XI29/XI12/MM2_g N_VSS_XI0/XI29/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM3 N_XI0/XI29/XI12/NET33_XI0/XI29/XI12/MM3_d
+ N_WL<54>_XI0/XI29/XI12/MM3_g N_BLN<3>_XI0/XI29/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM0 N_XI0/XI29/XI12/NET34_XI0/XI29/XI12/MM0_d
+ N_WL<54>_XI0/XI29/XI12/MM0_g N_BL<3>_XI0/XI29/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM1 N_XI0/XI29/XI12/NET33_XI0/XI29/XI12/MM1_d
+ N_XI0/XI29/XI12/NET34_XI0/XI29/XI12/MM1_g N_VSS_XI0/XI29/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM9 N_XI0/XI29/XI12/NET36_XI0/XI29/XI12/MM9_d
+ N_WL<55>_XI0/XI29/XI12/MM9_g N_BL<3>_XI0/XI29/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM6 N_XI0/XI29/XI12/NET35_XI0/XI29/XI12/MM6_d
+ N_XI0/XI29/XI12/NET36_XI0/XI29/XI12/MM6_g N_VSS_XI0/XI29/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM7 N_XI0/XI29/XI12/NET36_XI0/XI29/XI12/MM7_d
+ N_XI0/XI29/XI12/NET35_XI0/XI29/XI12/MM7_g N_VSS_XI0/XI29/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM8 N_XI0/XI29/XI12/NET35_XI0/XI29/XI12/MM8_d
+ N_WL<55>_XI0/XI29/XI12/MM8_g N_BLN<3>_XI0/XI29/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI12/MM5 N_XI0/XI29/XI12/NET34_XI0/XI29/XI12/MM5_d
+ N_XI0/XI29/XI12/NET33_XI0/XI29/XI12/MM5_g N_VDD_XI0/XI29/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI12/MM4 N_XI0/XI29/XI12/NET33_XI0/XI29/XI12/MM4_d
+ N_XI0/XI29/XI12/NET34_XI0/XI29/XI12/MM4_g N_VDD_XI0/XI29/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI12/MM10 N_XI0/XI29/XI12/NET35_XI0/XI29/XI12/MM10_d
+ N_XI0/XI29/XI12/NET36_XI0/XI29/XI12/MM10_g N_VDD_XI0/XI29/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI12/MM11 N_XI0/XI29/XI12/NET36_XI0/XI29/XI12/MM11_d
+ N_XI0/XI29/XI12/NET35_XI0/XI29/XI12/MM11_g N_VDD_XI0/XI29/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI13/MM2 N_XI0/XI29/XI13/NET34_XI0/XI29/XI13/MM2_d
+ N_XI0/XI29/XI13/NET33_XI0/XI29/XI13/MM2_g N_VSS_XI0/XI29/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM3 N_XI0/XI29/XI13/NET33_XI0/XI29/XI13/MM3_d
+ N_WL<54>_XI0/XI29/XI13/MM3_g N_BLN<2>_XI0/XI29/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM0 N_XI0/XI29/XI13/NET34_XI0/XI29/XI13/MM0_d
+ N_WL<54>_XI0/XI29/XI13/MM0_g N_BL<2>_XI0/XI29/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM1 N_XI0/XI29/XI13/NET33_XI0/XI29/XI13/MM1_d
+ N_XI0/XI29/XI13/NET34_XI0/XI29/XI13/MM1_g N_VSS_XI0/XI29/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM9 N_XI0/XI29/XI13/NET36_XI0/XI29/XI13/MM9_d
+ N_WL<55>_XI0/XI29/XI13/MM9_g N_BL<2>_XI0/XI29/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM6 N_XI0/XI29/XI13/NET35_XI0/XI29/XI13/MM6_d
+ N_XI0/XI29/XI13/NET36_XI0/XI29/XI13/MM6_g N_VSS_XI0/XI29/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM7 N_XI0/XI29/XI13/NET36_XI0/XI29/XI13/MM7_d
+ N_XI0/XI29/XI13/NET35_XI0/XI29/XI13/MM7_g N_VSS_XI0/XI29/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM8 N_XI0/XI29/XI13/NET35_XI0/XI29/XI13/MM8_d
+ N_WL<55>_XI0/XI29/XI13/MM8_g N_BLN<2>_XI0/XI29/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI13/MM5 N_XI0/XI29/XI13/NET34_XI0/XI29/XI13/MM5_d
+ N_XI0/XI29/XI13/NET33_XI0/XI29/XI13/MM5_g N_VDD_XI0/XI29/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI13/MM4 N_XI0/XI29/XI13/NET33_XI0/XI29/XI13/MM4_d
+ N_XI0/XI29/XI13/NET34_XI0/XI29/XI13/MM4_g N_VDD_XI0/XI29/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI13/MM10 N_XI0/XI29/XI13/NET35_XI0/XI29/XI13/MM10_d
+ N_XI0/XI29/XI13/NET36_XI0/XI29/XI13/MM10_g N_VDD_XI0/XI29/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI13/MM11 N_XI0/XI29/XI13/NET36_XI0/XI29/XI13/MM11_d
+ N_XI0/XI29/XI13/NET35_XI0/XI29/XI13/MM11_g N_VDD_XI0/XI29/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI14/MM2 N_XI0/XI29/XI14/NET34_XI0/XI29/XI14/MM2_d
+ N_XI0/XI29/XI14/NET33_XI0/XI29/XI14/MM2_g N_VSS_XI0/XI29/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM3 N_XI0/XI29/XI14/NET33_XI0/XI29/XI14/MM3_d
+ N_WL<54>_XI0/XI29/XI14/MM3_g N_BLN<1>_XI0/XI29/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM0 N_XI0/XI29/XI14/NET34_XI0/XI29/XI14/MM0_d
+ N_WL<54>_XI0/XI29/XI14/MM0_g N_BL<1>_XI0/XI29/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM1 N_XI0/XI29/XI14/NET33_XI0/XI29/XI14/MM1_d
+ N_XI0/XI29/XI14/NET34_XI0/XI29/XI14/MM1_g N_VSS_XI0/XI29/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM9 N_XI0/XI29/XI14/NET36_XI0/XI29/XI14/MM9_d
+ N_WL<55>_XI0/XI29/XI14/MM9_g N_BL<1>_XI0/XI29/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM6 N_XI0/XI29/XI14/NET35_XI0/XI29/XI14/MM6_d
+ N_XI0/XI29/XI14/NET36_XI0/XI29/XI14/MM6_g N_VSS_XI0/XI29/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM7 N_XI0/XI29/XI14/NET36_XI0/XI29/XI14/MM7_d
+ N_XI0/XI29/XI14/NET35_XI0/XI29/XI14/MM7_g N_VSS_XI0/XI29/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM8 N_XI0/XI29/XI14/NET35_XI0/XI29/XI14/MM8_d
+ N_WL<55>_XI0/XI29/XI14/MM8_g N_BLN<1>_XI0/XI29/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI14/MM5 N_XI0/XI29/XI14/NET34_XI0/XI29/XI14/MM5_d
+ N_XI0/XI29/XI14/NET33_XI0/XI29/XI14/MM5_g N_VDD_XI0/XI29/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI14/MM4 N_XI0/XI29/XI14/NET33_XI0/XI29/XI14/MM4_d
+ N_XI0/XI29/XI14/NET34_XI0/XI29/XI14/MM4_g N_VDD_XI0/XI29/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI14/MM10 N_XI0/XI29/XI14/NET35_XI0/XI29/XI14/MM10_d
+ N_XI0/XI29/XI14/NET36_XI0/XI29/XI14/MM10_g N_VDD_XI0/XI29/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI14/MM11 N_XI0/XI29/XI14/NET36_XI0/XI29/XI14/MM11_d
+ N_XI0/XI29/XI14/NET35_XI0/XI29/XI14/MM11_g N_VDD_XI0/XI29/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI15/MM2 N_XI0/XI29/XI15/NET34_XI0/XI29/XI15/MM2_d
+ N_XI0/XI29/XI15/NET33_XI0/XI29/XI15/MM2_g N_VSS_XI0/XI29/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM3 N_XI0/XI29/XI15/NET33_XI0/XI29/XI15/MM3_d
+ N_WL<54>_XI0/XI29/XI15/MM3_g N_BLN<0>_XI0/XI29/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM0 N_XI0/XI29/XI15/NET34_XI0/XI29/XI15/MM0_d
+ N_WL<54>_XI0/XI29/XI15/MM0_g N_BL<0>_XI0/XI29/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM1 N_XI0/XI29/XI15/NET33_XI0/XI29/XI15/MM1_d
+ N_XI0/XI29/XI15/NET34_XI0/XI29/XI15/MM1_g N_VSS_XI0/XI29/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM9 N_XI0/XI29/XI15/NET36_XI0/XI29/XI15/MM9_d
+ N_WL<55>_XI0/XI29/XI15/MM9_g N_BL<0>_XI0/XI29/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM6 N_XI0/XI29/XI15/NET35_XI0/XI29/XI15/MM6_d
+ N_XI0/XI29/XI15/NET36_XI0/XI29/XI15/MM6_g N_VSS_XI0/XI29/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM7 N_XI0/XI29/XI15/NET36_XI0/XI29/XI15/MM7_d
+ N_XI0/XI29/XI15/NET35_XI0/XI29/XI15/MM7_g N_VSS_XI0/XI29/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM8 N_XI0/XI29/XI15/NET35_XI0/XI29/XI15/MM8_d
+ N_WL<55>_XI0/XI29/XI15/MM8_g N_BLN<0>_XI0/XI29/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI29/XI15/MM5 N_XI0/XI29/XI15/NET34_XI0/XI29/XI15/MM5_d
+ N_XI0/XI29/XI15/NET33_XI0/XI29/XI15/MM5_g N_VDD_XI0/XI29/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI15/MM4 N_XI0/XI29/XI15/NET33_XI0/XI29/XI15/MM4_d
+ N_XI0/XI29/XI15/NET34_XI0/XI29/XI15/MM4_g N_VDD_XI0/XI29/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI15/MM10 N_XI0/XI29/XI15/NET35_XI0/XI29/XI15/MM10_d
+ N_XI0/XI29/XI15/NET36_XI0/XI29/XI15/MM10_g N_VDD_XI0/XI29/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI29/XI15/MM11 N_XI0/XI29/XI15/NET36_XI0/XI29/XI15/MM11_d
+ N_XI0/XI29/XI15/NET35_XI0/XI29/XI15/MM11_g N_VDD_XI0/XI29/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI0/MM2 N_XI0/XI30/XI0/NET34_XI0/XI30/XI0/MM2_d
+ N_XI0/XI30/XI0/NET33_XI0/XI30/XI0/MM2_g N_VSS_XI0/XI30/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM3 N_XI0/XI30/XI0/NET33_XI0/XI30/XI0/MM3_d
+ N_WL<56>_XI0/XI30/XI0/MM3_g N_BLN<15>_XI0/XI30/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM0 N_XI0/XI30/XI0/NET34_XI0/XI30/XI0/MM0_d
+ N_WL<56>_XI0/XI30/XI0/MM0_g N_BL<15>_XI0/XI30/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM1 N_XI0/XI30/XI0/NET33_XI0/XI30/XI0/MM1_d
+ N_XI0/XI30/XI0/NET34_XI0/XI30/XI0/MM1_g N_VSS_XI0/XI30/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM9 N_XI0/XI30/XI0/NET36_XI0/XI30/XI0/MM9_d
+ N_WL<57>_XI0/XI30/XI0/MM9_g N_BL<15>_XI0/XI30/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM6 N_XI0/XI30/XI0/NET35_XI0/XI30/XI0/MM6_d
+ N_XI0/XI30/XI0/NET36_XI0/XI30/XI0/MM6_g N_VSS_XI0/XI30/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM7 N_XI0/XI30/XI0/NET36_XI0/XI30/XI0/MM7_d
+ N_XI0/XI30/XI0/NET35_XI0/XI30/XI0/MM7_g N_VSS_XI0/XI30/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM8 N_XI0/XI30/XI0/NET35_XI0/XI30/XI0/MM8_d
+ N_WL<57>_XI0/XI30/XI0/MM8_g N_BLN<15>_XI0/XI30/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI0/MM5 N_XI0/XI30/XI0/NET34_XI0/XI30/XI0/MM5_d
+ N_XI0/XI30/XI0/NET33_XI0/XI30/XI0/MM5_g N_VDD_XI0/XI30/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI0/MM4 N_XI0/XI30/XI0/NET33_XI0/XI30/XI0/MM4_d
+ N_XI0/XI30/XI0/NET34_XI0/XI30/XI0/MM4_g N_VDD_XI0/XI30/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI0/MM10 N_XI0/XI30/XI0/NET35_XI0/XI30/XI0/MM10_d
+ N_XI0/XI30/XI0/NET36_XI0/XI30/XI0/MM10_g N_VDD_XI0/XI30/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI0/MM11 N_XI0/XI30/XI0/NET36_XI0/XI30/XI0/MM11_d
+ N_XI0/XI30/XI0/NET35_XI0/XI30/XI0/MM11_g N_VDD_XI0/XI30/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI1/MM2 N_XI0/XI30/XI1/NET34_XI0/XI30/XI1/MM2_d
+ N_XI0/XI30/XI1/NET33_XI0/XI30/XI1/MM2_g N_VSS_XI0/XI30/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM3 N_XI0/XI30/XI1/NET33_XI0/XI30/XI1/MM3_d
+ N_WL<56>_XI0/XI30/XI1/MM3_g N_BLN<14>_XI0/XI30/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM0 N_XI0/XI30/XI1/NET34_XI0/XI30/XI1/MM0_d
+ N_WL<56>_XI0/XI30/XI1/MM0_g N_BL<14>_XI0/XI30/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM1 N_XI0/XI30/XI1/NET33_XI0/XI30/XI1/MM1_d
+ N_XI0/XI30/XI1/NET34_XI0/XI30/XI1/MM1_g N_VSS_XI0/XI30/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM9 N_XI0/XI30/XI1/NET36_XI0/XI30/XI1/MM9_d
+ N_WL<57>_XI0/XI30/XI1/MM9_g N_BL<14>_XI0/XI30/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM6 N_XI0/XI30/XI1/NET35_XI0/XI30/XI1/MM6_d
+ N_XI0/XI30/XI1/NET36_XI0/XI30/XI1/MM6_g N_VSS_XI0/XI30/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM7 N_XI0/XI30/XI1/NET36_XI0/XI30/XI1/MM7_d
+ N_XI0/XI30/XI1/NET35_XI0/XI30/XI1/MM7_g N_VSS_XI0/XI30/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM8 N_XI0/XI30/XI1/NET35_XI0/XI30/XI1/MM8_d
+ N_WL<57>_XI0/XI30/XI1/MM8_g N_BLN<14>_XI0/XI30/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI1/MM5 N_XI0/XI30/XI1/NET34_XI0/XI30/XI1/MM5_d
+ N_XI0/XI30/XI1/NET33_XI0/XI30/XI1/MM5_g N_VDD_XI0/XI30/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI1/MM4 N_XI0/XI30/XI1/NET33_XI0/XI30/XI1/MM4_d
+ N_XI0/XI30/XI1/NET34_XI0/XI30/XI1/MM4_g N_VDD_XI0/XI30/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI1/MM10 N_XI0/XI30/XI1/NET35_XI0/XI30/XI1/MM10_d
+ N_XI0/XI30/XI1/NET36_XI0/XI30/XI1/MM10_g N_VDD_XI0/XI30/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI1/MM11 N_XI0/XI30/XI1/NET36_XI0/XI30/XI1/MM11_d
+ N_XI0/XI30/XI1/NET35_XI0/XI30/XI1/MM11_g N_VDD_XI0/XI30/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI2/MM2 N_XI0/XI30/XI2/NET34_XI0/XI30/XI2/MM2_d
+ N_XI0/XI30/XI2/NET33_XI0/XI30/XI2/MM2_g N_VSS_XI0/XI30/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM3 N_XI0/XI30/XI2/NET33_XI0/XI30/XI2/MM3_d
+ N_WL<56>_XI0/XI30/XI2/MM3_g N_BLN<13>_XI0/XI30/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM0 N_XI0/XI30/XI2/NET34_XI0/XI30/XI2/MM0_d
+ N_WL<56>_XI0/XI30/XI2/MM0_g N_BL<13>_XI0/XI30/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM1 N_XI0/XI30/XI2/NET33_XI0/XI30/XI2/MM1_d
+ N_XI0/XI30/XI2/NET34_XI0/XI30/XI2/MM1_g N_VSS_XI0/XI30/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM9 N_XI0/XI30/XI2/NET36_XI0/XI30/XI2/MM9_d
+ N_WL<57>_XI0/XI30/XI2/MM9_g N_BL<13>_XI0/XI30/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM6 N_XI0/XI30/XI2/NET35_XI0/XI30/XI2/MM6_d
+ N_XI0/XI30/XI2/NET36_XI0/XI30/XI2/MM6_g N_VSS_XI0/XI30/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM7 N_XI0/XI30/XI2/NET36_XI0/XI30/XI2/MM7_d
+ N_XI0/XI30/XI2/NET35_XI0/XI30/XI2/MM7_g N_VSS_XI0/XI30/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM8 N_XI0/XI30/XI2/NET35_XI0/XI30/XI2/MM8_d
+ N_WL<57>_XI0/XI30/XI2/MM8_g N_BLN<13>_XI0/XI30/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI2/MM5 N_XI0/XI30/XI2/NET34_XI0/XI30/XI2/MM5_d
+ N_XI0/XI30/XI2/NET33_XI0/XI30/XI2/MM5_g N_VDD_XI0/XI30/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI2/MM4 N_XI0/XI30/XI2/NET33_XI0/XI30/XI2/MM4_d
+ N_XI0/XI30/XI2/NET34_XI0/XI30/XI2/MM4_g N_VDD_XI0/XI30/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI2/MM10 N_XI0/XI30/XI2/NET35_XI0/XI30/XI2/MM10_d
+ N_XI0/XI30/XI2/NET36_XI0/XI30/XI2/MM10_g N_VDD_XI0/XI30/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI2/MM11 N_XI0/XI30/XI2/NET36_XI0/XI30/XI2/MM11_d
+ N_XI0/XI30/XI2/NET35_XI0/XI30/XI2/MM11_g N_VDD_XI0/XI30/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI3/MM2 N_XI0/XI30/XI3/NET34_XI0/XI30/XI3/MM2_d
+ N_XI0/XI30/XI3/NET33_XI0/XI30/XI3/MM2_g N_VSS_XI0/XI30/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM3 N_XI0/XI30/XI3/NET33_XI0/XI30/XI3/MM3_d
+ N_WL<56>_XI0/XI30/XI3/MM3_g N_BLN<12>_XI0/XI30/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM0 N_XI0/XI30/XI3/NET34_XI0/XI30/XI3/MM0_d
+ N_WL<56>_XI0/XI30/XI3/MM0_g N_BL<12>_XI0/XI30/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM1 N_XI0/XI30/XI3/NET33_XI0/XI30/XI3/MM1_d
+ N_XI0/XI30/XI3/NET34_XI0/XI30/XI3/MM1_g N_VSS_XI0/XI30/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM9 N_XI0/XI30/XI3/NET36_XI0/XI30/XI3/MM9_d
+ N_WL<57>_XI0/XI30/XI3/MM9_g N_BL<12>_XI0/XI30/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM6 N_XI0/XI30/XI3/NET35_XI0/XI30/XI3/MM6_d
+ N_XI0/XI30/XI3/NET36_XI0/XI30/XI3/MM6_g N_VSS_XI0/XI30/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM7 N_XI0/XI30/XI3/NET36_XI0/XI30/XI3/MM7_d
+ N_XI0/XI30/XI3/NET35_XI0/XI30/XI3/MM7_g N_VSS_XI0/XI30/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM8 N_XI0/XI30/XI3/NET35_XI0/XI30/XI3/MM8_d
+ N_WL<57>_XI0/XI30/XI3/MM8_g N_BLN<12>_XI0/XI30/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI3/MM5 N_XI0/XI30/XI3/NET34_XI0/XI30/XI3/MM5_d
+ N_XI0/XI30/XI3/NET33_XI0/XI30/XI3/MM5_g N_VDD_XI0/XI30/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI3/MM4 N_XI0/XI30/XI3/NET33_XI0/XI30/XI3/MM4_d
+ N_XI0/XI30/XI3/NET34_XI0/XI30/XI3/MM4_g N_VDD_XI0/XI30/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI3/MM10 N_XI0/XI30/XI3/NET35_XI0/XI30/XI3/MM10_d
+ N_XI0/XI30/XI3/NET36_XI0/XI30/XI3/MM10_g N_VDD_XI0/XI30/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI3/MM11 N_XI0/XI30/XI3/NET36_XI0/XI30/XI3/MM11_d
+ N_XI0/XI30/XI3/NET35_XI0/XI30/XI3/MM11_g N_VDD_XI0/XI30/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI4/MM2 N_XI0/XI30/XI4/NET34_XI0/XI30/XI4/MM2_d
+ N_XI0/XI30/XI4/NET33_XI0/XI30/XI4/MM2_g N_VSS_XI0/XI30/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM3 N_XI0/XI30/XI4/NET33_XI0/XI30/XI4/MM3_d
+ N_WL<56>_XI0/XI30/XI4/MM3_g N_BLN<11>_XI0/XI30/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM0 N_XI0/XI30/XI4/NET34_XI0/XI30/XI4/MM0_d
+ N_WL<56>_XI0/XI30/XI4/MM0_g N_BL<11>_XI0/XI30/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM1 N_XI0/XI30/XI4/NET33_XI0/XI30/XI4/MM1_d
+ N_XI0/XI30/XI4/NET34_XI0/XI30/XI4/MM1_g N_VSS_XI0/XI30/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM9 N_XI0/XI30/XI4/NET36_XI0/XI30/XI4/MM9_d
+ N_WL<57>_XI0/XI30/XI4/MM9_g N_BL<11>_XI0/XI30/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM6 N_XI0/XI30/XI4/NET35_XI0/XI30/XI4/MM6_d
+ N_XI0/XI30/XI4/NET36_XI0/XI30/XI4/MM6_g N_VSS_XI0/XI30/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM7 N_XI0/XI30/XI4/NET36_XI0/XI30/XI4/MM7_d
+ N_XI0/XI30/XI4/NET35_XI0/XI30/XI4/MM7_g N_VSS_XI0/XI30/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM8 N_XI0/XI30/XI4/NET35_XI0/XI30/XI4/MM8_d
+ N_WL<57>_XI0/XI30/XI4/MM8_g N_BLN<11>_XI0/XI30/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI4/MM5 N_XI0/XI30/XI4/NET34_XI0/XI30/XI4/MM5_d
+ N_XI0/XI30/XI4/NET33_XI0/XI30/XI4/MM5_g N_VDD_XI0/XI30/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI4/MM4 N_XI0/XI30/XI4/NET33_XI0/XI30/XI4/MM4_d
+ N_XI0/XI30/XI4/NET34_XI0/XI30/XI4/MM4_g N_VDD_XI0/XI30/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI4/MM10 N_XI0/XI30/XI4/NET35_XI0/XI30/XI4/MM10_d
+ N_XI0/XI30/XI4/NET36_XI0/XI30/XI4/MM10_g N_VDD_XI0/XI30/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI4/MM11 N_XI0/XI30/XI4/NET36_XI0/XI30/XI4/MM11_d
+ N_XI0/XI30/XI4/NET35_XI0/XI30/XI4/MM11_g N_VDD_XI0/XI30/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI5/MM2 N_XI0/XI30/XI5/NET34_XI0/XI30/XI5/MM2_d
+ N_XI0/XI30/XI5/NET33_XI0/XI30/XI5/MM2_g N_VSS_XI0/XI30/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM3 N_XI0/XI30/XI5/NET33_XI0/XI30/XI5/MM3_d
+ N_WL<56>_XI0/XI30/XI5/MM3_g N_BLN<10>_XI0/XI30/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM0 N_XI0/XI30/XI5/NET34_XI0/XI30/XI5/MM0_d
+ N_WL<56>_XI0/XI30/XI5/MM0_g N_BL<10>_XI0/XI30/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM1 N_XI0/XI30/XI5/NET33_XI0/XI30/XI5/MM1_d
+ N_XI0/XI30/XI5/NET34_XI0/XI30/XI5/MM1_g N_VSS_XI0/XI30/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM9 N_XI0/XI30/XI5/NET36_XI0/XI30/XI5/MM9_d
+ N_WL<57>_XI0/XI30/XI5/MM9_g N_BL<10>_XI0/XI30/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM6 N_XI0/XI30/XI5/NET35_XI0/XI30/XI5/MM6_d
+ N_XI0/XI30/XI5/NET36_XI0/XI30/XI5/MM6_g N_VSS_XI0/XI30/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM7 N_XI0/XI30/XI5/NET36_XI0/XI30/XI5/MM7_d
+ N_XI0/XI30/XI5/NET35_XI0/XI30/XI5/MM7_g N_VSS_XI0/XI30/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM8 N_XI0/XI30/XI5/NET35_XI0/XI30/XI5/MM8_d
+ N_WL<57>_XI0/XI30/XI5/MM8_g N_BLN<10>_XI0/XI30/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI5/MM5 N_XI0/XI30/XI5/NET34_XI0/XI30/XI5/MM5_d
+ N_XI0/XI30/XI5/NET33_XI0/XI30/XI5/MM5_g N_VDD_XI0/XI30/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI5/MM4 N_XI0/XI30/XI5/NET33_XI0/XI30/XI5/MM4_d
+ N_XI0/XI30/XI5/NET34_XI0/XI30/XI5/MM4_g N_VDD_XI0/XI30/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI5/MM10 N_XI0/XI30/XI5/NET35_XI0/XI30/XI5/MM10_d
+ N_XI0/XI30/XI5/NET36_XI0/XI30/XI5/MM10_g N_VDD_XI0/XI30/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI5/MM11 N_XI0/XI30/XI5/NET36_XI0/XI30/XI5/MM11_d
+ N_XI0/XI30/XI5/NET35_XI0/XI30/XI5/MM11_g N_VDD_XI0/XI30/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI6/MM2 N_XI0/XI30/XI6/NET34_XI0/XI30/XI6/MM2_d
+ N_XI0/XI30/XI6/NET33_XI0/XI30/XI6/MM2_g N_VSS_XI0/XI30/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM3 N_XI0/XI30/XI6/NET33_XI0/XI30/XI6/MM3_d
+ N_WL<56>_XI0/XI30/XI6/MM3_g N_BLN<9>_XI0/XI30/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM0 N_XI0/XI30/XI6/NET34_XI0/XI30/XI6/MM0_d
+ N_WL<56>_XI0/XI30/XI6/MM0_g N_BL<9>_XI0/XI30/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM1 N_XI0/XI30/XI6/NET33_XI0/XI30/XI6/MM1_d
+ N_XI0/XI30/XI6/NET34_XI0/XI30/XI6/MM1_g N_VSS_XI0/XI30/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM9 N_XI0/XI30/XI6/NET36_XI0/XI30/XI6/MM9_d
+ N_WL<57>_XI0/XI30/XI6/MM9_g N_BL<9>_XI0/XI30/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM6 N_XI0/XI30/XI6/NET35_XI0/XI30/XI6/MM6_d
+ N_XI0/XI30/XI6/NET36_XI0/XI30/XI6/MM6_g N_VSS_XI0/XI30/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM7 N_XI0/XI30/XI6/NET36_XI0/XI30/XI6/MM7_d
+ N_XI0/XI30/XI6/NET35_XI0/XI30/XI6/MM7_g N_VSS_XI0/XI30/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM8 N_XI0/XI30/XI6/NET35_XI0/XI30/XI6/MM8_d
+ N_WL<57>_XI0/XI30/XI6/MM8_g N_BLN<9>_XI0/XI30/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI6/MM5 N_XI0/XI30/XI6/NET34_XI0/XI30/XI6/MM5_d
+ N_XI0/XI30/XI6/NET33_XI0/XI30/XI6/MM5_g N_VDD_XI0/XI30/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI6/MM4 N_XI0/XI30/XI6/NET33_XI0/XI30/XI6/MM4_d
+ N_XI0/XI30/XI6/NET34_XI0/XI30/XI6/MM4_g N_VDD_XI0/XI30/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI6/MM10 N_XI0/XI30/XI6/NET35_XI0/XI30/XI6/MM10_d
+ N_XI0/XI30/XI6/NET36_XI0/XI30/XI6/MM10_g N_VDD_XI0/XI30/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI6/MM11 N_XI0/XI30/XI6/NET36_XI0/XI30/XI6/MM11_d
+ N_XI0/XI30/XI6/NET35_XI0/XI30/XI6/MM11_g N_VDD_XI0/XI30/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI7/MM2 N_XI0/XI30/XI7/NET34_XI0/XI30/XI7/MM2_d
+ N_XI0/XI30/XI7/NET33_XI0/XI30/XI7/MM2_g N_VSS_XI0/XI30/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM3 N_XI0/XI30/XI7/NET33_XI0/XI30/XI7/MM3_d
+ N_WL<56>_XI0/XI30/XI7/MM3_g N_BLN<8>_XI0/XI30/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM0 N_XI0/XI30/XI7/NET34_XI0/XI30/XI7/MM0_d
+ N_WL<56>_XI0/XI30/XI7/MM0_g N_BL<8>_XI0/XI30/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM1 N_XI0/XI30/XI7/NET33_XI0/XI30/XI7/MM1_d
+ N_XI0/XI30/XI7/NET34_XI0/XI30/XI7/MM1_g N_VSS_XI0/XI30/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM9 N_XI0/XI30/XI7/NET36_XI0/XI30/XI7/MM9_d
+ N_WL<57>_XI0/XI30/XI7/MM9_g N_BL<8>_XI0/XI30/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM6 N_XI0/XI30/XI7/NET35_XI0/XI30/XI7/MM6_d
+ N_XI0/XI30/XI7/NET36_XI0/XI30/XI7/MM6_g N_VSS_XI0/XI30/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM7 N_XI0/XI30/XI7/NET36_XI0/XI30/XI7/MM7_d
+ N_XI0/XI30/XI7/NET35_XI0/XI30/XI7/MM7_g N_VSS_XI0/XI30/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM8 N_XI0/XI30/XI7/NET35_XI0/XI30/XI7/MM8_d
+ N_WL<57>_XI0/XI30/XI7/MM8_g N_BLN<8>_XI0/XI30/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI7/MM5 N_XI0/XI30/XI7/NET34_XI0/XI30/XI7/MM5_d
+ N_XI0/XI30/XI7/NET33_XI0/XI30/XI7/MM5_g N_VDD_XI0/XI30/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI7/MM4 N_XI0/XI30/XI7/NET33_XI0/XI30/XI7/MM4_d
+ N_XI0/XI30/XI7/NET34_XI0/XI30/XI7/MM4_g N_VDD_XI0/XI30/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI7/MM10 N_XI0/XI30/XI7/NET35_XI0/XI30/XI7/MM10_d
+ N_XI0/XI30/XI7/NET36_XI0/XI30/XI7/MM10_g N_VDD_XI0/XI30/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI7/MM11 N_XI0/XI30/XI7/NET36_XI0/XI30/XI7/MM11_d
+ N_XI0/XI30/XI7/NET35_XI0/XI30/XI7/MM11_g N_VDD_XI0/XI30/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI8/MM2 N_XI0/XI30/XI8/NET34_XI0/XI30/XI8/MM2_d
+ N_XI0/XI30/XI8/NET33_XI0/XI30/XI8/MM2_g N_VSS_XI0/XI30/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM3 N_XI0/XI30/XI8/NET33_XI0/XI30/XI8/MM3_d
+ N_WL<56>_XI0/XI30/XI8/MM3_g N_BLN<7>_XI0/XI30/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM0 N_XI0/XI30/XI8/NET34_XI0/XI30/XI8/MM0_d
+ N_WL<56>_XI0/XI30/XI8/MM0_g N_BL<7>_XI0/XI30/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM1 N_XI0/XI30/XI8/NET33_XI0/XI30/XI8/MM1_d
+ N_XI0/XI30/XI8/NET34_XI0/XI30/XI8/MM1_g N_VSS_XI0/XI30/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM9 N_XI0/XI30/XI8/NET36_XI0/XI30/XI8/MM9_d
+ N_WL<57>_XI0/XI30/XI8/MM9_g N_BL<7>_XI0/XI30/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM6 N_XI0/XI30/XI8/NET35_XI0/XI30/XI8/MM6_d
+ N_XI0/XI30/XI8/NET36_XI0/XI30/XI8/MM6_g N_VSS_XI0/XI30/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM7 N_XI0/XI30/XI8/NET36_XI0/XI30/XI8/MM7_d
+ N_XI0/XI30/XI8/NET35_XI0/XI30/XI8/MM7_g N_VSS_XI0/XI30/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM8 N_XI0/XI30/XI8/NET35_XI0/XI30/XI8/MM8_d
+ N_WL<57>_XI0/XI30/XI8/MM8_g N_BLN<7>_XI0/XI30/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI8/MM5 N_XI0/XI30/XI8/NET34_XI0/XI30/XI8/MM5_d
+ N_XI0/XI30/XI8/NET33_XI0/XI30/XI8/MM5_g N_VDD_XI0/XI30/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI8/MM4 N_XI0/XI30/XI8/NET33_XI0/XI30/XI8/MM4_d
+ N_XI0/XI30/XI8/NET34_XI0/XI30/XI8/MM4_g N_VDD_XI0/XI30/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI8/MM10 N_XI0/XI30/XI8/NET35_XI0/XI30/XI8/MM10_d
+ N_XI0/XI30/XI8/NET36_XI0/XI30/XI8/MM10_g N_VDD_XI0/XI30/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI8/MM11 N_XI0/XI30/XI8/NET36_XI0/XI30/XI8/MM11_d
+ N_XI0/XI30/XI8/NET35_XI0/XI30/XI8/MM11_g N_VDD_XI0/XI30/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI9/MM2 N_XI0/XI30/XI9/NET34_XI0/XI30/XI9/MM2_d
+ N_XI0/XI30/XI9/NET33_XI0/XI30/XI9/MM2_g N_VSS_XI0/XI30/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM3 N_XI0/XI30/XI9/NET33_XI0/XI30/XI9/MM3_d
+ N_WL<56>_XI0/XI30/XI9/MM3_g N_BLN<6>_XI0/XI30/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM0 N_XI0/XI30/XI9/NET34_XI0/XI30/XI9/MM0_d
+ N_WL<56>_XI0/XI30/XI9/MM0_g N_BL<6>_XI0/XI30/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM1 N_XI0/XI30/XI9/NET33_XI0/XI30/XI9/MM1_d
+ N_XI0/XI30/XI9/NET34_XI0/XI30/XI9/MM1_g N_VSS_XI0/XI30/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM9 N_XI0/XI30/XI9/NET36_XI0/XI30/XI9/MM9_d
+ N_WL<57>_XI0/XI30/XI9/MM9_g N_BL<6>_XI0/XI30/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM6 N_XI0/XI30/XI9/NET35_XI0/XI30/XI9/MM6_d
+ N_XI0/XI30/XI9/NET36_XI0/XI30/XI9/MM6_g N_VSS_XI0/XI30/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM7 N_XI0/XI30/XI9/NET36_XI0/XI30/XI9/MM7_d
+ N_XI0/XI30/XI9/NET35_XI0/XI30/XI9/MM7_g N_VSS_XI0/XI30/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM8 N_XI0/XI30/XI9/NET35_XI0/XI30/XI9/MM8_d
+ N_WL<57>_XI0/XI30/XI9/MM8_g N_BLN<6>_XI0/XI30/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI9/MM5 N_XI0/XI30/XI9/NET34_XI0/XI30/XI9/MM5_d
+ N_XI0/XI30/XI9/NET33_XI0/XI30/XI9/MM5_g N_VDD_XI0/XI30/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI9/MM4 N_XI0/XI30/XI9/NET33_XI0/XI30/XI9/MM4_d
+ N_XI0/XI30/XI9/NET34_XI0/XI30/XI9/MM4_g N_VDD_XI0/XI30/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI9/MM10 N_XI0/XI30/XI9/NET35_XI0/XI30/XI9/MM10_d
+ N_XI0/XI30/XI9/NET36_XI0/XI30/XI9/MM10_g N_VDD_XI0/XI30/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI9/MM11 N_XI0/XI30/XI9/NET36_XI0/XI30/XI9/MM11_d
+ N_XI0/XI30/XI9/NET35_XI0/XI30/XI9/MM11_g N_VDD_XI0/XI30/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI10/MM2 N_XI0/XI30/XI10/NET34_XI0/XI30/XI10/MM2_d
+ N_XI0/XI30/XI10/NET33_XI0/XI30/XI10/MM2_g N_VSS_XI0/XI30/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM3 N_XI0/XI30/XI10/NET33_XI0/XI30/XI10/MM3_d
+ N_WL<56>_XI0/XI30/XI10/MM3_g N_BLN<5>_XI0/XI30/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM0 N_XI0/XI30/XI10/NET34_XI0/XI30/XI10/MM0_d
+ N_WL<56>_XI0/XI30/XI10/MM0_g N_BL<5>_XI0/XI30/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM1 N_XI0/XI30/XI10/NET33_XI0/XI30/XI10/MM1_d
+ N_XI0/XI30/XI10/NET34_XI0/XI30/XI10/MM1_g N_VSS_XI0/XI30/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM9 N_XI0/XI30/XI10/NET36_XI0/XI30/XI10/MM9_d
+ N_WL<57>_XI0/XI30/XI10/MM9_g N_BL<5>_XI0/XI30/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM6 N_XI0/XI30/XI10/NET35_XI0/XI30/XI10/MM6_d
+ N_XI0/XI30/XI10/NET36_XI0/XI30/XI10/MM6_g N_VSS_XI0/XI30/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM7 N_XI0/XI30/XI10/NET36_XI0/XI30/XI10/MM7_d
+ N_XI0/XI30/XI10/NET35_XI0/XI30/XI10/MM7_g N_VSS_XI0/XI30/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM8 N_XI0/XI30/XI10/NET35_XI0/XI30/XI10/MM8_d
+ N_WL<57>_XI0/XI30/XI10/MM8_g N_BLN<5>_XI0/XI30/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI10/MM5 N_XI0/XI30/XI10/NET34_XI0/XI30/XI10/MM5_d
+ N_XI0/XI30/XI10/NET33_XI0/XI30/XI10/MM5_g N_VDD_XI0/XI30/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI10/MM4 N_XI0/XI30/XI10/NET33_XI0/XI30/XI10/MM4_d
+ N_XI0/XI30/XI10/NET34_XI0/XI30/XI10/MM4_g N_VDD_XI0/XI30/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI10/MM10 N_XI0/XI30/XI10/NET35_XI0/XI30/XI10/MM10_d
+ N_XI0/XI30/XI10/NET36_XI0/XI30/XI10/MM10_g N_VDD_XI0/XI30/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI10/MM11 N_XI0/XI30/XI10/NET36_XI0/XI30/XI10/MM11_d
+ N_XI0/XI30/XI10/NET35_XI0/XI30/XI10/MM11_g N_VDD_XI0/XI30/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI11/MM2 N_XI0/XI30/XI11/NET34_XI0/XI30/XI11/MM2_d
+ N_XI0/XI30/XI11/NET33_XI0/XI30/XI11/MM2_g N_VSS_XI0/XI30/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM3 N_XI0/XI30/XI11/NET33_XI0/XI30/XI11/MM3_d
+ N_WL<56>_XI0/XI30/XI11/MM3_g N_BLN<4>_XI0/XI30/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM0 N_XI0/XI30/XI11/NET34_XI0/XI30/XI11/MM0_d
+ N_WL<56>_XI0/XI30/XI11/MM0_g N_BL<4>_XI0/XI30/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM1 N_XI0/XI30/XI11/NET33_XI0/XI30/XI11/MM1_d
+ N_XI0/XI30/XI11/NET34_XI0/XI30/XI11/MM1_g N_VSS_XI0/XI30/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM9 N_XI0/XI30/XI11/NET36_XI0/XI30/XI11/MM9_d
+ N_WL<57>_XI0/XI30/XI11/MM9_g N_BL<4>_XI0/XI30/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM6 N_XI0/XI30/XI11/NET35_XI0/XI30/XI11/MM6_d
+ N_XI0/XI30/XI11/NET36_XI0/XI30/XI11/MM6_g N_VSS_XI0/XI30/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM7 N_XI0/XI30/XI11/NET36_XI0/XI30/XI11/MM7_d
+ N_XI0/XI30/XI11/NET35_XI0/XI30/XI11/MM7_g N_VSS_XI0/XI30/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM8 N_XI0/XI30/XI11/NET35_XI0/XI30/XI11/MM8_d
+ N_WL<57>_XI0/XI30/XI11/MM8_g N_BLN<4>_XI0/XI30/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI11/MM5 N_XI0/XI30/XI11/NET34_XI0/XI30/XI11/MM5_d
+ N_XI0/XI30/XI11/NET33_XI0/XI30/XI11/MM5_g N_VDD_XI0/XI30/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI11/MM4 N_XI0/XI30/XI11/NET33_XI0/XI30/XI11/MM4_d
+ N_XI0/XI30/XI11/NET34_XI0/XI30/XI11/MM4_g N_VDD_XI0/XI30/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI11/MM10 N_XI0/XI30/XI11/NET35_XI0/XI30/XI11/MM10_d
+ N_XI0/XI30/XI11/NET36_XI0/XI30/XI11/MM10_g N_VDD_XI0/XI30/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI11/MM11 N_XI0/XI30/XI11/NET36_XI0/XI30/XI11/MM11_d
+ N_XI0/XI30/XI11/NET35_XI0/XI30/XI11/MM11_g N_VDD_XI0/XI30/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI12/MM2 N_XI0/XI30/XI12/NET34_XI0/XI30/XI12/MM2_d
+ N_XI0/XI30/XI12/NET33_XI0/XI30/XI12/MM2_g N_VSS_XI0/XI30/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM3 N_XI0/XI30/XI12/NET33_XI0/XI30/XI12/MM3_d
+ N_WL<56>_XI0/XI30/XI12/MM3_g N_BLN<3>_XI0/XI30/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM0 N_XI0/XI30/XI12/NET34_XI0/XI30/XI12/MM0_d
+ N_WL<56>_XI0/XI30/XI12/MM0_g N_BL<3>_XI0/XI30/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM1 N_XI0/XI30/XI12/NET33_XI0/XI30/XI12/MM1_d
+ N_XI0/XI30/XI12/NET34_XI0/XI30/XI12/MM1_g N_VSS_XI0/XI30/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM9 N_XI0/XI30/XI12/NET36_XI0/XI30/XI12/MM9_d
+ N_WL<57>_XI0/XI30/XI12/MM9_g N_BL<3>_XI0/XI30/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM6 N_XI0/XI30/XI12/NET35_XI0/XI30/XI12/MM6_d
+ N_XI0/XI30/XI12/NET36_XI0/XI30/XI12/MM6_g N_VSS_XI0/XI30/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM7 N_XI0/XI30/XI12/NET36_XI0/XI30/XI12/MM7_d
+ N_XI0/XI30/XI12/NET35_XI0/XI30/XI12/MM7_g N_VSS_XI0/XI30/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM8 N_XI0/XI30/XI12/NET35_XI0/XI30/XI12/MM8_d
+ N_WL<57>_XI0/XI30/XI12/MM8_g N_BLN<3>_XI0/XI30/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI12/MM5 N_XI0/XI30/XI12/NET34_XI0/XI30/XI12/MM5_d
+ N_XI0/XI30/XI12/NET33_XI0/XI30/XI12/MM5_g N_VDD_XI0/XI30/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI12/MM4 N_XI0/XI30/XI12/NET33_XI0/XI30/XI12/MM4_d
+ N_XI0/XI30/XI12/NET34_XI0/XI30/XI12/MM4_g N_VDD_XI0/XI30/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI12/MM10 N_XI0/XI30/XI12/NET35_XI0/XI30/XI12/MM10_d
+ N_XI0/XI30/XI12/NET36_XI0/XI30/XI12/MM10_g N_VDD_XI0/XI30/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI12/MM11 N_XI0/XI30/XI12/NET36_XI0/XI30/XI12/MM11_d
+ N_XI0/XI30/XI12/NET35_XI0/XI30/XI12/MM11_g N_VDD_XI0/XI30/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI13/MM2 N_XI0/XI30/XI13/NET34_XI0/XI30/XI13/MM2_d
+ N_XI0/XI30/XI13/NET33_XI0/XI30/XI13/MM2_g N_VSS_XI0/XI30/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM3 N_XI0/XI30/XI13/NET33_XI0/XI30/XI13/MM3_d
+ N_WL<56>_XI0/XI30/XI13/MM3_g N_BLN<2>_XI0/XI30/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM0 N_XI0/XI30/XI13/NET34_XI0/XI30/XI13/MM0_d
+ N_WL<56>_XI0/XI30/XI13/MM0_g N_BL<2>_XI0/XI30/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM1 N_XI0/XI30/XI13/NET33_XI0/XI30/XI13/MM1_d
+ N_XI0/XI30/XI13/NET34_XI0/XI30/XI13/MM1_g N_VSS_XI0/XI30/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM9 N_XI0/XI30/XI13/NET36_XI0/XI30/XI13/MM9_d
+ N_WL<57>_XI0/XI30/XI13/MM9_g N_BL<2>_XI0/XI30/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM6 N_XI0/XI30/XI13/NET35_XI0/XI30/XI13/MM6_d
+ N_XI0/XI30/XI13/NET36_XI0/XI30/XI13/MM6_g N_VSS_XI0/XI30/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM7 N_XI0/XI30/XI13/NET36_XI0/XI30/XI13/MM7_d
+ N_XI0/XI30/XI13/NET35_XI0/XI30/XI13/MM7_g N_VSS_XI0/XI30/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM8 N_XI0/XI30/XI13/NET35_XI0/XI30/XI13/MM8_d
+ N_WL<57>_XI0/XI30/XI13/MM8_g N_BLN<2>_XI0/XI30/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI13/MM5 N_XI0/XI30/XI13/NET34_XI0/XI30/XI13/MM5_d
+ N_XI0/XI30/XI13/NET33_XI0/XI30/XI13/MM5_g N_VDD_XI0/XI30/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI13/MM4 N_XI0/XI30/XI13/NET33_XI0/XI30/XI13/MM4_d
+ N_XI0/XI30/XI13/NET34_XI0/XI30/XI13/MM4_g N_VDD_XI0/XI30/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI13/MM10 N_XI0/XI30/XI13/NET35_XI0/XI30/XI13/MM10_d
+ N_XI0/XI30/XI13/NET36_XI0/XI30/XI13/MM10_g N_VDD_XI0/XI30/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI13/MM11 N_XI0/XI30/XI13/NET36_XI0/XI30/XI13/MM11_d
+ N_XI0/XI30/XI13/NET35_XI0/XI30/XI13/MM11_g N_VDD_XI0/XI30/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI14/MM2 N_XI0/XI30/XI14/NET34_XI0/XI30/XI14/MM2_d
+ N_XI0/XI30/XI14/NET33_XI0/XI30/XI14/MM2_g N_VSS_XI0/XI30/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM3 N_XI0/XI30/XI14/NET33_XI0/XI30/XI14/MM3_d
+ N_WL<56>_XI0/XI30/XI14/MM3_g N_BLN<1>_XI0/XI30/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM0 N_XI0/XI30/XI14/NET34_XI0/XI30/XI14/MM0_d
+ N_WL<56>_XI0/XI30/XI14/MM0_g N_BL<1>_XI0/XI30/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM1 N_XI0/XI30/XI14/NET33_XI0/XI30/XI14/MM1_d
+ N_XI0/XI30/XI14/NET34_XI0/XI30/XI14/MM1_g N_VSS_XI0/XI30/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM9 N_XI0/XI30/XI14/NET36_XI0/XI30/XI14/MM9_d
+ N_WL<57>_XI0/XI30/XI14/MM9_g N_BL<1>_XI0/XI30/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM6 N_XI0/XI30/XI14/NET35_XI0/XI30/XI14/MM6_d
+ N_XI0/XI30/XI14/NET36_XI0/XI30/XI14/MM6_g N_VSS_XI0/XI30/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM7 N_XI0/XI30/XI14/NET36_XI0/XI30/XI14/MM7_d
+ N_XI0/XI30/XI14/NET35_XI0/XI30/XI14/MM7_g N_VSS_XI0/XI30/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM8 N_XI0/XI30/XI14/NET35_XI0/XI30/XI14/MM8_d
+ N_WL<57>_XI0/XI30/XI14/MM8_g N_BLN<1>_XI0/XI30/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI14/MM5 N_XI0/XI30/XI14/NET34_XI0/XI30/XI14/MM5_d
+ N_XI0/XI30/XI14/NET33_XI0/XI30/XI14/MM5_g N_VDD_XI0/XI30/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI14/MM4 N_XI0/XI30/XI14/NET33_XI0/XI30/XI14/MM4_d
+ N_XI0/XI30/XI14/NET34_XI0/XI30/XI14/MM4_g N_VDD_XI0/XI30/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI14/MM10 N_XI0/XI30/XI14/NET35_XI0/XI30/XI14/MM10_d
+ N_XI0/XI30/XI14/NET36_XI0/XI30/XI14/MM10_g N_VDD_XI0/XI30/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI14/MM11 N_XI0/XI30/XI14/NET36_XI0/XI30/XI14/MM11_d
+ N_XI0/XI30/XI14/NET35_XI0/XI30/XI14/MM11_g N_VDD_XI0/XI30/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI15/MM2 N_XI0/XI30/XI15/NET34_XI0/XI30/XI15/MM2_d
+ N_XI0/XI30/XI15/NET33_XI0/XI30/XI15/MM2_g N_VSS_XI0/XI30/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM3 N_XI0/XI30/XI15/NET33_XI0/XI30/XI15/MM3_d
+ N_WL<56>_XI0/XI30/XI15/MM3_g N_BLN<0>_XI0/XI30/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM0 N_XI0/XI30/XI15/NET34_XI0/XI30/XI15/MM0_d
+ N_WL<56>_XI0/XI30/XI15/MM0_g N_BL<0>_XI0/XI30/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM1 N_XI0/XI30/XI15/NET33_XI0/XI30/XI15/MM1_d
+ N_XI0/XI30/XI15/NET34_XI0/XI30/XI15/MM1_g N_VSS_XI0/XI30/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM9 N_XI0/XI30/XI15/NET36_XI0/XI30/XI15/MM9_d
+ N_WL<57>_XI0/XI30/XI15/MM9_g N_BL<0>_XI0/XI30/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM6 N_XI0/XI30/XI15/NET35_XI0/XI30/XI15/MM6_d
+ N_XI0/XI30/XI15/NET36_XI0/XI30/XI15/MM6_g N_VSS_XI0/XI30/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM7 N_XI0/XI30/XI15/NET36_XI0/XI30/XI15/MM7_d
+ N_XI0/XI30/XI15/NET35_XI0/XI30/XI15/MM7_g N_VSS_XI0/XI30/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM8 N_XI0/XI30/XI15/NET35_XI0/XI30/XI15/MM8_d
+ N_WL<57>_XI0/XI30/XI15/MM8_g N_BLN<0>_XI0/XI30/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI30/XI15/MM5 N_XI0/XI30/XI15/NET34_XI0/XI30/XI15/MM5_d
+ N_XI0/XI30/XI15/NET33_XI0/XI30/XI15/MM5_g N_VDD_XI0/XI30/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI15/MM4 N_XI0/XI30/XI15/NET33_XI0/XI30/XI15/MM4_d
+ N_XI0/XI30/XI15/NET34_XI0/XI30/XI15/MM4_g N_VDD_XI0/XI30/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI15/MM10 N_XI0/XI30/XI15/NET35_XI0/XI30/XI15/MM10_d
+ N_XI0/XI30/XI15/NET36_XI0/XI30/XI15/MM10_g N_VDD_XI0/XI30/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI30/XI15/MM11 N_XI0/XI30/XI15/NET36_XI0/XI30/XI15/MM11_d
+ N_XI0/XI30/XI15/NET35_XI0/XI30/XI15/MM11_g N_VDD_XI0/XI30/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI0/MM2 N_XI0/XI31/XI0/NET34_XI0/XI31/XI0/MM2_d
+ N_XI0/XI31/XI0/NET33_XI0/XI31/XI0/MM2_g N_VSS_XI0/XI31/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM3 N_XI0/XI31/XI0/NET33_XI0/XI31/XI0/MM3_d
+ N_WL<58>_XI0/XI31/XI0/MM3_g N_BLN<15>_XI0/XI31/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM0 N_XI0/XI31/XI0/NET34_XI0/XI31/XI0/MM0_d
+ N_WL<58>_XI0/XI31/XI0/MM0_g N_BL<15>_XI0/XI31/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM1 N_XI0/XI31/XI0/NET33_XI0/XI31/XI0/MM1_d
+ N_XI0/XI31/XI0/NET34_XI0/XI31/XI0/MM1_g N_VSS_XI0/XI31/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM9 N_XI0/XI31/XI0/NET36_XI0/XI31/XI0/MM9_d
+ N_WL<59>_XI0/XI31/XI0/MM9_g N_BL<15>_XI0/XI31/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM6 N_XI0/XI31/XI0/NET35_XI0/XI31/XI0/MM6_d
+ N_XI0/XI31/XI0/NET36_XI0/XI31/XI0/MM6_g N_VSS_XI0/XI31/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM7 N_XI0/XI31/XI0/NET36_XI0/XI31/XI0/MM7_d
+ N_XI0/XI31/XI0/NET35_XI0/XI31/XI0/MM7_g N_VSS_XI0/XI31/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM8 N_XI0/XI31/XI0/NET35_XI0/XI31/XI0/MM8_d
+ N_WL<59>_XI0/XI31/XI0/MM8_g N_BLN<15>_XI0/XI31/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI0/MM5 N_XI0/XI31/XI0/NET34_XI0/XI31/XI0/MM5_d
+ N_XI0/XI31/XI0/NET33_XI0/XI31/XI0/MM5_g N_VDD_XI0/XI31/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI0/MM4 N_XI0/XI31/XI0/NET33_XI0/XI31/XI0/MM4_d
+ N_XI0/XI31/XI0/NET34_XI0/XI31/XI0/MM4_g N_VDD_XI0/XI31/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI0/MM10 N_XI0/XI31/XI0/NET35_XI0/XI31/XI0/MM10_d
+ N_XI0/XI31/XI0/NET36_XI0/XI31/XI0/MM10_g N_VDD_XI0/XI31/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI0/MM11 N_XI0/XI31/XI0/NET36_XI0/XI31/XI0/MM11_d
+ N_XI0/XI31/XI0/NET35_XI0/XI31/XI0/MM11_g N_VDD_XI0/XI31/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI1/MM2 N_XI0/XI31/XI1/NET34_XI0/XI31/XI1/MM2_d
+ N_XI0/XI31/XI1/NET33_XI0/XI31/XI1/MM2_g N_VSS_XI0/XI31/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM3 N_XI0/XI31/XI1/NET33_XI0/XI31/XI1/MM3_d
+ N_WL<58>_XI0/XI31/XI1/MM3_g N_BLN<14>_XI0/XI31/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM0 N_XI0/XI31/XI1/NET34_XI0/XI31/XI1/MM0_d
+ N_WL<58>_XI0/XI31/XI1/MM0_g N_BL<14>_XI0/XI31/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM1 N_XI0/XI31/XI1/NET33_XI0/XI31/XI1/MM1_d
+ N_XI0/XI31/XI1/NET34_XI0/XI31/XI1/MM1_g N_VSS_XI0/XI31/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM9 N_XI0/XI31/XI1/NET36_XI0/XI31/XI1/MM9_d
+ N_WL<59>_XI0/XI31/XI1/MM9_g N_BL<14>_XI0/XI31/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM6 N_XI0/XI31/XI1/NET35_XI0/XI31/XI1/MM6_d
+ N_XI0/XI31/XI1/NET36_XI0/XI31/XI1/MM6_g N_VSS_XI0/XI31/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM7 N_XI0/XI31/XI1/NET36_XI0/XI31/XI1/MM7_d
+ N_XI0/XI31/XI1/NET35_XI0/XI31/XI1/MM7_g N_VSS_XI0/XI31/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM8 N_XI0/XI31/XI1/NET35_XI0/XI31/XI1/MM8_d
+ N_WL<59>_XI0/XI31/XI1/MM8_g N_BLN<14>_XI0/XI31/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI1/MM5 N_XI0/XI31/XI1/NET34_XI0/XI31/XI1/MM5_d
+ N_XI0/XI31/XI1/NET33_XI0/XI31/XI1/MM5_g N_VDD_XI0/XI31/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI1/MM4 N_XI0/XI31/XI1/NET33_XI0/XI31/XI1/MM4_d
+ N_XI0/XI31/XI1/NET34_XI0/XI31/XI1/MM4_g N_VDD_XI0/XI31/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI1/MM10 N_XI0/XI31/XI1/NET35_XI0/XI31/XI1/MM10_d
+ N_XI0/XI31/XI1/NET36_XI0/XI31/XI1/MM10_g N_VDD_XI0/XI31/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI1/MM11 N_XI0/XI31/XI1/NET36_XI0/XI31/XI1/MM11_d
+ N_XI0/XI31/XI1/NET35_XI0/XI31/XI1/MM11_g N_VDD_XI0/XI31/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI2/MM2 N_XI0/XI31/XI2/NET34_XI0/XI31/XI2/MM2_d
+ N_XI0/XI31/XI2/NET33_XI0/XI31/XI2/MM2_g N_VSS_XI0/XI31/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM3 N_XI0/XI31/XI2/NET33_XI0/XI31/XI2/MM3_d
+ N_WL<58>_XI0/XI31/XI2/MM3_g N_BLN<13>_XI0/XI31/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM0 N_XI0/XI31/XI2/NET34_XI0/XI31/XI2/MM0_d
+ N_WL<58>_XI0/XI31/XI2/MM0_g N_BL<13>_XI0/XI31/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM1 N_XI0/XI31/XI2/NET33_XI0/XI31/XI2/MM1_d
+ N_XI0/XI31/XI2/NET34_XI0/XI31/XI2/MM1_g N_VSS_XI0/XI31/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM9 N_XI0/XI31/XI2/NET36_XI0/XI31/XI2/MM9_d
+ N_WL<59>_XI0/XI31/XI2/MM9_g N_BL<13>_XI0/XI31/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM6 N_XI0/XI31/XI2/NET35_XI0/XI31/XI2/MM6_d
+ N_XI0/XI31/XI2/NET36_XI0/XI31/XI2/MM6_g N_VSS_XI0/XI31/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM7 N_XI0/XI31/XI2/NET36_XI0/XI31/XI2/MM7_d
+ N_XI0/XI31/XI2/NET35_XI0/XI31/XI2/MM7_g N_VSS_XI0/XI31/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM8 N_XI0/XI31/XI2/NET35_XI0/XI31/XI2/MM8_d
+ N_WL<59>_XI0/XI31/XI2/MM8_g N_BLN<13>_XI0/XI31/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI2/MM5 N_XI0/XI31/XI2/NET34_XI0/XI31/XI2/MM5_d
+ N_XI0/XI31/XI2/NET33_XI0/XI31/XI2/MM5_g N_VDD_XI0/XI31/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI2/MM4 N_XI0/XI31/XI2/NET33_XI0/XI31/XI2/MM4_d
+ N_XI0/XI31/XI2/NET34_XI0/XI31/XI2/MM4_g N_VDD_XI0/XI31/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI2/MM10 N_XI0/XI31/XI2/NET35_XI0/XI31/XI2/MM10_d
+ N_XI0/XI31/XI2/NET36_XI0/XI31/XI2/MM10_g N_VDD_XI0/XI31/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI2/MM11 N_XI0/XI31/XI2/NET36_XI0/XI31/XI2/MM11_d
+ N_XI0/XI31/XI2/NET35_XI0/XI31/XI2/MM11_g N_VDD_XI0/XI31/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI3/MM2 N_XI0/XI31/XI3/NET34_XI0/XI31/XI3/MM2_d
+ N_XI0/XI31/XI3/NET33_XI0/XI31/XI3/MM2_g N_VSS_XI0/XI31/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM3 N_XI0/XI31/XI3/NET33_XI0/XI31/XI3/MM3_d
+ N_WL<58>_XI0/XI31/XI3/MM3_g N_BLN<12>_XI0/XI31/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM0 N_XI0/XI31/XI3/NET34_XI0/XI31/XI3/MM0_d
+ N_WL<58>_XI0/XI31/XI3/MM0_g N_BL<12>_XI0/XI31/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM1 N_XI0/XI31/XI3/NET33_XI0/XI31/XI3/MM1_d
+ N_XI0/XI31/XI3/NET34_XI0/XI31/XI3/MM1_g N_VSS_XI0/XI31/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM9 N_XI0/XI31/XI3/NET36_XI0/XI31/XI3/MM9_d
+ N_WL<59>_XI0/XI31/XI3/MM9_g N_BL<12>_XI0/XI31/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM6 N_XI0/XI31/XI3/NET35_XI0/XI31/XI3/MM6_d
+ N_XI0/XI31/XI3/NET36_XI0/XI31/XI3/MM6_g N_VSS_XI0/XI31/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM7 N_XI0/XI31/XI3/NET36_XI0/XI31/XI3/MM7_d
+ N_XI0/XI31/XI3/NET35_XI0/XI31/XI3/MM7_g N_VSS_XI0/XI31/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM8 N_XI0/XI31/XI3/NET35_XI0/XI31/XI3/MM8_d
+ N_WL<59>_XI0/XI31/XI3/MM8_g N_BLN<12>_XI0/XI31/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI3/MM5 N_XI0/XI31/XI3/NET34_XI0/XI31/XI3/MM5_d
+ N_XI0/XI31/XI3/NET33_XI0/XI31/XI3/MM5_g N_VDD_XI0/XI31/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI3/MM4 N_XI0/XI31/XI3/NET33_XI0/XI31/XI3/MM4_d
+ N_XI0/XI31/XI3/NET34_XI0/XI31/XI3/MM4_g N_VDD_XI0/XI31/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI3/MM10 N_XI0/XI31/XI3/NET35_XI0/XI31/XI3/MM10_d
+ N_XI0/XI31/XI3/NET36_XI0/XI31/XI3/MM10_g N_VDD_XI0/XI31/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI3/MM11 N_XI0/XI31/XI3/NET36_XI0/XI31/XI3/MM11_d
+ N_XI0/XI31/XI3/NET35_XI0/XI31/XI3/MM11_g N_VDD_XI0/XI31/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI4/MM2 N_XI0/XI31/XI4/NET34_XI0/XI31/XI4/MM2_d
+ N_XI0/XI31/XI4/NET33_XI0/XI31/XI4/MM2_g N_VSS_XI0/XI31/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM3 N_XI0/XI31/XI4/NET33_XI0/XI31/XI4/MM3_d
+ N_WL<58>_XI0/XI31/XI4/MM3_g N_BLN<11>_XI0/XI31/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM0 N_XI0/XI31/XI4/NET34_XI0/XI31/XI4/MM0_d
+ N_WL<58>_XI0/XI31/XI4/MM0_g N_BL<11>_XI0/XI31/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM1 N_XI0/XI31/XI4/NET33_XI0/XI31/XI4/MM1_d
+ N_XI0/XI31/XI4/NET34_XI0/XI31/XI4/MM1_g N_VSS_XI0/XI31/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM9 N_XI0/XI31/XI4/NET36_XI0/XI31/XI4/MM9_d
+ N_WL<59>_XI0/XI31/XI4/MM9_g N_BL<11>_XI0/XI31/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM6 N_XI0/XI31/XI4/NET35_XI0/XI31/XI4/MM6_d
+ N_XI0/XI31/XI4/NET36_XI0/XI31/XI4/MM6_g N_VSS_XI0/XI31/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM7 N_XI0/XI31/XI4/NET36_XI0/XI31/XI4/MM7_d
+ N_XI0/XI31/XI4/NET35_XI0/XI31/XI4/MM7_g N_VSS_XI0/XI31/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM8 N_XI0/XI31/XI4/NET35_XI0/XI31/XI4/MM8_d
+ N_WL<59>_XI0/XI31/XI4/MM8_g N_BLN<11>_XI0/XI31/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI4/MM5 N_XI0/XI31/XI4/NET34_XI0/XI31/XI4/MM5_d
+ N_XI0/XI31/XI4/NET33_XI0/XI31/XI4/MM5_g N_VDD_XI0/XI31/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI4/MM4 N_XI0/XI31/XI4/NET33_XI0/XI31/XI4/MM4_d
+ N_XI0/XI31/XI4/NET34_XI0/XI31/XI4/MM4_g N_VDD_XI0/XI31/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI4/MM10 N_XI0/XI31/XI4/NET35_XI0/XI31/XI4/MM10_d
+ N_XI0/XI31/XI4/NET36_XI0/XI31/XI4/MM10_g N_VDD_XI0/XI31/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI4/MM11 N_XI0/XI31/XI4/NET36_XI0/XI31/XI4/MM11_d
+ N_XI0/XI31/XI4/NET35_XI0/XI31/XI4/MM11_g N_VDD_XI0/XI31/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI5/MM2 N_XI0/XI31/XI5/NET34_XI0/XI31/XI5/MM2_d
+ N_XI0/XI31/XI5/NET33_XI0/XI31/XI5/MM2_g N_VSS_XI0/XI31/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM3 N_XI0/XI31/XI5/NET33_XI0/XI31/XI5/MM3_d
+ N_WL<58>_XI0/XI31/XI5/MM3_g N_BLN<10>_XI0/XI31/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM0 N_XI0/XI31/XI5/NET34_XI0/XI31/XI5/MM0_d
+ N_WL<58>_XI0/XI31/XI5/MM0_g N_BL<10>_XI0/XI31/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM1 N_XI0/XI31/XI5/NET33_XI0/XI31/XI5/MM1_d
+ N_XI0/XI31/XI5/NET34_XI0/XI31/XI5/MM1_g N_VSS_XI0/XI31/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM9 N_XI0/XI31/XI5/NET36_XI0/XI31/XI5/MM9_d
+ N_WL<59>_XI0/XI31/XI5/MM9_g N_BL<10>_XI0/XI31/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM6 N_XI0/XI31/XI5/NET35_XI0/XI31/XI5/MM6_d
+ N_XI0/XI31/XI5/NET36_XI0/XI31/XI5/MM6_g N_VSS_XI0/XI31/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM7 N_XI0/XI31/XI5/NET36_XI0/XI31/XI5/MM7_d
+ N_XI0/XI31/XI5/NET35_XI0/XI31/XI5/MM7_g N_VSS_XI0/XI31/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM8 N_XI0/XI31/XI5/NET35_XI0/XI31/XI5/MM8_d
+ N_WL<59>_XI0/XI31/XI5/MM8_g N_BLN<10>_XI0/XI31/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI5/MM5 N_XI0/XI31/XI5/NET34_XI0/XI31/XI5/MM5_d
+ N_XI0/XI31/XI5/NET33_XI0/XI31/XI5/MM5_g N_VDD_XI0/XI31/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI5/MM4 N_XI0/XI31/XI5/NET33_XI0/XI31/XI5/MM4_d
+ N_XI0/XI31/XI5/NET34_XI0/XI31/XI5/MM4_g N_VDD_XI0/XI31/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI5/MM10 N_XI0/XI31/XI5/NET35_XI0/XI31/XI5/MM10_d
+ N_XI0/XI31/XI5/NET36_XI0/XI31/XI5/MM10_g N_VDD_XI0/XI31/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI5/MM11 N_XI0/XI31/XI5/NET36_XI0/XI31/XI5/MM11_d
+ N_XI0/XI31/XI5/NET35_XI0/XI31/XI5/MM11_g N_VDD_XI0/XI31/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI6/MM2 N_XI0/XI31/XI6/NET34_XI0/XI31/XI6/MM2_d
+ N_XI0/XI31/XI6/NET33_XI0/XI31/XI6/MM2_g N_VSS_XI0/XI31/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM3 N_XI0/XI31/XI6/NET33_XI0/XI31/XI6/MM3_d
+ N_WL<58>_XI0/XI31/XI6/MM3_g N_BLN<9>_XI0/XI31/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM0 N_XI0/XI31/XI6/NET34_XI0/XI31/XI6/MM0_d
+ N_WL<58>_XI0/XI31/XI6/MM0_g N_BL<9>_XI0/XI31/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM1 N_XI0/XI31/XI6/NET33_XI0/XI31/XI6/MM1_d
+ N_XI0/XI31/XI6/NET34_XI0/XI31/XI6/MM1_g N_VSS_XI0/XI31/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM9 N_XI0/XI31/XI6/NET36_XI0/XI31/XI6/MM9_d
+ N_WL<59>_XI0/XI31/XI6/MM9_g N_BL<9>_XI0/XI31/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM6 N_XI0/XI31/XI6/NET35_XI0/XI31/XI6/MM6_d
+ N_XI0/XI31/XI6/NET36_XI0/XI31/XI6/MM6_g N_VSS_XI0/XI31/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM7 N_XI0/XI31/XI6/NET36_XI0/XI31/XI6/MM7_d
+ N_XI0/XI31/XI6/NET35_XI0/XI31/XI6/MM7_g N_VSS_XI0/XI31/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM8 N_XI0/XI31/XI6/NET35_XI0/XI31/XI6/MM8_d
+ N_WL<59>_XI0/XI31/XI6/MM8_g N_BLN<9>_XI0/XI31/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI6/MM5 N_XI0/XI31/XI6/NET34_XI0/XI31/XI6/MM5_d
+ N_XI0/XI31/XI6/NET33_XI0/XI31/XI6/MM5_g N_VDD_XI0/XI31/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI6/MM4 N_XI0/XI31/XI6/NET33_XI0/XI31/XI6/MM4_d
+ N_XI0/XI31/XI6/NET34_XI0/XI31/XI6/MM4_g N_VDD_XI0/XI31/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI6/MM10 N_XI0/XI31/XI6/NET35_XI0/XI31/XI6/MM10_d
+ N_XI0/XI31/XI6/NET36_XI0/XI31/XI6/MM10_g N_VDD_XI0/XI31/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI6/MM11 N_XI0/XI31/XI6/NET36_XI0/XI31/XI6/MM11_d
+ N_XI0/XI31/XI6/NET35_XI0/XI31/XI6/MM11_g N_VDD_XI0/XI31/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI7/MM2 N_XI0/XI31/XI7/NET34_XI0/XI31/XI7/MM2_d
+ N_XI0/XI31/XI7/NET33_XI0/XI31/XI7/MM2_g N_VSS_XI0/XI31/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM3 N_XI0/XI31/XI7/NET33_XI0/XI31/XI7/MM3_d
+ N_WL<58>_XI0/XI31/XI7/MM3_g N_BLN<8>_XI0/XI31/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM0 N_XI0/XI31/XI7/NET34_XI0/XI31/XI7/MM0_d
+ N_WL<58>_XI0/XI31/XI7/MM0_g N_BL<8>_XI0/XI31/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM1 N_XI0/XI31/XI7/NET33_XI0/XI31/XI7/MM1_d
+ N_XI0/XI31/XI7/NET34_XI0/XI31/XI7/MM1_g N_VSS_XI0/XI31/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM9 N_XI0/XI31/XI7/NET36_XI0/XI31/XI7/MM9_d
+ N_WL<59>_XI0/XI31/XI7/MM9_g N_BL<8>_XI0/XI31/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM6 N_XI0/XI31/XI7/NET35_XI0/XI31/XI7/MM6_d
+ N_XI0/XI31/XI7/NET36_XI0/XI31/XI7/MM6_g N_VSS_XI0/XI31/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM7 N_XI0/XI31/XI7/NET36_XI0/XI31/XI7/MM7_d
+ N_XI0/XI31/XI7/NET35_XI0/XI31/XI7/MM7_g N_VSS_XI0/XI31/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM8 N_XI0/XI31/XI7/NET35_XI0/XI31/XI7/MM8_d
+ N_WL<59>_XI0/XI31/XI7/MM8_g N_BLN<8>_XI0/XI31/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI7/MM5 N_XI0/XI31/XI7/NET34_XI0/XI31/XI7/MM5_d
+ N_XI0/XI31/XI7/NET33_XI0/XI31/XI7/MM5_g N_VDD_XI0/XI31/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI7/MM4 N_XI0/XI31/XI7/NET33_XI0/XI31/XI7/MM4_d
+ N_XI0/XI31/XI7/NET34_XI0/XI31/XI7/MM4_g N_VDD_XI0/XI31/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI7/MM10 N_XI0/XI31/XI7/NET35_XI0/XI31/XI7/MM10_d
+ N_XI0/XI31/XI7/NET36_XI0/XI31/XI7/MM10_g N_VDD_XI0/XI31/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI7/MM11 N_XI0/XI31/XI7/NET36_XI0/XI31/XI7/MM11_d
+ N_XI0/XI31/XI7/NET35_XI0/XI31/XI7/MM11_g N_VDD_XI0/XI31/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI8/MM2 N_XI0/XI31/XI8/NET34_XI0/XI31/XI8/MM2_d
+ N_XI0/XI31/XI8/NET33_XI0/XI31/XI8/MM2_g N_VSS_XI0/XI31/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM3 N_XI0/XI31/XI8/NET33_XI0/XI31/XI8/MM3_d
+ N_WL<58>_XI0/XI31/XI8/MM3_g N_BLN<7>_XI0/XI31/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM0 N_XI0/XI31/XI8/NET34_XI0/XI31/XI8/MM0_d
+ N_WL<58>_XI0/XI31/XI8/MM0_g N_BL<7>_XI0/XI31/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM1 N_XI0/XI31/XI8/NET33_XI0/XI31/XI8/MM1_d
+ N_XI0/XI31/XI8/NET34_XI0/XI31/XI8/MM1_g N_VSS_XI0/XI31/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM9 N_XI0/XI31/XI8/NET36_XI0/XI31/XI8/MM9_d
+ N_WL<59>_XI0/XI31/XI8/MM9_g N_BL<7>_XI0/XI31/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM6 N_XI0/XI31/XI8/NET35_XI0/XI31/XI8/MM6_d
+ N_XI0/XI31/XI8/NET36_XI0/XI31/XI8/MM6_g N_VSS_XI0/XI31/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM7 N_XI0/XI31/XI8/NET36_XI0/XI31/XI8/MM7_d
+ N_XI0/XI31/XI8/NET35_XI0/XI31/XI8/MM7_g N_VSS_XI0/XI31/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM8 N_XI0/XI31/XI8/NET35_XI0/XI31/XI8/MM8_d
+ N_WL<59>_XI0/XI31/XI8/MM8_g N_BLN<7>_XI0/XI31/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI8/MM5 N_XI0/XI31/XI8/NET34_XI0/XI31/XI8/MM5_d
+ N_XI0/XI31/XI8/NET33_XI0/XI31/XI8/MM5_g N_VDD_XI0/XI31/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI8/MM4 N_XI0/XI31/XI8/NET33_XI0/XI31/XI8/MM4_d
+ N_XI0/XI31/XI8/NET34_XI0/XI31/XI8/MM4_g N_VDD_XI0/XI31/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI8/MM10 N_XI0/XI31/XI8/NET35_XI0/XI31/XI8/MM10_d
+ N_XI0/XI31/XI8/NET36_XI0/XI31/XI8/MM10_g N_VDD_XI0/XI31/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI8/MM11 N_XI0/XI31/XI8/NET36_XI0/XI31/XI8/MM11_d
+ N_XI0/XI31/XI8/NET35_XI0/XI31/XI8/MM11_g N_VDD_XI0/XI31/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI9/MM2 N_XI0/XI31/XI9/NET34_XI0/XI31/XI9/MM2_d
+ N_XI0/XI31/XI9/NET33_XI0/XI31/XI9/MM2_g N_VSS_XI0/XI31/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM3 N_XI0/XI31/XI9/NET33_XI0/XI31/XI9/MM3_d
+ N_WL<58>_XI0/XI31/XI9/MM3_g N_BLN<6>_XI0/XI31/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM0 N_XI0/XI31/XI9/NET34_XI0/XI31/XI9/MM0_d
+ N_WL<58>_XI0/XI31/XI9/MM0_g N_BL<6>_XI0/XI31/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM1 N_XI0/XI31/XI9/NET33_XI0/XI31/XI9/MM1_d
+ N_XI0/XI31/XI9/NET34_XI0/XI31/XI9/MM1_g N_VSS_XI0/XI31/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM9 N_XI0/XI31/XI9/NET36_XI0/XI31/XI9/MM9_d
+ N_WL<59>_XI0/XI31/XI9/MM9_g N_BL<6>_XI0/XI31/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM6 N_XI0/XI31/XI9/NET35_XI0/XI31/XI9/MM6_d
+ N_XI0/XI31/XI9/NET36_XI0/XI31/XI9/MM6_g N_VSS_XI0/XI31/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM7 N_XI0/XI31/XI9/NET36_XI0/XI31/XI9/MM7_d
+ N_XI0/XI31/XI9/NET35_XI0/XI31/XI9/MM7_g N_VSS_XI0/XI31/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM8 N_XI0/XI31/XI9/NET35_XI0/XI31/XI9/MM8_d
+ N_WL<59>_XI0/XI31/XI9/MM8_g N_BLN<6>_XI0/XI31/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI9/MM5 N_XI0/XI31/XI9/NET34_XI0/XI31/XI9/MM5_d
+ N_XI0/XI31/XI9/NET33_XI0/XI31/XI9/MM5_g N_VDD_XI0/XI31/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI9/MM4 N_XI0/XI31/XI9/NET33_XI0/XI31/XI9/MM4_d
+ N_XI0/XI31/XI9/NET34_XI0/XI31/XI9/MM4_g N_VDD_XI0/XI31/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI9/MM10 N_XI0/XI31/XI9/NET35_XI0/XI31/XI9/MM10_d
+ N_XI0/XI31/XI9/NET36_XI0/XI31/XI9/MM10_g N_VDD_XI0/XI31/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI9/MM11 N_XI0/XI31/XI9/NET36_XI0/XI31/XI9/MM11_d
+ N_XI0/XI31/XI9/NET35_XI0/XI31/XI9/MM11_g N_VDD_XI0/XI31/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI10/MM2 N_XI0/XI31/XI10/NET34_XI0/XI31/XI10/MM2_d
+ N_XI0/XI31/XI10/NET33_XI0/XI31/XI10/MM2_g N_VSS_XI0/XI31/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM3 N_XI0/XI31/XI10/NET33_XI0/XI31/XI10/MM3_d
+ N_WL<58>_XI0/XI31/XI10/MM3_g N_BLN<5>_XI0/XI31/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM0 N_XI0/XI31/XI10/NET34_XI0/XI31/XI10/MM0_d
+ N_WL<58>_XI0/XI31/XI10/MM0_g N_BL<5>_XI0/XI31/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM1 N_XI0/XI31/XI10/NET33_XI0/XI31/XI10/MM1_d
+ N_XI0/XI31/XI10/NET34_XI0/XI31/XI10/MM1_g N_VSS_XI0/XI31/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM9 N_XI0/XI31/XI10/NET36_XI0/XI31/XI10/MM9_d
+ N_WL<59>_XI0/XI31/XI10/MM9_g N_BL<5>_XI0/XI31/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM6 N_XI0/XI31/XI10/NET35_XI0/XI31/XI10/MM6_d
+ N_XI0/XI31/XI10/NET36_XI0/XI31/XI10/MM6_g N_VSS_XI0/XI31/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM7 N_XI0/XI31/XI10/NET36_XI0/XI31/XI10/MM7_d
+ N_XI0/XI31/XI10/NET35_XI0/XI31/XI10/MM7_g N_VSS_XI0/XI31/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM8 N_XI0/XI31/XI10/NET35_XI0/XI31/XI10/MM8_d
+ N_WL<59>_XI0/XI31/XI10/MM8_g N_BLN<5>_XI0/XI31/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI10/MM5 N_XI0/XI31/XI10/NET34_XI0/XI31/XI10/MM5_d
+ N_XI0/XI31/XI10/NET33_XI0/XI31/XI10/MM5_g N_VDD_XI0/XI31/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI10/MM4 N_XI0/XI31/XI10/NET33_XI0/XI31/XI10/MM4_d
+ N_XI0/XI31/XI10/NET34_XI0/XI31/XI10/MM4_g N_VDD_XI0/XI31/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI10/MM10 N_XI0/XI31/XI10/NET35_XI0/XI31/XI10/MM10_d
+ N_XI0/XI31/XI10/NET36_XI0/XI31/XI10/MM10_g N_VDD_XI0/XI31/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI10/MM11 N_XI0/XI31/XI10/NET36_XI0/XI31/XI10/MM11_d
+ N_XI0/XI31/XI10/NET35_XI0/XI31/XI10/MM11_g N_VDD_XI0/XI31/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI11/MM2 N_XI0/XI31/XI11/NET34_XI0/XI31/XI11/MM2_d
+ N_XI0/XI31/XI11/NET33_XI0/XI31/XI11/MM2_g N_VSS_XI0/XI31/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM3 N_XI0/XI31/XI11/NET33_XI0/XI31/XI11/MM3_d
+ N_WL<58>_XI0/XI31/XI11/MM3_g N_BLN<4>_XI0/XI31/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM0 N_XI0/XI31/XI11/NET34_XI0/XI31/XI11/MM0_d
+ N_WL<58>_XI0/XI31/XI11/MM0_g N_BL<4>_XI0/XI31/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM1 N_XI0/XI31/XI11/NET33_XI0/XI31/XI11/MM1_d
+ N_XI0/XI31/XI11/NET34_XI0/XI31/XI11/MM1_g N_VSS_XI0/XI31/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM9 N_XI0/XI31/XI11/NET36_XI0/XI31/XI11/MM9_d
+ N_WL<59>_XI0/XI31/XI11/MM9_g N_BL<4>_XI0/XI31/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM6 N_XI0/XI31/XI11/NET35_XI0/XI31/XI11/MM6_d
+ N_XI0/XI31/XI11/NET36_XI0/XI31/XI11/MM6_g N_VSS_XI0/XI31/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM7 N_XI0/XI31/XI11/NET36_XI0/XI31/XI11/MM7_d
+ N_XI0/XI31/XI11/NET35_XI0/XI31/XI11/MM7_g N_VSS_XI0/XI31/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM8 N_XI0/XI31/XI11/NET35_XI0/XI31/XI11/MM8_d
+ N_WL<59>_XI0/XI31/XI11/MM8_g N_BLN<4>_XI0/XI31/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI11/MM5 N_XI0/XI31/XI11/NET34_XI0/XI31/XI11/MM5_d
+ N_XI0/XI31/XI11/NET33_XI0/XI31/XI11/MM5_g N_VDD_XI0/XI31/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI11/MM4 N_XI0/XI31/XI11/NET33_XI0/XI31/XI11/MM4_d
+ N_XI0/XI31/XI11/NET34_XI0/XI31/XI11/MM4_g N_VDD_XI0/XI31/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI11/MM10 N_XI0/XI31/XI11/NET35_XI0/XI31/XI11/MM10_d
+ N_XI0/XI31/XI11/NET36_XI0/XI31/XI11/MM10_g N_VDD_XI0/XI31/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI11/MM11 N_XI0/XI31/XI11/NET36_XI0/XI31/XI11/MM11_d
+ N_XI0/XI31/XI11/NET35_XI0/XI31/XI11/MM11_g N_VDD_XI0/XI31/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI12/MM2 N_XI0/XI31/XI12/NET34_XI0/XI31/XI12/MM2_d
+ N_XI0/XI31/XI12/NET33_XI0/XI31/XI12/MM2_g N_VSS_XI0/XI31/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM3 N_XI0/XI31/XI12/NET33_XI0/XI31/XI12/MM3_d
+ N_WL<58>_XI0/XI31/XI12/MM3_g N_BLN<3>_XI0/XI31/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM0 N_XI0/XI31/XI12/NET34_XI0/XI31/XI12/MM0_d
+ N_WL<58>_XI0/XI31/XI12/MM0_g N_BL<3>_XI0/XI31/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM1 N_XI0/XI31/XI12/NET33_XI0/XI31/XI12/MM1_d
+ N_XI0/XI31/XI12/NET34_XI0/XI31/XI12/MM1_g N_VSS_XI0/XI31/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM9 N_XI0/XI31/XI12/NET36_XI0/XI31/XI12/MM9_d
+ N_WL<59>_XI0/XI31/XI12/MM9_g N_BL<3>_XI0/XI31/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM6 N_XI0/XI31/XI12/NET35_XI0/XI31/XI12/MM6_d
+ N_XI0/XI31/XI12/NET36_XI0/XI31/XI12/MM6_g N_VSS_XI0/XI31/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM7 N_XI0/XI31/XI12/NET36_XI0/XI31/XI12/MM7_d
+ N_XI0/XI31/XI12/NET35_XI0/XI31/XI12/MM7_g N_VSS_XI0/XI31/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM8 N_XI0/XI31/XI12/NET35_XI0/XI31/XI12/MM8_d
+ N_WL<59>_XI0/XI31/XI12/MM8_g N_BLN<3>_XI0/XI31/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI12/MM5 N_XI0/XI31/XI12/NET34_XI0/XI31/XI12/MM5_d
+ N_XI0/XI31/XI12/NET33_XI0/XI31/XI12/MM5_g N_VDD_XI0/XI31/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI12/MM4 N_XI0/XI31/XI12/NET33_XI0/XI31/XI12/MM4_d
+ N_XI0/XI31/XI12/NET34_XI0/XI31/XI12/MM4_g N_VDD_XI0/XI31/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI12/MM10 N_XI0/XI31/XI12/NET35_XI0/XI31/XI12/MM10_d
+ N_XI0/XI31/XI12/NET36_XI0/XI31/XI12/MM10_g N_VDD_XI0/XI31/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI12/MM11 N_XI0/XI31/XI12/NET36_XI0/XI31/XI12/MM11_d
+ N_XI0/XI31/XI12/NET35_XI0/XI31/XI12/MM11_g N_VDD_XI0/XI31/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI13/MM2 N_XI0/XI31/XI13/NET34_XI0/XI31/XI13/MM2_d
+ N_XI0/XI31/XI13/NET33_XI0/XI31/XI13/MM2_g N_VSS_XI0/XI31/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM3 N_XI0/XI31/XI13/NET33_XI0/XI31/XI13/MM3_d
+ N_WL<58>_XI0/XI31/XI13/MM3_g N_BLN<2>_XI0/XI31/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM0 N_XI0/XI31/XI13/NET34_XI0/XI31/XI13/MM0_d
+ N_WL<58>_XI0/XI31/XI13/MM0_g N_BL<2>_XI0/XI31/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM1 N_XI0/XI31/XI13/NET33_XI0/XI31/XI13/MM1_d
+ N_XI0/XI31/XI13/NET34_XI0/XI31/XI13/MM1_g N_VSS_XI0/XI31/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM9 N_XI0/XI31/XI13/NET36_XI0/XI31/XI13/MM9_d
+ N_WL<59>_XI0/XI31/XI13/MM9_g N_BL<2>_XI0/XI31/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM6 N_XI0/XI31/XI13/NET35_XI0/XI31/XI13/MM6_d
+ N_XI0/XI31/XI13/NET36_XI0/XI31/XI13/MM6_g N_VSS_XI0/XI31/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM7 N_XI0/XI31/XI13/NET36_XI0/XI31/XI13/MM7_d
+ N_XI0/XI31/XI13/NET35_XI0/XI31/XI13/MM7_g N_VSS_XI0/XI31/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM8 N_XI0/XI31/XI13/NET35_XI0/XI31/XI13/MM8_d
+ N_WL<59>_XI0/XI31/XI13/MM8_g N_BLN<2>_XI0/XI31/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI13/MM5 N_XI0/XI31/XI13/NET34_XI0/XI31/XI13/MM5_d
+ N_XI0/XI31/XI13/NET33_XI0/XI31/XI13/MM5_g N_VDD_XI0/XI31/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI13/MM4 N_XI0/XI31/XI13/NET33_XI0/XI31/XI13/MM4_d
+ N_XI0/XI31/XI13/NET34_XI0/XI31/XI13/MM4_g N_VDD_XI0/XI31/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI13/MM10 N_XI0/XI31/XI13/NET35_XI0/XI31/XI13/MM10_d
+ N_XI0/XI31/XI13/NET36_XI0/XI31/XI13/MM10_g N_VDD_XI0/XI31/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI13/MM11 N_XI0/XI31/XI13/NET36_XI0/XI31/XI13/MM11_d
+ N_XI0/XI31/XI13/NET35_XI0/XI31/XI13/MM11_g N_VDD_XI0/XI31/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI14/MM2 N_XI0/XI31/XI14/NET34_XI0/XI31/XI14/MM2_d
+ N_XI0/XI31/XI14/NET33_XI0/XI31/XI14/MM2_g N_VSS_XI0/XI31/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM3 N_XI0/XI31/XI14/NET33_XI0/XI31/XI14/MM3_d
+ N_WL<58>_XI0/XI31/XI14/MM3_g N_BLN<1>_XI0/XI31/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM0 N_XI0/XI31/XI14/NET34_XI0/XI31/XI14/MM0_d
+ N_WL<58>_XI0/XI31/XI14/MM0_g N_BL<1>_XI0/XI31/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM1 N_XI0/XI31/XI14/NET33_XI0/XI31/XI14/MM1_d
+ N_XI0/XI31/XI14/NET34_XI0/XI31/XI14/MM1_g N_VSS_XI0/XI31/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM9 N_XI0/XI31/XI14/NET36_XI0/XI31/XI14/MM9_d
+ N_WL<59>_XI0/XI31/XI14/MM9_g N_BL<1>_XI0/XI31/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM6 N_XI0/XI31/XI14/NET35_XI0/XI31/XI14/MM6_d
+ N_XI0/XI31/XI14/NET36_XI0/XI31/XI14/MM6_g N_VSS_XI0/XI31/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM7 N_XI0/XI31/XI14/NET36_XI0/XI31/XI14/MM7_d
+ N_XI0/XI31/XI14/NET35_XI0/XI31/XI14/MM7_g N_VSS_XI0/XI31/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM8 N_XI0/XI31/XI14/NET35_XI0/XI31/XI14/MM8_d
+ N_WL<59>_XI0/XI31/XI14/MM8_g N_BLN<1>_XI0/XI31/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI14/MM5 N_XI0/XI31/XI14/NET34_XI0/XI31/XI14/MM5_d
+ N_XI0/XI31/XI14/NET33_XI0/XI31/XI14/MM5_g N_VDD_XI0/XI31/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI14/MM4 N_XI0/XI31/XI14/NET33_XI0/XI31/XI14/MM4_d
+ N_XI0/XI31/XI14/NET34_XI0/XI31/XI14/MM4_g N_VDD_XI0/XI31/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI14/MM10 N_XI0/XI31/XI14/NET35_XI0/XI31/XI14/MM10_d
+ N_XI0/XI31/XI14/NET36_XI0/XI31/XI14/MM10_g N_VDD_XI0/XI31/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI14/MM11 N_XI0/XI31/XI14/NET36_XI0/XI31/XI14/MM11_d
+ N_XI0/XI31/XI14/NET35_XI0/XI31/XI14/MM11_g N_VDD_XI0/XI31/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI15/MM2 N_XI0/XI31/XI15/NET34_XI0/XI31/XI15/MM2_d
+ N_XI0/XI31/XI15/NET33_XI0/XI31/XI15/MM2_g N_VSS_XI0/XI31/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM3 N_XI0/XI31/XI15/NET33_XI0/XI31/XI15/MM3_d
+ N_WL<58>_XI0/XI31/XI15/MM3_g N_BLN<0>_XI0/XI31/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM0 N_XI0/XI31/XI15/NET34_XI0/XI31/XI15/MM0_d
+ N_WL<58>_XI0/XI31/XI15/MM0_g N_BL<0>_XI0/XI31/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM1 N_XI0/XI31/XI15/NET33_XI0/XI31/XI15/MM1_d
+ N_XI0/XI31/XI15/NET34_XI0/XI31/XI15/MM1_g N_VSS_XI0/XI31/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM9 N_XI0/XI31/XI15/NET36_XI0/XI31/XI15/MM9_d
+ N_WL<59>_XI0/XI31/XI15/MM9_g N_BL<0>_XI0/XI31/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM6 N_XI0/XI31/XI15/NET35_XI0/XI31/XI15/MM6_d
+ N_XI0/XI31/XI15/NET36_XI0/XI31/XI15/MM6_g N_VSS_XI0/XI31/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM7 N_XI0/XI31/XI15/NET36_XI0/XI31/XI15/MM7_d
+ N_XI0/XI31/XI15/NET35_XI0/XI31/XI15/MM7_g N_VSS_XI0/XI31/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM8 N_XI0/XI31/XI15/NET35_XI0/XI31/XI15/MM8_d
+ N_WL<59>_XI0/XI31/XI15/MM8_g N_BLN<0>_XI0/XI31/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI31/XI15/MM5 N_XI0/XI31/XI15/NET34_XI0/XI31/XI15/MM5_d
+ N_XI0/XI31/XI15/NET33_XI0/XI31/XI15/MM5_g N_VDD_XI0/XI31/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI15/MM4 N_XI0/XI31/XI15/NET33_XI0/XI31/XI15/MM4_d
+ N_XI0/XI31/XI15/NET34_XI0/XI31/XI15/MM4_g N_VDD_XI0/XI31/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI15/MM10 N_XI0/XI31/XI15/NET35_XI0/XI31/XI15/MM10_d
+ N_XI0/XI31/XI15/NET36_XI0/XI31/XI15/MM10_g N_VDD_XI0/XI31/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI31/XI15/MM11 N_XI0/XI31/XI15/NET36_XI0/XI31/XI15/MM11_d
+ N_XI0/XI31/XI15/NET35_XI0/XI31/XI15/MM11_g N_VDD_XI0/XI31/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI0/MM2 N_XI0/XI32/XI0/NET34_XI0/XI32/XI0/MM2_d
+ N_XI0/XI32/XI0/NET33_XI0/XI32/XI0/MM2_g N_VSS_XI0/XI32/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM3 N_XI0/XI32/XI0/NET33_XI0/XI32/XI0/MM3_d
+ N_WL<60>_XI0/XI32/XI0/MM3_g N_BLN<15>_XI0/XI32/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM0 N_XI0/XI32/XI0/NET34_XI0/XI32/XI0/MM0_d
+ N_WL<60>_XI0/XI32/XI0/MM0_g N_BL<15>_XI0/XI32/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM1 N_XI0/XI32/XI0/NET33_XI0/XI32/XI0/MM1_d
+ N_XI0/XI32/XI0/NET34_XI0/XI32/XI0/MM1_g N_VSS_XI0/XI32/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM9 N_XI0/XI32/XI0/NET36_XI0/XI32/XI0/MM9_d
+ N_WL<61>_XI0/XI32/XI0/MM9_g N_BL<15>_XI0/XI32/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM6 N_XI0/XI32/XI0/NET35_XI0/XI32/XI0/MM6_d
+ N_XI0/XI32/XI0/NET36_XI0/XI32/XI0/MM6_g N_VSS_XI0/XI32/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM7 N_XI0/XI32/XI0/NET36_XI0/XI32/XI0/MM7_d
+ N_XI0/XI32/XI0/NET35_XI0/XI32/XI0/MM7_g N_VSS_XI0/XI32/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM8 N_XI0/XI32/XI0/NET35_XI0/XI32/XI0/MM8_d
+ N_WL<61>_XI0/XI32/XI0/MM8_g N_BLN<15>_XI0/XI32/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI0/MM5 N_XI0/XI32/XI0/NET34_XI0/XI32/XI0/MM5_d
+ N_XI0/XI32/XI0/NET33_XI0/XI32/XI0/MM5_g N_VDD_XI0/XI32/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI0/MM4 N_XI0/XI32/XI0/NET33_XI0/XI32/XI0/MM4_d
+ N_XI0/XI32/XI0/NET34_XI0/XI32/XI0/MM4_g N_VDD_XI0/XI32/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI0/MM10 N_XI0/XI32/XI0/NET35_XI0/XI32/XI0/MM10_d
+ N_XI0/XI32/XI0/NET36_XI0/XI32/XI0/MM10_g N_VDD_XI0/XI32/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI0/MM11 N_XI0/XI32/XI0/NET36_XI0/XI32/XI0/MM11_d
+ N_XI0/XI32/XI0/NET35_XI0/XI32/XI0/MM11_g N_VDD_XI0/XI32/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI1/MM2 N_XI0/XI32/XI1/NET34_XI0/XI32/XI1/MM2_d
+ N_XI0/XI32/XI1/NET33_XI0/XI32/XI1/MM2_g N_VSS_XI0/XI32/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM3 N_XI0/XI32/XI1/NET33_XI0/XI32/XI1/MM3_d
+ N_WL<60>_XI0/XI32/XI1/MM3_g N_BLN<14>_XI0/XI32/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM0 N_XI0/XI32/XI1/NET34_XI0/XI32/XI1/MM0_d
+ N_WL<60>_XI0/XI32/XI1/MM0_g N_BL<14>_XI0/XI32/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM1 N_XI0/XI32/XI1/NET33_XI0/XI32/XI1/MM1_d
+ N_XI0/XI32/XI1/NET34_XI0/XI32/XI1/MM1_g N_VSS_XI0/XI32/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM9 N_XI0/XI32/XI1/NET36_XI0/XI32/XI1/MM9_d
+ N_WL<61>_XI0/XI32/XI1/MM9_g N_BL<14>_XI0/XI32/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM6 N_XI0/XI32/XI1/NET35_XI0/XI32/XI1/MM6_d
+ N_XI0/XI32/XI1/NET36_XI0/XI32/XI1/MM6_g N_VSS_XI0/XI32/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM7 N_XI0/XI32/XI1/NET36_XI0/XI32/XI1/MM7_d
+ N_XI0/XI32/XI1/NET35_XI0/XI32/XI1/MM7_g N_VSS_XI0/XI32/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM8 N_XI0/XI32/XI1/NET35_XI0/XI32/XI1/MM8_d
+ N_WL<61>_XI0/XI32/XI1/MM8_g N_BLN<14>_XI0/XI32/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI1/MM5 N_XI0/XI32/XI1/NET34_XI0/XI32/XI1/MM5_d
+ N_XI0/XI32/XI1/NET33_XI0/XI32/XI1/MM5_g N_VDD_XI0/XI32/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI1/MM4 N_XI0/XI32/XI1/NET33_XI0/XI32/XI1/MM4_d
+ N_XI0/XI32/XI1/NET34_XI0/XI32/XI1/MM4_g N_VDD_XI0/XI32/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI1/MM10 N_XI0/XI32/XI1/NET35_XI0/XI32/XI1/MM10_d
+ N_XI0/XI32/XI1/NET36_XI0/XI32/XI1/MM10_g N_VDD_XI0/XI32/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI1/MM11 N_XI0/XI32/XI1/NET36_XI0/XI32/XI1/MM11_d
+ N_XI0/XI32/XI1/NET35_XI0/XI32/XI1/MM11_g N_VDD_XI0/XI32/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI2/MM2 N_XI0/XI32/XI2/NET34_XI0/XI32/XI2/MM2_d
+ N_XI0/XI32/XI2/NET33_XI0/XI32/XI2/MM2_g N_VSS_XI0/XI32/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM3 N_XI0/XI32/XI2/NET33_XI0/XI32/XI2/MM3_d
+ N_WL<60>_XI0/XI32/XI2/MM3_g N_BLN<13>_XI0/XI32/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM0 N_XI0/XI32/XI2/NET34_XI0/XI32/XI2/MM0_d
+ N_WL<60>_XI0/XI32/XI2/MM0_g N_BL<13>_XI0/XI32/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM1 N_XI0/XI32/XI2/NET33_XI0/XI32/XI2/MM1_d
+ N_XI0/XI32/XI2/NET34_XI0/XI32/XI2/MM1_g N_VSS_XI0/XI32/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM9 N_XI0/XI32/XI2/NET36_XI0/XI32/XI2/MM9_d
+ N_WL<61>_XI0/XI32/XI2/MM9_g N_BL<13>_XI0/XI32/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM6 N_XI0/XI32/XI2/NET35_XI0/XI32/XI2/MM6_d
+ N_XI0/XI32/XI2/NET36_XI0/XI32/XI2/MM6_g N_VSS_XI0/XI32/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM7 N_XI0/XI32/XI2/NET36_XI0/XI32/XI2/MM7_d
+ N_XI0/XI32/XI2/NET35_XI0/XI32/XI2/MM7_g N_VSS_XI0/XI32/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM8 N_XI0/XI32/XI2/NET35_XI0/XI32/XI2/MM8_d
+ N_WL<61>_XI0/XI32/XI2/MM8_g N_BLN<13>_XI0/XI32/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI2/MM5 N_XI0/XI32/XI2/NET34_XI0/XI32/XI2/MM5_d
+ N_XI0/XI32/XI2/NET33_XI0/XI32/XI2/MM5_g N_VDD_XI0/XI32/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI2/MM4 N_XI0/XI32/XI2/NET33_XI0/XI32/XI2/MM4_d
+ N_XI0/XI32/XI2/NET34_XI0/XI32/XI2/MM4_g N_VDD_XI0/XI32/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI2/MM10 N_XI0/XI32/XI2/NET35_XI0/XI32/XI2/MM10_d
+ N_XI0/XI32/XI2/NET36_XI0/XI32/XI2/MM10_g N_VDD_XI0/XI32/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI2/MM11 N_XI0/XI32/XI2/NET36_XI0/XI32/XI2/MM11_d
+ N_XI0/XI32/XI2/NET35_XI0/XI32/XI2/MM11_g N_VDD_XI0/XI32/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI3/MM2 N_XI0/XI32/XI3/NET34_XI0/XI32/XI3/MM2_d
+ N_XI0/XI32/XI3/NET33_XI0/XI32/XI3/MM2_g N_VSS_XI0/XI32/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM3 N_XI0/XI32/XI3/NET33_XI0/XI32/XI3/MM3_d
+ N_WL<60>_XI0/XI32/XI3/MM3_g N_BLN<12>_XI0/XI32/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM0 N_XI0/XI32/XI3/NET34_XI0/XI32/XI3/MM0_d
+ N_WL<60>_XI0/XI32/XI3/MM0_g N_BL<12>_XI0/XI32/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM1 N_XI0/XI32/XI3/NET33_XI0/XI32/XI3/MM1_d
+ N_XI0/XI32/XI3/NET34_XI0/XI32/XI3/MM1_g N_VSS_XI0/XI32/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM9 N_XI0/XI32/XI3/NET36_XI0/XI32/XI3/MM9_d
+ N_WL<61>_XI0/XI32/XI3/MM9_g N_BL<12>_XI0/XI32/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM6 N_XI0/XI32/XI3/NET35_XI0/XI32/XI3/MM6_d
+ N_XI0/XI32/XI3/NET36_XI0/XI32/XI3/MM6_g N_VSS_XI0/XI32/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM7 N_XI0/XI32/XI3/NET36_XI0/XI32/XI3/MM7_d
+ N_XI0/XI32/XI3/NET35_XI0/XI32/XI3/MM7_g N_VSS_XI0/XI32/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM8 N_XI0/XI32/XI3/NET35_XI0/XI32/XI3/MM8_d
+ N_WL<61>_XI0/XI32/XI3/MM8_g N_BLN<12>_XI0/XI32/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI3/MM5 N_XI0/XI32/XI3/NET34_XI0/XI32/XI3/MM5_d
+ N_XI0/XI32/XI3/NET33_XI0/XI32/XI3/MM5_g N_VDD_XI0/XI32/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI3/MM4 N_XI0/XI32/XI3/NET33_XI0/XI32/XI3/MM4_d
+ N_XI0/XI32/XI3/NET34_XI0/XI32/XI3/MM4_g N_VDD_XI0/XI32/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI3/MM10 N_XI0/XI32/XI3/NET35_XI0/XI32/XI3/MM10_d
+ N_XI0/XI32/XI3/NET36_XI0/XI32/XI3/MM10_g N_VDD_XI0/XI32/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI3/MM11 N_XI0/XI32/XI3/NET36_XI0/XI32/XI3/MM11_d
+ N_XI0/XI32/XI3/NET35_XI0/XI32/XI3/MM11_g N_VDD_XI0/XI32/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI4/MM2 N_XI0/XI32/XI4/NET34_XI0/XI32/XI4/MM2_d
+ N_XI0/XI32/XI4/NET33_XI0/XI32/XI4/MM2_g N_VSS_XI0/XI32/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM3 N_XI0/XI32/XI4/NET33_XI0/XI32/XI4/MM3_d
+ N_WL<60>_XI0/XI32/XI4/MM3_g N_BLN<11>_XI0/XI32/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM0 N_XI0/XI32/XI4/NET34_XI0/XI32/XI4/MM0_d
+ N_WL<60>_XI0/XI32/XI4/MM0_g N_BL<11>_XI0/XI32/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM1 N_XI0/XI32/XI4/NET33_XI0/XI32/XI4/MM1_d
+ N_XI0/XI32/XI4/NET34_XI0/XI32/XI4/MM1_g N_VSS_XI0/XI32/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM9 N_XI0/XI32/XI4/NET36_XI0/XI32/XI4/MM9_d
+ N_WL<61>_XI0/XI32/XI4/MM9_g N_BL<11>_XI0/XI32/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM6 N_XI0/XI32/XI4/NET35_XI0/XI32/XI4/MM6_d
+ N_XI0/XI32/XI4/NET36_XI0/XI32/XI4/MM6_g N_VSS_XI0/XI32/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM7 N_XI0/XI32/XI4/NET36_XI0/XI32/XI4/MM7_d
+ N_XI0/XI32/XI4/NET35_XI0/XI32/XI4/MM7_g N_VSS_XI0/XI32/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM8 N_XI0/XI32/XI4/NET35_XI0/XI32/XI4/MM8_d
+ N_WL<61>_XI0/XI32/XI4/MM8_g N_BLN<11>_XI0/XI32/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI4/MM5 N_XI0/XI32/XI4/NET34_XI0/XI32/XI4/MM5_d
+ N_XI0/XI32/XI4/NET33_XI0/XI32/XI4/MM5_g N_VDD_XI0/XI32/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI4/MM4 N_XI0/XI32/XI4/NET33_XI0/XI32/XI4/MM4_d
+ N_XI0/XI32/XI4/NET34_XI0/XI32/XI4/MM4_g N_VDD_XI0/XI32/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI4/MM10 N_XI0/XI32/XI4/NET35_XI0/XI32/XI4/MM10_d
+ N_XI0/XI32/XI4/NET36_XI0/XI32/XI4/MM10_g N_VDD_XI0/XI32/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI4/MM11 N_XI0/XI32/XI4/NET36_XI0/XI32/XI4/MM11_d
+ N_XI0/XI32/XI4/NET35_XI0/XI32/XI4/MM11_g N_VDD_XI0/XI32/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI5/MM2 N_XI0/XI32/XI5/NET34_XI0/XI32/XI5/MM2_d
+ N_XI0/XI32/XI5/NET33_XI0/XI32/XI5/MM2_g N_VSS_XI0/XI32/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM3 N_XI0/XI32/XI5/NET33_XI0/XI32/XI5/MM3_d
+ N_WL<60>_XI0/XI32/XI5/MM3_g N_BLN<10>_XI0/XI32/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM0 N_XI0/XI32/XI5/NET34_XI0/XI32/XI5/MM0_d
+ N_WL<60>_XI0/XI32/XI5/MM0_g N_BL<10>_XI0/XI32/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM1 N_XI0/XI32/XI5/NET33_XI0/XI32/XI5/MM1_d
+ N_XI0/XI32/XI5/NET34_XI0/XI32/XI5/MM1_g N_VSS_XI0/XI32/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM9 N_XI0/XI32/XI5/NET36_XI0/XI32/XI5/MM9_d
+ N_WL<61>_XI0/XI32/XI5/MM9_g N_BL<10>_XI0/XI32/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM6 N_XI0/XI32/XI5/NET35_XI0/XI32/XI5/MM6_d
+ N_XI0/XI32/XI5/NET36_XI0/XI32/XI5/MM6_g N_VSS_XI0/XI32/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM7 N_XI0/XI32/XI5/NET36_XI0/XI32/XI5/MM7_d
+ N_XI0/XI32/XI5/NET35_XI0/XI32/XI5/MM7_g N_VSS_XI0/XI32/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM8 N_XI0/XI32/XI5/NET35_XI0/XI32/XI5/MM8_d
+ N_WL<61>_XI0/XI32/XI5/MM8_g N_BLN<10>_XI0/XI32/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI5/MM5 N_XI0/XI32/XI5/NET34_XI0/XI32/XI5/MM5_d
+ N_XI0/XI32/XI5/NET33_XI0/XI32/XI5/MM5_g N_VDD_XI0/XI32/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI5/MM4 N_XI0/XI32/XI5/NET33_XI0/XI32/XI5/MM4_d
+ N_XI0/XI32/XI5/NET34_XI0/XI32/XI5/MM4_g N_VDD_XI0/XI32/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI5/MM10 N_XI0/XI32/XI5/NET35_XI0/XI32/XI5/MM10_d
+ N_XI0/XI32/XI5/NET36_XI0/XI32/XI5/MM10_g N_VDD_XI0/XI32/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI5/MM11 N_XI0/XI32/XI5/NET36_XI0/XI32/XI5/MM11_d
+ N_XI0/XI32/XI5/NET35_XI0/XI32/XI5/MM11_g N_VDD_XI0/XI32/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI6/MM2 N_XI0/XI32/XI6/NET34_XI0/XI32/XI6/MM2_d
+ N_XI0/XI32/XI6/NET33_XI0/XI32/XI6/MM2_g N_VSS_XI0/XI32/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM3 N_XI0/XI32/XI6/NET33_XI0/XI32/XI6/MM3_d
+ N_WL<60>_XI0/XI32/XI6/MM3_g N_BLN<9>_XI0/XI32/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM0 N_XI0/XI32/XI6/NET34_XI0/XI32/XI6/MM0_d
+ N_WL<60>_XI0/XI32/XI6/MM0_g N_BL<9>_XI0/XI32/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM1 N_XI0/XI32/XI6/NET33_XI0/XI32/XI6/MM1_d
+ N_XI0/XI32/XI6/NET34_XI0/XI32/XI6/MM1_g N_VSS_XI0/XI32/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM9 N_XI0/XI32/XI6/NET36_XI0/XI32/XI6/MM9_d
+ N_WL<61>_XI0/XI32/XI6/MM9_g N_BL<9>_XI0/XI32/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM6 N_XI0/XI32/XI6/NET35_XI0/XI32/XI6/MM6_d
+ N_XI0/XI32/XI6/NET36_XI0/XI32/XI6/MM6_g N_VSS_XI0/XI32/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM7 N_XI0/XI32/XI6/NET36_XI0/XI32/XI6/MM7_d
+ N_XI0/XI32/XI6/NET35_XI0/XI32/XI6/MM7_g N_VSS_XI0/XI32/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM8 N_XI0/XI32/XI6/NET35_XI0/XI32/XI6/MM8_d
+ N_WL<61>_XI0/XI32/XI6/MM8_g N_BLN<9>_XI0/XI32/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI6/MM5 N_XI0/XI32/XI6/NET34_XI0/XI32/XI6/MM5_d
+ N_XI0/XI32/XI6/NET33_XI0/XI32/XI6/MM5_g N_VDD_XI0/XI32/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI6/MM4 N_XI0/XI32/XI6/NET33_XI0/XI32/XI6/MM4_d
+ N_XI0/XI32/XI6/NET34_XI0/XI32/XI6/MM4_g N_VDD_XI0/XI32/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI6/MM10 N_XI0/XI32/XI6/NET35_XI0/XI32/XI6/MM10_d
+ N_XI0/XI32/XI6/NET36_XI0/XI32/XI6/MM10_g N_VDD_XI0/XI32/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI6/MM11 N_XI0/XI32/XI6/NET36_XI0/XI32/XI6/MM11_d
+ N_XI0/XI32/XI6/NET35_XI0/XI32/XI6/MM11_g N_VDD_XI0/XI32/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI7/MM2 N_XI0/XI32/XI7/NET34_XI0/XI32/XI7/MM2_d
+ N_XI0/XI32/XI7/NET33_XI0/XI32/XI7/MM2_g N_VSS_XI0/XI32/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM3 N_XI0/XI32/XI7/NET33_XI0/XI32/XI7/MM3_d
+ N_WL<60>_XI0/XI32/XI7/MM3_g N_BLN<8>_XI0/XI32/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM0 N_XI0/XI32/XI7/NET34_XI0/XI32/XI7/MM0_d
+ N_WL<60>_XI0/XI32/XI7/MM0_g N_BL<8>_XI0/XI32/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM1 N_XI0/XI32/XI7/NET33_XI0/XI32/XI7/MM1_d
+ N_XI0/XI32/XI7/NET34_XI0/XI32/XI7/MM1_g N_VSS_XI0/XI32/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM9 N_XI0/XI32/XI7/NET36_XI0/XI32/XI7/MM9_d
+ N_WL<61>_XI0/XI32/XI7/MM9_g N_BL<8>_XI0/XI32/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM6 N_XI0/XI32/XI7/NET35_XI0/XI32/XI7/MM6_d
+ N_XI0/XI32/XI7/NET36_XI0/XI32/XI7/MM6_g N_VSS_XI0/XI32/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM7 N_XI0/XI32/XI7/NET36_XI0/XI32/XI7/MM7_d
+ N_XI0/XI32/XI7/NET35_XI0/XI32/XI7/MM7_g N_VSS_XI0/XI32/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM8 N_XI0/XI32/XI7/NET35_XI0/XI32/XI7/MM8_d
+ N_WL<61>_XI0/XI32/XI7/MM8_g N_BLN<8>_XI0/XI32/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI7/MM5 N_XI0/XI32/XI7/NET34_XI0/XI32/XI7/MM5_d
+ N_XI0/XI32/XI7/NET33_XI0/XI32/XI7/MM5_g N_VDD_XI0/XI32/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI7/MM4 N_XI0/XI32/XI7/NET33_XI0/XI32/XI7/MM4_d
+ N_XI0/XI32/XI7/NET34_XI0/XI32/XI7/MM4_g N_VDD_XI0/XI32/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI7/MM10 N_XI0/XI32/XI7/NET35_XI0/XI32/XI7/MM10_d
+ N_XI0/XI32/XI7/NET36_XI0/XI32/XI7/MM10_g N_VDD_XI0/XI32/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI7/MM11 N_XI0/XI32/XI7/NET36_XI0/XI32/XI7/MM11_d
+ N_XI0/XI32/XI7/NET35_XI0/XI32/XI7/MM11_g N_VDD_XI0/XI32/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI8/MM2 N_XI0/XI32/XI8/NET34_XI0/XI32/XI8/MM2_d
+ N_XI0/XI32/XI8/NET33_XI0/XI32/XI8/MM2_g N_VSS_XI0/XI32/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM3 N_XI0/XI32/XI8/NET33_XI0/XI32/XI8/MM3_d
+ N_WL<60>_XI0/XI32/XI8/MM3_g N_BLN<7>_XI0/XI32/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM0 N_XI0/XI32/XI8/NET34_XI0/XI32/XI8/MM0_d
+ N_WL<60>_XI0/XI32/XI8/MM0_g N_BL<7>_XI0/XI32/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM1 N_XI0/XI32/XI8/NET33_XI0/XI32/XI8/MM1_d
+ N_XI0/XI32/XI8/NET34_XI0/XI32/XI8/MM1_g N_VSS_XI0/XI32/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM9 N_XI0/XI32/XI8/NET36_XI0/XI32/XI8/MM9_d
+ N_WL<61>_XI0/XI32/XI8/MM9_g N_BL<7>_XI0/XI32/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM6 N_XI0/XI32/XI8/NET35_XI0/XI32/XI8/MM6_d
+ N_XI0/XI32/XI8/NET36_XI0/XI32/XI8/MM6_g N_VSS_XI0/XI32/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM7 N_XI0/XI32/XI8/NET36_XI0/XI32/XI8/MM7_d
+ N_XI0/XI32/XI8/NET35_XI0/XI32/XI8/MM7_g N_VSS_XI0/XI32/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM8 N_XI0/XI32/XI8/NET35_XI0/XI32/XI8/MM8_d
+ N_WL<61>_XI0/XI32/XI8/MM8_g N_BLN<7>_XI0/XI32/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI8/MM5 N_XI0/XI32/XI8/NET34_XI0/XI32/XI8/MM5_d
+ N_XI0/XI32/XI8/NET33_XI0/XI32/XI8/MM5_g N_VDD_XI0/XI32/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI8/MM4 N_XI0/XI32/XI8/NET33_XI0/XI32/XI8/MM4_d
+ N_XI0/XI32/XI8/NET34_XI0/XI32/XI8/MM4_g N_VDD_XI0/XI32/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI8/MM10 N_XI0/XI32/XI8/NET35_XI0/XI32/XI8/MM10_d
+ N_XI0/XI32/XI8/NET36_XI0/XI32/XI8/MM10_g N_VDD_XI0/XI32/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI8/MM11 N_XI0/XI32/XI8/NET36_XI0/XI32/XI8/MM11_d
+ N_XI0/XI32/XI8/NET35_XI0/XI32/XI8/MM11_g N_VDD_XI0/XI32/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI9/MM2 N_XI0/XI32/XI9/NET34_XI0/XI32/XI9/MM2_d
+ N_XI0/XI32/XI9/NET33_XI0/XI32/XI9/MM2_g N_VSS_XI0/XI32/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM3 N_XI0/XI32/XI9/NET33_XI0/XI32/XI9/MM3_d
+ N_WL<60>_XI0/XI32/XI9/MM3_g N_BLN<6>_XI0/XI32/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM0 N_XI0/XI32/XI9/NET34_XI0/XI32/XI9/MM0_d
+ N_WL<60>_XI0/XI32/XI9/MM0_g N_BL<6>_XI0/XI32/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM1 N_XI0/XI32/XI9/NET33_XI0/XI32/XI9/MM1_d
+ N_XI0/XI32/XI9/NET34_XI0/XI32/XI9/MM1_g N_VSS_XI0/XI32/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM9 N_XI0/XI32/XI9/NET36_XI0/XI32/XI9/MM9_d
+ N_WL<61>_XI0/XI32/XI9/MM9_g N_BL<6>_XI0/XI32/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM6 N_XI0/XI32/XI9/NET35_XI0/XI32/XI9/MM6_d
+ N_XI0/XI32/XI9/NET36_XI0/XI32/XI9/MM6_g N_VSS_XI0/XI32/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM7 N_XI0/XI32/XI9/NET36_XI0/XI32/XI9/MM7_d
+ N_XI0/XI32/XI9/NET35_XI0/XI32/XI9/MM7_g N_VSS_XI0/XI32/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM8 N_XI0/XI32/XI9/NET35_XI0/XI32/XI9/MM8_d
+ N_WL<61>_XI0/XI32/XI9/MM8_g N_BLN<6>_XI0/XI32/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI9/MM5 N_XI0/XI32/XI9/NET34_XI0/XI32/XI9/MM5_d
+ N_XI0/XI32/XI9/NET33_XI0/XI32/XI9/MM5_g N_VDD_XI0/XI32/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI9/MM4 N_XI0/XI32/XI9/NET33_XI0/XI32/XI9/MM4_d
+ N_XI0/XI32/XI9/NET34_XI0/XI32/XI9/MM4_g N_VDD_XI0/XI32/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI9/MM10 N_XI0/XI32/XI9/NET35_XI0/XI32/XI9/MM10_d
+ N_XI0/XI32/XI9/NET36_XI0/XI32/XI9/MM10_g N_VDD_XI0/XI32/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI9/MM11 N_XI0/XI32/XI9/NET36_XI0/XI32/XI9/MM11_d
+ N_XI0/XI32/XI9/NET35_XI0/XI32/XI9/MM11_g N_VDD_XI0/XI32/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI10/MM2 N_XI0/XI32/XI10/NET34_XI0/XI32/XI10/MM2_d
+ N_XI0/XI32/XI10/NET33_XI0/XI32/XI10/MM2_g N_VSS_XI0/XI32/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM3 N_XI0/XI32/XI10/NET33_XI0/XI32/XI10/MM3_d
+ N_WL<60>_XI0/XI32/XI10/MM3_g N_BLN<5>_XI0/XI32/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM0 N_XI0/XI32/XI10/NET34_XI0/XI32/XI10/MM0_d
+ N_WL<60>_XI0/XI32/XI10/MM0_g N_BL<5>_XI0/XI32/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM1 N_XI0/XI32/XI10/NET33_XI0/XI32/XI10/MM1_d
+ N_XI0/XI32/XI10/NET34_XI0/XI32/XI10/MM1_g N_VSS_XI0/XI32/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM9 N_XI0/XI32/XI10/NET36_XI0/XI32/XI10/MM9_d
+ N_WL<61>_XI0/XI32/XI10/MM9_g N_BL<5>_XI0/XI32/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM6 N_XI0/XI32/XI10/NET35_XI0/XI32/XI10/MM6_d
+ N_XI0/XI32/XI10/NET36_XI0/XI32/XI10/MM6_g N_VSS_XI0/XI32/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM7 N_XI0/XI32/XI10/NET36_XI0/XI32/XI10/MM7_d
+ N_XI0/XI32/XI10/NET35_XI0/XI32/XI10/MM7_g N_VSS_XI0/XI32/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM8 N_XI0/XI32/XI10/NET35_XI0/XI32/XI10/MM8_d
+ N_WL<61>_XI0/XI32/XI10/MM8_g N_BLN<5>_XI0/XI32/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI10/MM5 N_XI0/XI32/XI10/NET34_XI0/XI32/XI10/MM5_d
+ N_XI0/XI32/XI10/NET33_XI0/XI32/XI10/MM5_g N_VDD_XI0/XI32/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI10/MM4 N_XI0/XI32/XI10/NET33_XI0/XI32/XI10/MM4_d
+ N_XI0/XI32/XI10/NET34_XI0/XI32/XI10/MM4_g N_VDD_XI0/XI32/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI10/MM10 N_XI0/XI32/XI10/NET35_XI0/XI32/XI10/MM10_d
+ N_XI0/XI32/XI10/NET36_XI0/XI32/XI10/MM10_g N_VDD_XI0/XI32/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI10/MM11 N_XI0/XI32/XI10/NET36_XI0/XI32/XI10/MM11_d
+ N_XI0/XI32/XI10/NET35_XI0/XI32/XI10/MM11_g N_VDD_XI0/XI32/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI11/MM2 N_XI0/XI32/XI11/NET34_XI0/XI32/XI11/MM2_d
+ N_XI0/XI32/XI11/NET33_XI0/XI32/XI11/MM2_g N_VSS_XI0/XI32/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM3 N_XI0/XI32/XI11/NET33_XI0/XI32/XI11/MM3_d
+ N_WL<60>_XI0/XI32/XI11/MM3_g N_BLN<4>_XI0/XI32/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM0 N_XI0/XI32/XI11/NET34_XI0/XI32/XI11/MM0_d
+ N_WL<60>_XI0/XI32/XI11/MM0_g N_BL<4>_XI0/XI32/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM1 N_XI0/XI32/XI11/NET33_XI0/XI32/XI11/MM1_d
+ N_XI0/XI32/XI11/NET34_XI0/XI32/XI11/MM1_g N_VSS_XI0/XI32/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM9 N_XI0/XI32/XI11/NET36_XI0/XI32/XI11/MM9_d
+ N_WL<61>_XI0/XI32/XI11/MM9_g N_BL<4>_XI0/XI32/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM6 N_XI0/XI32/XI11/NET35_XI0/XI32/XI11/MM6_d
+ N_XI0/XI32/XI11/NET36_XI0/XI32/XI11/MM6_g N_VSS_XI0/XI32/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM7 N_XI0/XI32/XI11/NET36_XI0/XI32/XI11/MM7_d
+ N_XI0/XI32/XI11/NET35_XI0/XI32/XI11/MM7_g N_VSS_XI0/XI32/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM8 N_XI0/XI32/XI11/NET35_XI0/XI32/XI11/MM8_d
+ N_WL<61>_XI0/XI32/XI11/MM8_g N_BLN<4>_XI0/XI32/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI11/MM5 N_XI0/XI32/XI11/NET34_XI0/XI32/XI11/MM5_d
+ N_XI0/XI32/XI11/NET33_XI0/XI32/XI11/MM5_g N_VDD_XI0/XI32/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI11/MM4 N_XI0/XI32/XI11/NET33_XI0/XI32/XI11/MM4_d
+ N_XI0/XI32/XI11/NET34_XI0/XI32/XI11/MM4_g N_VDD_XI0/XI32/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI11/MM10 N_XI0/XI32/XI11/NET35_XI0/XI32/XI11/MM10_d
+ N_XI0/XI32/XI11/NET36_XI0/XI32/XI11/MM10_g N_VDD_XI0/XI32/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI11/MM11 N_XI0/XI32/XI11/NET36_XI0/XI32/XI11/MM11_d
+ N_XI0/XI32/XI11/NET35_XI0/XI32/XI11/MM11_g N_VDD_XI0/XI32/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI12/MM2 N_XI0/XI32/XI12/NET34_XI0/XI32/XI12/MM2_d
+ N_XI0/XI32/XI12/NET33_XI0/XI32/XI12/MM2_g N_VSS_XI0/XI32/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM3 N_XI0/XI32/XI12/NET33_XI0/XI32/XI12/MM3_d
+ N_WL<60>_XI0/XI32/XI12/MM3_g N_BLN<3>_XI0/XI32/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM0 N_XI0/XI32/XI12/NET34_XI0/XI32/XI12/MM0_d
+ N_WL<60>_XI0/XI32/XI12/MM0_g N_BL<3>_XI0/XI32/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM1 N_XI0/XI32/XI12/NET33_XI0/XI32/XI12/MM1_d
+ N_XI0/XI32/XI12/NET34_XI0/XI32/XI12/MM1_g N_VSS_XI0/XI32/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM9 N_XI0/XI32/XI12/NET36_XI0/XI32/XI12/MM9_d
+ N_WL<61>_XI0/XI32/XI12/MM9_g N_BL<3>_XI0/XI32/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM6 N_XI0/XI32/XI12/NET35_XI0/XI32/XI12/MM6_d
+ N_XI0/XI32/XI12/NET36_XI0/XI32/XI12/MM6_g N_VSS_XI0/XI32/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM7 N_XI0/XI32/XI12/NET36_XI0/XI32/XI12/MM7_d
+ N_XI0/XI32/XI12/NET35_XI0/XI32/XI12/MM7_g N_VSS_XI0/XI32/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM8 N_XI0/XI32/XI12/NET35_XI0/XI32/XI12/MM8_d
+ N_WL<61>_XI0/XI32/XI12/MM8_g N_BLN<3>_XI0/XI32/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI12/MM5 N_XI0/XI32/XI12/NET34_XI0/XI32/XI12/MM5_d
+ N_XI0/XI32/XI12/NET33_XI0/XI32/XI12/MM5_g N_VDD_XI0/XI32/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI12/MM4 N_XI0/XI32/XI12/NET33_XI0/XI32/XI12/MM4_d
+ N_XI0/XI32/XI12/NET34_XI0/XI32/XI12/MM4_g N_VDD_XI0/XI32/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI12/MM10 N_XI0/XI32/XI12/NET35_XI0/XI32/XI12/MM10_d
+ N_XI0/XI32/XI12/NET36_XI0/XI32/XI12/MM10_g N_VDD_XI0/XI32/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI12/MM11 N_XI0/XI32/XI12/NET36_XI0/XI32/XI12/MM11_d
+ N_XI0/XI32/XI12/NET35_XI0/XI32/XI12/MM11_g N_VDD_XI0/XI32/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI13/MM2 N_XI0/XI32/XI13/NET34_XI0/XI32/XI13/MM2_d
+ N_XI0/XI32/XI13/NET33_XI0/XI32/XI13/MM2_g N_VSS_XI0/XI32/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM3 N_XI0/XI32/XI13/NET33_XI0/XI32/XI13/MM3_d
+ N_WL<60>_XI0/XI32/XI13/MM3_g N_BLN<2>_XI0/XI32/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM0 N_XI0/XI32/XI13/NET34_XI0/XI32/XI13/MM0_d
+ N_WL<60>_XI0/XI32/XI13/MM0_g N_BL<2>_XI0/XI32/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM1 N_XI0/XI32/XI13/NET33_XI0/XI32/XI13/MM1_d
+ N_XI0/XI32/XI13/NET34_XI0/XI32/XI13/MM1_g N_VSS_XI0/XI32/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM9 N_XI0/XI32/XI13/NET36_XI0/XI32/XI13/MM9_d
+ N_WL<61>_XI0/XI32/XI13/MM9_g N_BL<2>_XI0/XI32/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM6 N_XI0/XI32/XI13/NET35_XI0/XI32/XI13/MM6_d
+ N_XI0/XI32/XI13/NET36_XI0/XI32/XI13/MM6_g N_VSS_XI0/XI32/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM7 N_XI0/XI32/XI13/NET36_XI0/XI32/XI13/MM7_d
+ N_XI0/XI32/XI13/NET35_XI0/XI32/XI13/MM7_g N_VSS_XI0/XI32/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM8 N_XI0/XI32/XI13/NET35_XI0/XI32/XI13/MM8_d
+ N_WL<61>_XI0/XI32/XI13/MM8_g N_BLN<2>_XI0/XI32/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI13/MM5 N_XI0/XI32/XI13/NET34_XI0/XI32/XI13/MM5_d
+ N_XI0/XI32/XI13/NET33_XI0/XI32/XI13/MM5_g N_VDD_XI0/XI32/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI13/MM4 N_XI0/XI32/XI13/NET33_XI0/XI32/XI13/MM4_d
+ N_XI0/XI32/XI13/NET34_XI0/XI32/XI13/MM4_g N_VDD_XI0/XI32/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI13/MM10 N_XI0/XI32/XI13/NET35_XI0/XI32/XI13/MM10_d
+ N_XI0/XI32/XI13/NET36_XI0/XI32/XI13/MM10_g N_VDD_XI0/XI32/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI13/MM11 N_XI0/XI32/XI13/NET36_XI0/XI32/XI13/MM11_d
+ N_XI0/XI32/XI13/NET35_XI0/XI32/XI13/MM11_g N_VDD_XI0/XI32/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI14/MM2 N_XI0/XI32/XI14/NET34_XI0/XI32/XI14/MM2_d
+ N_XI0/XI32/XI14/NET33_XI0/XI32/XI14/MM2_g N_VSS_XI0/XI32/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM3 N_XI0/XI32/XI14/NET33_XI0/XI32/XI14/MM3_d
+ N_WL<60>_XI0/XI32/XI14/MM3_g N_BLN<1>_XI0/XI32/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM0 N_XI0/XI32/XI14/NET34_XI0/XI32/XI14/MM0_d
+ N_WL<60>_XI0/XI32/XI14/MM0_g N_BL<1>_XI0/XI32/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM1 N_XI0/XI32/XI14/NET33_XI0/XI32/XI14/MM1_d
+ N_XI0/XI32/XI14/NET34_XI0/XI32/XI14/MM1_g N_VSS_XI0/XI32/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM9 N_XI0/XI32/XI14/NET36_XI0/XI32/XI14/MM9_d
+ N_WL<61>_XI0/XI32/XI14/MM9_g N_BL<1>_XI0/XI32/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM6 N_XI0/XI32/XI14/NET35_XI0/XI32/XI14/MM6_d
+ N_XI0/XI32/XI14/NET36_XI0/XI32/XI14/MM6_g N_VSS_XI0/XI32/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM7 N_XI0/XI32/XI14/NET36_XI0/XI32/XI14/MM7_d
+ N_XI0/XI32/XI14/NET35_XI0/XI32/XI14/MM7_g N_VSS_XI0/XI32/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM8 N_XI0/XI32/XI14/NET35_XI0/XI32/XI14/MM8_d
+ N_WL<61>_XI0/XI32/XI14/MM8_g N_BLN<1>_XI0/XI32/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI14/MM5 N_XI0/XI32/XI14/NET34_XI0/XI32/XI14/MM5_d
+ N_XI0/XI32/XI14/NET33_XI0/XI32/XI14/MM5_g N_VDD_XI0/XI32/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI14/MM4 N_XI0/XI32/XI14/NET33_XI0/XI32/XI14/MM4_d
+ N_XI0/XI32/XI14/NET34_XI0/XI32/XI14/MM4_g N_VDD_XI0/XI32/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI14/MM10 N_XI0/XI32/XI14/NET35_XI0/XI32/XI14/MM10_d
+ N_XI0/XI32/XI14/NET36_XI0/XI32/XI14/MM10_g N_VDD_XI0/XI32/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI14/MM11 N_XI0/XI32/XI14/NET36_XI0/XI32/XI14/MM11_d
+ N_XI0/XI32/XI14/NET35_XI0/XI32/XI14/MM11_g N_VDD_XI0/XI32/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI15/MM2 N_XI0/XI32/XI15/NET34_XI0/XI32/XI15/MM2_d
+ N_XI0/XI32/XI15/NET33_XI0/XI32/XI15/MM2_g N_VSS_XI0/XI32/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM3 N_XI0/XI32/XI15/NET33_XI0/XI32/XI15/MM3_d
+ N_WL<60>_XI0/XI32/XI15/MM3_g N_BLN<0>_XI0/XI32/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM0 N_XI0/XI32/XI15/NET34_XI0/XI32/XI15/MM0_d
+ N_WL<60>_XI0/XI32/XI15/MM0_g N_BL<0>_XI0/XI32/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM1 N_XI0/XI32/XI15/NET33_XI0/XI32/XI15/MM1_d
+ N_XI0/XI32/XI15/NET34_XI0/XI32/XI15/MM1_g N_VSS_XI0/XI32/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM9 N_XI0/XI32/XI15/NET36_XI0/XI32/XI15/MM9_d
+ N_WL<61>_XI0/XI32/XI15/MM9_g N_BL<0>_XI0/XI32/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM6 N_XI0/XI32/XI15/NET35_XI0/XI32/XI15/MM6_d
+ N_XI0/XI32/XI15/NET36_XI0/XI32/XI15/MM6_g N_VSS_XI0/XI32/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM7 N_XI0/XI32/XI15/NET36_XI0/XI32/XI15/MM7_d
+ N_XI0/XI32/XI15/NET35_XI0/XI32/XI15/MM7_g N_VSS_XI0/XI32/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM8 N_XI0/XI32/XI15/NET35_XI0/XI32/XI15/MM8_d
+ N_WL<61>_XI0/XI32/XI15/MM8_g N_BLN<0>_XI0/XI32/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI32/XI15/MM5 N_XI0/XI32/XI15/NET34_XI0/XI32/XI15/MM5_d
+ N_XI0/XI32/XI15/NET33_XI0/XI32/XI15/MM5_g N_VDD_XI0/XI32/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI15/MM4 N_XI0/XI32/XI15/NET33_XI0/XI32/XI15/MM4_d
+ N_XI0/XI32/XI15/NET34_XI0/XI32/XI15/MM4_g N_VDD_XI0/XI32/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI15/MM10 N_XI0/XI32/XI15/NET35_XI0/XI32/XI15/MM10_d
+ N_XI0/XI32/XI15/NET36_XI0/XI32/XI15/MM10_g N_VDD_XI0/XI32/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI32/XI15/MM11 N_XI0/XI32/XI15/NET36_XI0/XI32/XI15/MM11_d
+ N_XI0/XI32/XI15/NET35_XI0/XI32/XI15/MM11_g N_VDD_XI0/XI32/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI0/MM2 N_XI0/XI33/XI0/NET34_XI0/XI33/XI0/MM2_d
+ N_XI0/XI33/XI0/NET33_XI0/XI33/XI0/MM2_g N_VSS_XI0/XI33/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM3 N_XI0/XI33/XI0/NET33_XI0/XI33/XI0/MM3_d
+ N_WL<62>_XI0/XI33/XI0/MM3_g N_BLN<15>_XI0/XI33/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM0 N_XI0/XI33/XI0/NET34_XI0/XI33/XI0/MM0_d
+ N_WL<62>_XI0/XI33/XI0/MM0_g N_BL<15>_XI0/XI33/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM1 N_XI0/XI33/XI0/NET33_XI0/XI33/XI0/MM1_d
+ N_XI0/XI33/XI0/NET34_XI0/XI33/XI0/MM1_g N_VSS_XI0/XI33/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM9 N_XI0/XI33/XI0/NET36_XI0/XI33/XI0/MM9_d
+ N_WL<63>_XI0/XI33/XI0/MM9_g N_BL<15>_XI0/XI33/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM6 N_XI0/XI33/XI0/NET35_XI0/XI33/XI0/MM6_d
+ N_XI0/XI33/XI0/NET36_XI0/XI33/XI0/MM6_g N_VSS_XI0/XI33/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM7 N_XI0/XI33/XI0/NET36_XI0/XI33/XI0/MM7_d
+ N_XI0/XI33/XI0/NET35_XI0/XI33/XI0/MM7_g N_VSS_XI0/XI33/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM8 N_XI0/XI33/XI0/NET35_XI0/XI33/XI0/MM8_d
+ N_WL<63>_XI0/XI33/XI0/MM8_g N_BLN<15>_XI0/XI33/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI0/MM5 N_XI0/XI33/XI0/NET34_XI0/XI33/XI0/MM5_d
+ N_XI0/XI33/XI0/NET33_XI0/XI33/XI0/MM5_g N_VDD_XI0/XI33/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI0/MM4 N_XI0/XI33/XI0/NET33_XI0/XI33/XI0/MM4_d
+ N_XI0/XI33/XI0/NET34_XI0/XI33/XI0/MM4_g N_VDD_XI0/XI33/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI0/MM10 N_XI0/XI33/XI0/NET35_XI0/XI33/XI0/MM10_d
+ N_XI0/XI33/XI0/NET36_XI0/XI33/XI0/MM10_g N_VDD_XI0/XI33/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI0/MM11 N_XI0/XI33/XI0/NET36_XI0/XI33/XI0/MM11_d
+ N_XI0/XI33/XI0/NET35_XI0/XI33/XI0/MM11_g N_VDD_XI0/XI33/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI1/MM2 N_XI0/XI33/XI1/NET34_XI0/XI33/XI1/MM2_d
+ N_XI0/XI33/XI1/NET33_XI0/XI33/XI1/MM2_g N_VSS_XI0/XI33/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM3 N_XI0/XI33/XI1/NET33_XI0/XI33/XI1/MM3_d
+ N_WL<62>_XI0/XI33/XI1/MM3_g N_BLN<14>_XI0/XI33/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM0 N_XI0/XI33/XI1/NET34_XI0/XI33/XI1/MM0_d
+ N_WL<62>_XI0/XI33/XI1/MM0_g N_BL<14>_XI0/XI33/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM1 N_XI0/XI33/XI1/NET33_XI0/XI33/XI1/MM1_d
+ N_XI0/XI33/XI1/NET34_XI0/XI33/XI1/MM1_g N_VSS_XI0/XI33/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM9 N_XI0/XI33/XI1/NET36_XI0/XI33/XI1/MM9_d
+ N_WL<63>_XI0/XI33/XI1/MM9_g N_BL<14>_XI0/XI33/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM6 N_XI0/XI33/XI1/NET35_XI0/XI33/XI1/MM6_d
+ N_XI0/XI33/XI1/NET36_XI0/XI33/XI1/MM6_g N_VSS_XI0/XI33/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM7 N_XI0/XI33/XI1/NET36_XI0/XI33/XI1/MM7_d
+ N_XI0/XI33/XI1/NET35_XI0/XI33/XI1/MM7_g N_VSS_XI0/XI33/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM8 N_XI0/XI33/XI1/NET35_XI0/XI33/XI1/MM8_d
+ N_WL<63>_XI0/XI33/XI1/MM8_g N_BLN<14>_XI0/XI33/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI1/MM5 N_XI0/XI33/XI1/NET34_XI0/XI33/XI1/MM5_d
+ N_XI0/XI33/XI1/NET33_XI0/XI33/XI1/MM5_g N_VDD_XI0/XI33/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI1/MM4 N_XI0/XI33/XI1/NET33_XI0/XI33/XI1/MM4_d
+ N_XI0/XI33/XI1/NET34_XI0/XI33/XI1/MM4_g N_VDD_XI0/XI33/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI1/MM10 N_XI0/XI33/XI1/NET35_XI0/XI33/XI1/MM10_d
+ N_XI0/XI33/XI1/NET36_XI0/XI33/XI1/MM10_g N_VDD_XI0/XI33/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI1/MM11 N_XI0/XI33/XI1/NET36_XI0/XI33/XI1/MM11_d
+ N_XI0/XI33/XI1/NET35_XI0/XI33/XI1/MM11_g N_VDD_XI0/XI33/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI2/MM2 N_XI0/XI33/XI2/NET34_XI0/XI33/XI2/MM2_d
+ N_XI0/XI33/XI2/NET33_XI0/XI33/XI2/MM2_g N_VSS_XI0/XI33/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM3 N_XI0/XI33/XI2/NET33_XI0/XI33/XI2/MM3_d
+ N_WL<62>_XI0/XI33/XI2/MM3_g N_BLN<13>_XI0/XI33/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM0 N_XI0/XI33/XI2/NET34_XI0/XI33/XI2/MM0_d
+ N_WL<62>_XI0/XI33/XI2/MM0_g N_BL<13>_XI0/XI33/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM1 N_XI0/XI33/XI2/NET33_XI0/XI33/XI2/MM1_d
+ N_XI0/XI33/XI2/NET34_XI0/XI33/XI2/MM1_g N_VSS_XI0/XI33/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM9 N_XI0/XI33/XI2/NET36_XI0/XI33/XI2/MM9_d
+ N_WL<63>_XI0/XI33/XI2/MM9_g N_BL<13>_XI0/XI33/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM6 N_XI0/XI33/XI2/NET35_XI0/XI33/XI2/MM6_d
+ N_XI0/XI33/XI2/NET36_XI0/XI33/XI2/MM6_g N_VSS_XI0/XI33/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM7 N_XI0/XI33/XI2/NET36_XI0/XI33/XI2/MM7_d
+ N_XI0/XI33/XI2/NET35_XI0/XI33/XI2/MM7_g N_VSS_XI0/XI33/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM8 N_XI0/XI33/XI2/NET35_XI0/XI33/XI2/MM8_d
+ N_WL<63>_XI0/XI33/XI2/MM8_g N_BLN<13>_XI0/XI33/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI2/MM5 N_XI0/XI33/XI2/NET34_XI0/XI33/XI2/MM5_d
+ N_XI0/XI33/XI2/NET33_XI0/XI33/XI2/MM5_g N_VDD_XI0/XI33/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI2/MM4 N_XI0/XI33/XI2/NET33_XI0/XI33/XI2/MM4_d
+ N_XI0/XI33/XI2/NET34_XI0/XI33/XI2/MM4_g N_VDD_XI0/XI33/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI2/MM10 N_XI0/XI33/XI2/NET35_XI0/XI33/XI2/MM10_d
+ N_XI0/XI33/XI2/NET36_XI0/XI33/XI2/MM10_g N_VDD_XI0/XI33/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI2/MM11 N_XI0/XI33/XI2/NET36_XI0/XI33/XI2/MM11_d
+ N_XI0/XI33/XI2/NET35_XI0/XI33/XI2/MM11_g N_VDD_XI0/XI33/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI3/MM2 N_XI0/XI33/XI3/NET34_XI0/XI33/XI3/MM2_d
+ N_XI0/XI33/XI3/NET33_XI0/XI33/XI3/MM2_g N_VSS_XI0/XI33/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM3 N_XI0/XI33/XI3/NET33_XI0/XI33/XI3/MM3_d
+ N_WL<62>_XI0/XI33/XI3/MM3_g N_BLN<12>_XI0/XI33/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM0 N_XI0/XI33/XI3/NET34_XI0/XI33/XI3/MM0_d
+ N_WL<62>_XI0/XI33/XI3/MM0_g N_BL<12>_XI0/XI33/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM1 N_XI0/XI33/XI3/NET33_XI0/XI33/XI3/MM1_d
+ N_XI0/XI33/XI3/NET34_XI0/XI33/XI3/MM1_g N_VSS_XI0/XI33/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM9 N_XI0/XI33/XI3/NET36_XI0/XI33/XI3/MM9_d
+ N_WL<63>_XI0/XI33/XI3/MM9_g N_BL<12>_XI0/XI33/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM6 N_XI0/XI33/XI3/NET35_XI0/XI33/XI3/MM6_d
+ N_XI0/XI33/XI3/NET36_XI0/XI33/XI3/MM6_g N_VSS_XI0/XI33/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM7 N_XI0/XI33/XI3/NET36_XI0/XI33/XI3/MM7_d
+ N_XI0/XI33/XI3/NET35_XI0/XI33/XI3/MM7_g N_VSS_XI0/XI33/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM8 N_XI0/XI33/XI3/NET35_XI0/XI33/XI3/MM8_d
+ N_WL<63>_XI0/XI33/XI3/MM8_g N_BLN<12>_XI0/XI33/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI3/MM5 N_XI0/XI33/XI3/NET34_XI0/XI33/XI3/MM5_d
+ N_XI0/XI33/XI3/NET33_XI0/XI33/XI3/MM5_g N_VDD_XI0/XI33/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI3/MM4 N_XI0/XI33/XI3/NET33_XI0/XI33/XI3/MM4_d
+ N_XI0/XI33/XI3/NET34_XI0/XI33/XI3/MM4_g N_VDD_XI0/XI33/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI3/MM10 N_XI0/XI33/XI3/NET35_XI0/XI33/XI3/MM10_d
+ N_XI0/XI33/XI3/NET36_XI0/XI33/XI3/MM10_g N_VDD_XI0/XI33/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI3/MM11 N_XI0/XI33/XI3/NET36_XI0/XI33/XI3/MM11_d
+ N_XI0/XI33/XI3/NET35_XI0/XI33/XI3/MM11_g N_VDD_XI0/XI33/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI4/MM2 N_XI0/XI33/XI4/NET34_XI0/XI33/XI4/MM2_d
+ N_XI0/XI33/XI4/NET33_XI0/XI33/XI4/MM2_g N_VSS_XI0/XI33/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM3 N_XI0/XI33/XI4/NET33_XI0/XI33/XI4/MM3_d
+ N_WL<62>_XI0/XI33/XI4/MM3_g N_BLN<11>_XI0/XI33/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM0 N_XI0/XI33/XI4/NET34_XI0/XI33/XI4/MM0_d
+ N_WL<62>_XI0/XI33/XI4/MM0_g N_BL<11>_XI0/XI33/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM1 N_XI0/XI33/XI4/NET33_XI0/XI33/XI4/MM1_d
+ N_XI0/XI33/XI4/NET34_XI0/XI33/XI4/MM1_g N_VSS_XI0/XI33/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM9 N_XI0/XI33/XI4/NET36_XI0/XI33/XI4/MM9_d
+ N_WL<63>_XI0/XI33/XI4/MM9_g N_BL<11>_XI0/XI33/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM6 N_XI0/XI33/XI4/NET35_XI0/XI33/XI4/MM6_d
+ N_XI0/XI33/XI4/NET36_XI0/XI33/XI4/MM6_g N_VSS_XI0/XI33/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM7 N_XI0/XI33/XI4/NET36_XI0/XI33/XI4/MM7_d
+ N_XI0/XI33/XI4/NET35_XI0/XI33/XI4/MM7_g N_VSS_XI0/XI33/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM8 N_XI0/XI33/XI4/NET35_XI0/XI33/XI4/MM8_d
+ N_WL<63>_XI0/XI33/XI4/MM8_g N_BLN<11>_XI0/XI33/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI4/MM5 N_XI0/XI33/XI4/NET34_XI0/XI33/XI4/MM5_d
+ N_XI0/XI33/XI4/NET33_XI0/XI33/XI4/MM5_g N_VDD_XI0/XI33/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI4/MM4 N_XI0/XI33/XI4/NET33_XI0/XI33/XI4/MM4_d
+ N_XI0/XI33/XI4/NET34_XI0/XI33/XI4/MM4_g N_VDD_XI0/XI33/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI4/MM10 N_XI0/XI33/XI4/NET35_XI0/XI33/XI4/MM10_d
+ N_XI0/XI33/XI4/NET36_XI0/XI33/XI4/MM10_g N_VDD_XI0/XI33/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI4/MM11 N_XI0/XI33/XI4/NET36_XI0/XI33/XI4/MM11_d
+ N_XI0/XI33/XI4/NET35_XI0/XI33/XI4/MM11_g N_VDD_XI0/XI33/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI5/MM2 N_XI0/XI33/XI5/NET34_XI0/XI33/XI5/MM2_d
+ N_XI0/XI33/XI5/NET33_XI0/XI33/XI5/MM2_g N_VSS_XI0/XI33/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM3 N_XI0/XI33/XI5/NET33_XI0/XI33/XI5/MM3_d
+ N_WL<62>_XI0/XI33/XI5/MM3_g N_BLN<10>_XI0/XI33/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM0 N_XI0/XI33/XI5/NET34_XI0/XI33/XI5/MM0_d
+ N_WL<62>_XI0/XI33/XI5/MM0_g N_BL<10>_XI0/XI33/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM1 N_XI0/XI33/XI5/NET33_XI0/XI33/XI5/MM1_d
+ N_XI0/XI33/XI5/NET34_XI0/XI33/XI5/MM1_g N_VSS_XI0/XI33/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM9 N_XI0/XI33/XI5/NET36_XI0/XI33/XI5/MM9_d
+ N_WL<63>_XI0/XI33/XI5/MM9_g N_BL<10>_XI0/XI33/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM6 N_XI0/XI33/XI5/NET35_XI0/XI33/XI5/MM6_d
+ N_XI0/XI33/XI5/NET36_XI0/XI33/XI5/MM6_g N_VSS_XI0/XI33/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM7 N_XI0/XI33/XI5/NET36_XI0/XI33/XI5/MM7_d
+ N_XI0/XI33/XI5/NET35_XI0/XI33/XI5/MM7_g N_VSS_XI0/XI33/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM8 N_XI0/XI33/XI5/NET35_XI0/XI33/XI5/MM8_d
+ N_WL<63>_XI0/XI33/XI5/MM8_g N_BLN<10>_XI0/XI33/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI5/MM5 N_XI0/XI33/XI5/NET34_XI0/XI33/XI5/MM5_d
+ N_XI0/XI33/XI5/NET33_XI0/XI33/XI5/MM5_g N_VDD_XI0/XI33/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI5/MM4 N_XI0/XI33/XI5/NET33_XI0/XI33/XI5/MM4_d
+ N_XI0/XI33/XI5/NET34_XI0/XI33/XI5/MM4_g N_VDD_XI0/XI33/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI5/MM10 N_XI0/XI33/XI5/NET35_XI0/XI33/XI5/MM10_d
+ N_XI0/XI33/XI5/NET36_XI0/XI33/XI5/MM10_g N_VDD_XI0/XI33/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI5/MM11 N_XI0/XI33/XI5/NET36_XI0/XI33/XI5/MM11_d
+ N_XI0/XI33/XI5/NET35_XI0/XI33/XI5/MM11_g N_VDD_XI0/XI33/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI6/MM2 N_XI0/XI33/XI6/NET34_XI0/XI33/XI6/MM2_d
+ N_XI0/XI33/XI6/NET33_XI0/XI33/XI6/MM2_g N_VSS_XI0/XI33/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM3 N_XI0/XI33/XI6/NET33_XI0/XI33/XI6/MM3_d
+ N_WL<62>_XI0/XI33/XI6/MM3_g N_BLN<9>_XI0/XI33/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM0 N_XI0/XI33/XI6/NET34_XI0/XI33/XI6/MM0_d
+ N_WL<62>_XI0/XI33/XI6/MM0_g N_BL<9>_XI0/XI33/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM1 N_XI0/XI33/XI6/NET33_XI0/XI33/XI6/MM1_d
+ N_XI0/XI33/XI6/NET34_XI0/XI33/XI6/MM1_g N_VSS_XI0/XI33/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM9 N_XI0/XI33/XI6/NET36_XI0/XI33/XI6/MM9_d
+ N_WL<63>_XI0/XI33/XI6/MM9_g N_BL<9>_XI0/XI33/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM6 N_XI0/XI33/XI6/NET35_XI0/XI33/XI6/MM6_d
+ N_XI0/XI33/XI6/NET36_XI0/XI33/XI6/MM6_g N_VSS_XI0/XI33/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM7 N_XI0/XI33/XI6/NET36_XI0/XI33/XI6/MM7_d
+ N_XI0/XI33/XI6/NET35_XI0/XI33/XI6/MM7_g N_VSS_XI0/XI33/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM8 N_XI0/XI33/XI6/NET35_XI0/XI33/XI6/MM8_d
+ N_WL<63>_XI0/XI33/XI6/MM8_g N_BLN<9>_XI0/XI33/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI6/MM5 N_XI0/XI33/XI6/NET34_XI0/XI33/XI6/MM5_d
+ N_XI0/XI33/XI6/NET33_XI0/XI33/XI6/MM5_g N_VDD_XI0/XI33/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI6/MM4 N_XI0/XI33/XI6/NET33_XI0/XI33/XI6/MM4_d
+ N_XI0/XI33/XI6/NET34_XI0/XI33/XI6/MM4_g N_VDD_XI0/XI33/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI6/MM10 N_XI0/XI33/XI6/NET35_XI0/XI33/XI6/MM10_d
+ N_XI0/XI33/XI6/NET36_XI0/XI33/XI6/MM10_g N_VDD_XI0/XI33/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI6/MM11 N_XI0/XI33/XI6/NET36_XI0/XI33/XI6/MM11_d
+ N_XI0/XI33/XI6/NET35_XI0/XI33/XI6/MM11_g N_VDD_XI0/XI33/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI7/MM2 N_XI0/XI33/XI7/NET34_XI0/XI33/XI7/MM2_d
+ N_XI0/XI33/XI7/NET33_XI0/XI33/XI7/MM2_g N_VSS_XI0/XI33/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM3 N_XI0/XI33/XI7/NET33_XI0/XI33/XI7/MM3_d
+ N_WL<62>_XI0/XI33/XI7/MM3_g N_BLN<8>_XI0/XI33/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM0 N_XI0/XI33/XI7/NET34_XI0/XI33/XI7/MM0_d
+ N_WL<62>_XI0/XI33/XI7/MM0_g N_BL<8>_XI0/XI33/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM1 N_XI0/XI33/XI7/NET33_XI0/XI33/XI7/MM1_d
+ N_XI0/XI33/XI7/NET34_XI0/XI33/XI7/MM1_g N_VSS_XI0/XI33/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM9 N_XI0/XI33/XI7/NET36_XI0/XI33/XI7/MM9_d
+ N_WL<63>_XI0/XI33/XI7/MM9_g N_BL<8>_XI0/XI33/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM6 N_XI0/XI33/XI7/NET35_XI0/XI33/XI7/MM6_d
+ N_XI0/XI33/XI7/NET36_XI0/XI33/XI7/MM6_g N_VSS_XI0/XI33/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM7 N_XI0/XI33/XI7/NET36_XI0/XI33/XI7/MM7_d
+ N_XI0/XI33/XI7/NET35_XI0/XI33/XI7/MM7_g N_VSS_XI0/XI33/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM8 N_XI0/XI33/XI7/NET35_XI0/XI33/XI7/MM8_d
+ N_WL<63>_XI0/XI33/XI7/MM8_g N_BLN<8>_XI0/XI33/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI7/MM5 N_XI0/XI33/XI7/NET34_XI0/XI33/XI7/MM5_d
+ N_XI0/XI33/XI7/NET33_XI0/XI33/XI7/MM5_g N_VDD_XI0/XI33/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI7/MM4 N_XI0/XI33/XI7/NET33_XI0/XI33/XI7/MM4_d
+ N_XI0/XI33/XI7/NET34_XI0/XI33/XI7/MM4_g N_VDD_XI0/XI33/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI7/MM10 N_XI0/XI33/XI7/NET35_XI0/XI33/XI7/MM10_d
+ N_XI0/XI33/XI7/NET36_XI0/XI33/XI7/MM10_g N_VDD_XI0/XI33/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI7/MM11 N_XI0/XI33/XI7/NET36_XI0/XI33/XI7/MM11_d
+ N_XI0/XI33/XI7/NET35_XI0/XI33/XI7/MM11_g N_VDD_XI0/XI33/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI8/MM2 N_XI0/XI33/XI8/NET34_XI0/XI33/XI8/MM2_d
+ N_XI0/XI33/XI8/NET33_XI0/XI33/XI8/MM2_g N_VSS_XI0/XI33/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM3 N_XI0/XI33/XI8/NET33_XI0/XI33/XI8/MM3_d
+ N_WL<62>_XI0/XI33/XI8/MM3_g N_BLN<7>_XI0/XI33/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM0 N_XI0/XI33/XI8/NET34_XI0/XI33/XI8/MM0_d
+ N_WL<62>_XI0/XI33/XI8/MM0_g N_BL<7>_XI0/XI33/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM1 N_XI0/XI33/XI8/NET33_XI0/XI33/XI8/MM1_d
+ N_XI0/XI33/XI8/NET34_XI0/XI33/XI8/MM1_g N_VSS_XI0/XI33/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM9 N_XI0/XI33/XI8/NET36_XI0/XI33/XI8/MM9_d
+ N_WL<63>_XI0/XI33/XI8/MM9_g N_BL<7>_XI0/XI33/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM6 N_XI0/XI33/XI8/NET35_XI0/XI33/XI8/MM6_d
+ N_XI0/XI33/XI8/NET36_XI0/XI33/XI8/MM6_g N_VSS_XI0/XI33/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM7 N_XI0/XI33/XI8/NET36_XI0/XI33/XI8/MM7_d
+ N_XI0/XI33/XI8/NET35_XI0/XI33/XI8/MM7_g N_VSS_XI0/XI33/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM8 N_XI0/XI33/XI8/NET35_XI0/XI33/XI8/MM8_d
+ N_WL<63>_XI0/XI33/XI8/MM8_g N_BLN<7>_XI0/XI33/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI8/MM5 N_XI0/XI33/XI8/NET34_XI0/XI33/XI8/MM5_d
+ N_XI0/XI33/XI8/NET33_XI0/XI33/XI8/MM5_g N_VDD_XI0/XI33/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI8/MM4 N_XI0/XI33/XI8/NET33_XI0/XI33/XI8/MM4_d
+ N_XI0/XI33/XI8/NET34_XI0/XI33/XI8/MM4_g N_VDD_XI0/XI33/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI8/MM10 N_XI0/XI33/XI8/NET35_XI0/XI33/XI8/MM10_d
+ N_XI0/XI33/XI8/NET36_XI0/XI33/XI8/MM10_g N_VDD_XI0/XI33/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI8/MM11 N_XI0/XI33/XI8/NET36_XI0/XI33/XI8/MM11_d
+ N_XI0/XI33/XI8/NET35_XI0/XI33/XI8/MM11_g N_VDD_XI0/XI33/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI9/MM2 N_XI0/XI33/XI9/NET34_XI0/XI33/XI9/MM2_d
+ N_XI0/XI33/XI9/NET33_XI0/XI33/XI9/MM2_g N_VSS_XI0/XI33/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM3 N_XI0/XI33/XI9/NET33_XI0/XI33/XI9/MM3_d
+ N_WL<62>_XI0/XI33/XI9/MM3_g N_BLN<6>_XI0/XI33/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM0 N_XI0/XI33/XI9/NET34_XI0/XI33/XI9/MM0_d
+ N_WL<62>_XI0/XI33/XI9/MM0_g N_BL<6>_XI0/XI33/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM1 N_XI0/XI33/XI9/NET33_XI0/XI33/XI9/MM1_d
+ N_XI0/XI33/XI9/NET34_XI0/XI33/XI9/MM1_g N_VSS_XI0/XI33/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM9 N_XI0/XI33/XI9/NET36_XI0/XI33/XI9/MM9_d
+ N_WL<63>_XI0/XI33/XI9/MM9_g N_BL<6>_XI0/XI33/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM6 N_XI0/XI33/XI9/NET35_XI0/XI33/XI9/MM6_d
+ N_XI0/XI33/XI9/NET36_XI0/XI33/XI9/MM6_g N_VSS_XI0/XI33/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM7 N_XI0/XI33/XI9/NET36_XI0/XI33/XI9/MM7_d
+ N_XI0/XI33/XI9/NET35_XI0/XI33/XI9/MM7_g N_VSS_XI0/XI33/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM8 N_XI0/XI33/XI9/NET35_XI0/XI33/XI9/MM8_d
+ N_WL<63>_XI0/XI33/XI9/MM8_g N_BLN<6>_XI0/XI33/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI9/MM5 N_XI0/XI33/XI9/NET34_XI0/XI33/XI9/MM5_d
+ N_XI0/XI33/XI9/NET33_XI0/XI33/XI9/MM5_g N_VDD_XI0/XI33/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI9/MM4 N_XI0/XI33/XI9/NET33_XI0/XI33/XI9/MM4_d
+ N_XI0/XI33/XI9/NET34_XI0/XI33/XI9/MM4_g N_VDD_XI0/XI33/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI9/MM10 N_XI0/XI33/XI9/NET35_XI0/XI33/XI9/MM10_d
+ N_XI0/XI33/XI9/NET36_XI0/XI33/XI9/MM10_g N_VDD_XI0/XI33/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI9/MM11 N_XI0/XI33/XI9/NET36_XI0/XI33/XI9/MM11_d
+ N_XI0/XI33/XI9/NET35_XI0/XI33/XI9/MM11_g N_VDD_XI0/XI33/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI10/MM2 N_XI0/XI33/XI10/NET34_XI0/XI33/XI10/MM2_d
+ N_XI0/XI33/XI10/NET33_XI0/XI33/XI10/MM2_g N_VSS_XI0/XI33/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM3 N_XI0/XI33/XI10/NET33_XI0/XI33/XI10/MM3_d
+ N_WL<62>_XI0/XI33/XI10/MM3_g N_BLN<5>_XI0/XI33/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM0 N_XI0/XI33/XI10/NET34_XI0/XI33/XI10/MM0_d
+ N_WL<62>_XI0/XI33/XI10/MM0_g N_BL<5>_XI0/XI33/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM1 N_XI0/XI33/XI10/NET33_XI0/XI33/XI10/MM1_d
+ N_XI0/XI33/XI10/NET34_XI0/XI33/XI10/MM1_g N_VSS_XI0/XI33/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM9 N_XI0/XI33/XI10/NET36_XI0/XI33/XI10/MM9_d
+ N_WL<63>_XI0/XI33/XI10/MM9_g N_BL<5>_XI0/XI33/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM6 N_XI0/XI33/XI10/NET35_XI0/XI33/XI10/MM6_d
+ N_XI0/XI33/XI10/NET36_XI0/XI33/XI10/MM6_g N_VSS_XI0/XI33/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM7 N_XI0/XI33/XI10/NET36_XI0/XI33/XI10/MM7_d
+ N_XI0/XI33/XI10/NET35_XI0/XI33/XI10/MM7_g N_VSS_XI0/XI33/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM8 N_XI0/XI33/XI10/NET35_XI0/XI33/XI10/MM8_d
+ N_WL<63>_XI0/XI33/XI10/MM8_g N_BLN<5>_XI0/XI33/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI10/MM5 N_XI0/XI33/XI10/NET34_XI0/XI33/XI10/MM5_d
+ N_XI0/XI33/XI10/NET33_XI0/XI33/XI10/MM5_g N_VDD_XI0/XI33/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI10/MM4 N_XI0/XI33/XI10/NET33_XI0/XI33/XI10/MM4_d
+ N_XI0/XI33/XI10/NET34_XI0/XI33/XI10/MM4_g N_VDD_XI0/XI33/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI10/MM10 N_XI0/XI33/XI10/NET35_XI0/XI33/XI10/MM10_d
+ N_XI0/XI33/XI10/NET36_XI0/XI33/XI10/MM10_g N_VDD_XI0/XI33/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI10/MM11 N_XI0/XI33/XI10/NET36_XI0/XI33/XI10/MM11_d
+ N_XI0/XI33/XI10/NET35_XI0/XI33/XI10/MM11_g N_VDD_XI0/XI33/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI11/MM2 N_XI0/XI33/XI11/NET34_XI0/XI33/XI11/MM2_d
+ N_XI0/XI33/XI11/NET33_XI0/XI33/XI11/MM2_g N_VSS_XI0/XI33/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM3 N_XI0/XI33/XI11/NET33_XI0/XI33/XI11/MM3_d
+ N_WL<62>_XI0/XI33/XI11/MM3_g N_BLN<4>_XI0/XI33/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM0 N_XI0/XI33/XI11/NET34_XI0/XI33/XI11/MM0_d
+ N_WL<62>_XI0/XI33/XI11/MM0_g N_BL<4>_XI0/XI33/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM1 N_XI0/XI33/XI11/NET33_XI0/XI33/XI11/MM1_d
+ N_XI0/XI33/XI11/NET34_XI0/XI33/XI11/MM1_g N_VSS_XI0/XI33/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM9 N_XI0/XI33/XI11/NET36_XI0/XI33/XI11/MM9_d
+ N_WL<63>_XI0/XI33/XI11/MM9_g N_BL<4>_XI0/XI33/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM6 N_XI0/XI33/XI11/NET35_XI0/XI33/XI11/MM6_d
+ N_XI0/XI33/XI11/NET36_XI0/XI33/XI11/MM6_g N_VSS_XI0/XI33/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM7 N_XI0/XI33/XI11/NET36_XI0/XI33/XI11/MM7_d
+ N_XI0/XI33/XI11/NET35_XI0/XI33/XI11/MM7_g N_VSS_XI0/XI33/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM8 N_XI0/XI33/XI11/NET35_XI0/XI33/XI11/MM8_d
+ N_WL<63>_XI0/XI33/XI11/MM8_g N_BLN<4>_XI0/XI33/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI11/MM5 N_XI0/XI33/XI11/NET34_XI0/XI33/XI11/MM5_d
+ N_XI0/XI33/XI11/NET33_XI0/XI33/XI11/MM5_g N_VDD_XI0/XI33/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI11/MM4 N_XI0/XI33/XI11/NET33_XI0/XI33/XI11/MM4_d
+ N_XI0/XI33/XI11/NET34_XI0/XI33/XI11/MM4_g N_VDD_XI0/XI33/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI11/MM10 N_XI0/XI33/XI11/NET35_XI0/XI33/XI11/MM10_d
+ N_XI0/XI33/XI11/NET36_XI0/XI33/XI11/MM10_g N_VDD_XI0/XI33/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI11/MM11 N_XI0/XI33/XI11/NET36_XI0/XI33/XI11/MM11_d
+ N_XI0/XI33/XI11/NET35_XI0/XI33/XI11/MM11_g N_VDD_XI0/XI33/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI12/MM2 N_XI0/XI33/XI12/NET34_XI0/XI33/XI12/MM2_d
+ N_XI0/XI33/XI12/NET33_XI0/XI33/XI12/MM2_g N_VSS_XI0/XI33/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM3 N_XI0/XI33/XI12/NET33_XI0/XI33/XI12/MM3_d
+ N_WL<62>_XI0/XI33/XI12/MM3_g N_BLN<3>_XI0/XI33/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM0 N_XI0/XI33/XI12/NET34_XI0/XI33/XI12/MM0_d
+ N_WL<62>_XI0/XI33/XI12/MM0_g N_BL<3>_XI0/XI33/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM1 N_XI0/XI33/XI12/NET33_XI0/XI33/XI12/MM1_d
+ N_XI0/XI33/XI12/NET34_XI0/XI33/XI12/MM1_g N_VSS_XI0/XI33/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM9 N_XI0/XI33/XI12/NET36_XI0/XI33/XI12/MM9_d
+ N_WL<63>_XI0/XI33/XI12/MM9_g N_BL<3>_XI0/XI33/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM6 N_XI0/XI33/XI12/NET35_XI0/XI33/XI12/MM6_d
+ N_XI0/XI33/XI12/NET36_XI0/XI33/XI12/MM6_g N_VSS_XI0/XI33/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM7 N_XI0/XI33/XI12/NET36_XI0/XI33/XI12/MM7_d
+ N_XI0/XI33/XI12/NET35_XI0/XI33/XI12/MM7_g N_VSS_XI0/XI33/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM8 N_XI0/XI33/XI12/NET35_XI0/XI33/XI12/MM8_d
+ N_WL<63>_XI0/XI33/XI12/MM8_g N_BLN<3>_XI0/XI33/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI12/MM5 N_XI0/XI33/XI12/NET34_XI0/XI33/XI12/MM5_d
+ N_XI0/XI33/XI12/NET33_XI0/XI33/XI12/MM5_g N_VDD_XI0/XI33/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI12/MM4 N_XI0/XI33/XI12/NET33_XI0/XI33/XI12/MM4_d
+ N_XI0/XI33/XI12/NET34_XI0/XI33/XI12/MM4_g N_VDD_XI0/XI33/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI12/MM10 N_XI0/XI33/XI12/NET35_XI0/XI33/XI12/MM10_d
+ N_XI0/XI33/XI12/NET36_XI0/XI33/XI12/MM10_g N_VDD_XI0/XI33/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI12/MM11 N_XI0/XI33/XI12/NET36_XI0/XI33/XI12/MM11_d
+ N_XI0/XI33/XI12/NET35_XI0/XI33/XI12/MM11_g N_VDD_XI0/XI33/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI13/MM2 N_XI0/XI33/XI13/NET34_XI0/XI33/XI13/MM2_d
+ N_XI0/XI33/XI13/NET33_XI0/XI33/XI13/MM2_g N_VSS_XI0/XI33/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM3 N_XI0/XI33/XI13/NET33_XI0/XI33/XI13/MM3_d
+ N_WL<62>_XI0/XI33/XI13/MM3_g N_BLN<2>_XI0/XI33/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM0 N_XI0/XI33/XI13/NET34_XI0/XI33/XI13/MM0_d
+ N_WL<62>_XI0/XI33/XI13/MM0_g N_BL<2>_XI0/XI33/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM1 N_XI0/XI33/XI13/NET33_XI0/XI33/XI13/MM1_d
+ N_XI0/XI33/XI13/NET34_XI0/XI33/XI13/MM1_g N_VSS_XI0/XI33/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM9 N_XI0/XI33/XI13/NET36_XI0/XI33/XI13/MM9_d
+ N_WL<63>_XI0/XI33/XI13/MM9_g N_BL<2>_XI0/XI33/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM6 N_XI0/XI33/XI13/NET35_XI0/XI33/XI13/MM6_d
+ N_XI0/XI33/XI13/NET36_XI0/XI33/XI13/MM6_g N_VSS_XI0/XI33/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM7 N_XI0/XI33/XI13/NET36_XI0/XI33/XI13/MM7_d
+ N_XI0/XI33/XI13/NET35_XI0/XI33/XI13/MM7_g N_VSS_XI0/XI33/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM8 N_XI0/XI33/XI13/NET35_XI0/XI33/XI13/MM8_d
+ N_WL<63>_XI0/XI33/XI13/MM8_g N_BLN<2>_XI0/XI33/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI13/MM5 N_XI0/XI33/XI13/NET34_XI0/XI33/XI13/MM5_d
+ N_XI0/XI33/XI13/NET33_XI0/XI33/XI13/MM5_g N_VDD_XI0/XI33/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI13/MM4 N_XI0/XI33/XI13/NET33_XI0/XI33/XI13/MM4_d
+ N_XI0/XI33/XI13/NET34_XI0/XI33/XI13/MM4_g N_VDD_XI0/XI33/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI13/MM10 N_XI0/XI33/XI13/NET35_XI0/XI33/XI13/MM10_d
+ N_XI0/XI33/XI13/NET36_XI0/XI33/XI13/MM10_g N_VDD_XI0/XI33/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI13/MM11 N_XI0/XI33/XI13/NET36_XI0/XI33/XI13/MM11_d
+ N_XI0/XI33/XI13/NET35_XI0/XI33/XI13/MM11_g N_VDD_XI0/XI33/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI14/MM2 N_XI0/XI33/XI14/NET34_XI0/XI33/XI14/MM2_d
+ N_XI0/XI33/XI14/NET33_XI0/XI33/XI14/MM2_g N_VSS_XI0/XI33/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM3 N_XI0/XI33/XI14/NET33_XI0/XI33/XI14/MM3_d
+ N_WL<62>_XI0/XI33/XI14/MM3_g N_BLN<1>_XI0/XI33/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM0 N_XI0/XI33/XI14/NET34_XI0/XI33/XI14/MM0_d
+ N_WL<62>_XI0/XI33/XI14/MM0_g N_BL<1>_XI0/XI33/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM1 N_XI0/XI33/XI14/NET33_XI0/XI33/XI14/MM1_d
+ N_XI0/XI33/XI14/NET34_XI0/XI33/XI14/MM1_g N_VSS_XI0/XI33/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM9 N_XI0/XI33/XI14/NET36_XI0/XI33/XI14/MM9_d
+ N_WL<63>_XI0/XI33/XI14/MM9_g N_BL<1>_XI0/XI33/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM6 N_XI0/XI33/XI14/NET35_XI0/XI33/XI14/MM6_d
+ N_XI0/XI33/XI14/NET36_XI0/XI33/XI14/MM6_g N_VSS_XI0/XI33/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM7 N_XI0/XI33/XI14/NET36_XI0/XI33/XI14/MM7_d
+ N_XI0/XI33/XI14/NET35_XI0/XI33/XI14/MM7_g N_VSS_XI0/XI33/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM8 N_XI0/XI33/XI14/NET35_XI0/XI33/XI14/MM8_d
+ N_WL<63>_XI0/XI33/XI14/MM8_g N_BLN<1>_XI0/XI33/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI14/MM5 N_XI0/XI33/XI14/NET34_XI0/XI33/XI14/MM5_d
+ N_XI0/XI33/XI14/NET33_XI0/XI33/XI14/MM5_g N_VDD_XI0/XI33/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI14/MM4 N_XI0/XI33/XI14/NET33_XI0/XI33/XI14/MM4_d
+ N_XI0/XI33/XI14/NET34_XI0/XI33/XI14/MM4_g N_VDD_XI0/XI33/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI14/MM10 N_XI0/XI33/XI14/NET35_XI0/XI33/XI14/MM10_d
+ N_XI0/XI33/XI14/NET36_XI0/XI33/XI14/MM10_g N_VDD_XI0/XI33/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI14/MM11 N_XI0/XI33/XI14/NET36_XI0/XI33/XI14/MM11_d
+ N_XI0/XI33/XI14/NET35_XI0/XI33/XI14/MM11_g N_VDD_XI0/XI33/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI15/MM2 N_XI0/XI33/XI15/NET34_XI0/XI33/XI15/MM2_d
+ N_XI0/XI33/XI15/NET33_XI0/XI33/XI15/MM2_g N_VSS_XI0/XI33/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM3 N_XI0/XI33/XI15/NET33_XI0/XI33/XI15/MM3_d
+ N_WL<62>_XI0/XI33/XI15/MM3_g N_BLN<0>_XI0/XI33/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM0 N_XI0/XI33/XI15/NET34_XI0/XI33/XI15/MM0_d
+ N_WL<62>_XI0/XI33/XI15/MM0_g N_BL<0>_XI0/XI33/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM1 N_XI0/XI33/XI15/NET33_XI0/XI33/XI15/MM1_d
+ N_XI0/XI33/XI15/NET34_XI0/XI33/XI15/MM1_g N_VSS_XI0/XI33/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM9 N_XI0/XI33/XI15/NET36_XI0/XI33/XI15/MM9_d
+ N_WL<63>_XI0/XI33/XI15/MM9_g N_BL<0>_XI0/XI33/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM6 N_XI0/XI33/XI15/NET35_XI0/XI33/XI15/MM6_d
+ N_XI0/XI33/XI15/NET36_XI0/XI33/XI15/MM6_g N_VSS_XI0/XI33/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM7 N_XI0/XI33/XI15/NET36_XI0/XI33/XI15/MM7_d
+ N_XI0/XI33/XI15/NET35_XI0/XI33/XI15/MM7_g N_VSS_XI0/XI33/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM8 N_XI0/XI33/XI15/NET35_XI0/XI33/XI15/MM8_d
+ N_WL<63>_XI0/XI33/XI15/MM8_g N_BLN<0>_XI0/XI33/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI33/XI15/MM5 N_XI0/XI33/XI15/NET34_XI0/XI33/XI15/MM5_d
+ N_XI0/XI33/XI15/NET33_XI0/XI33/XI15/MM5_g N_VDD_XI0/XI33/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI15/MM4 N_XI0/XI33/XI15/NET33_XI0/XI33/XI15/MM4_d
+ N_XI0/XI33/XI15/NET34_XI0/XI33/XI15/MM4_g N_VDD_XI0/XI33/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI15/MM10 N_XI0/XI33/XI15/NET35_XI0/XI33/XI15/MM10_d
+ N_XI0/XI33/XI15/NET36_XI0/XI33/XI15/MM10_g N_VDD_XI0/XI33/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI33/XI15/MM11 N_XI0/XI33/XI15/NET36_XI0/XI33/XI15/MM11_d
+ N_XI0/XI33/XI15/NET35_XI0/XI33/XI15/MM11_g N_VDD_XI0/XI33/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI0/MM2 N_XI0/XI34/XI0/NET34_XI0/XI34/XI0/MM2_d
+ N_XI0/XI34/XI0/NET33_XI0/XI34/XI0/MM2_g N_VSS_XI0/XI34/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM3 N_XI0/XI34/XI0/NET33_XI0/XI34/XI0/MM3_d
+ N_WL<64>_XI0/XI34/XI0/MM3_g N_BLN<15>_XI0/XI34/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM0 N_XI0/XI34/XI0/NET34_XI0/XI34/XI0/MM0_d
+ N_WL<64>_XI0/XI34/XI0/MM0_g N_BL<15>_XI0/XI34/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM1 N_XI0/XI34/XI0/NET33_XI0/XI34/XI0/MM1_d
+ N_XI0/XI34/XI0/NET34_XI0/XI34/XI0/MM1_g N_VSS_XI0/XI34/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM9 N_XI0/XI34/XI0/NET36_XI0/XI34/XI0/MM9_d
+ N_WL<65>_XI0/XI34/XI0/MM9_g N_BL<15>_XI0/XI34/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM6 N_XI0/XI34/XI0/NET35_XI0/XI34/XI0/MM6_d
+ N_XI0/XI34/XI0/NET36_XI0/XI34/XI0/MM6_g N_VSS_XI0/XI34/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM7 N_XI0/XI34/XI0/NET36_XI0/XI34/XI0/MM7_d
+ N_XI0/XI34/XI0/NET35_XI0/XI34/XI0/MM7_g N_VSS_XI0/XI34/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM8 N_XI0/XI34/XI0/NET35_XI0/XI34/XI0/MM8_d
+ N_WL<65>_XI0/XI34/XI0/MM8_g N_BLN<15>_XI0/XI34/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI0/MM5 N_XI0/XI34/XI0/NET34_XI0/XI34/XI0/MM5_d
+ N_XI0/XI34/XI0/NET33_XI0/XI34/XI0/MM5_g N_VDD_XI0/XI34/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI0/MM4 N_XI0/XI34/XI0/NET33_XI0/XI34/XI0/MM4_d
+ N_XI0/XI34/XI0/NET34_XI0/XI34/XI0/MM4_g N_VDD_XI0/XI34/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI0/MM10 N_XI0/XI34/XI0/NET35_XI0/XI34/XI0/MM10_d
+ N_XI0/XI34/XI0/NET36_XI0/XI34/XI0/MM10_g N_VDD_XI0/XI34/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI0/MM11 N_XI0/XI34/XI0/NET36_XI0/XI34/XI0/MM11_d
+ N_XI0/XI34/XI0/NET35_XI0/XI34/XI0/MM11_g N_VDD_XI0/XI34/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI1/MM2 N_XI0/XI34/XI1/NET34_XI0/XI34/XI1/MM2_d
+ N_XI0/XI34/XI1/NET33_XI0/XI34/XI1/MM2_g N_VSS_XI0/XI34/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM3 N_XI0/XI34/XI1/NET33_XI0/XI34/XI1/MM3_d
+ N_WL<64>_XI0/XI34/XI1/MM3_g N_BLN<14>_XI0/XI34/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM0 N_XI0/XI34/XI1/NET34_XI0/XI34/XI1/MM0_d
+ N_WL<64>_XI0/XI34/XI1/MM0_g N_BL<14>_XI0/XI34/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM1 N_XI0/XI34/XI1/NET33_XI0/XI34/XI1/MM1_d
+ N_XI0/XI34/XI1/NET34_XI0/XI34/XI1/MM1_g N_VSS_XI0/XI34/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM9 N_XI0/XI34/XI1/NET36_XI0/XI34/XI1/MM9_d
+ N_WL<65>_XI0/XI34/XI1/MM9_g N_BL<14>_XI0/XI34/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM6 N_XI0/XI34/XI1/NET35_XI0/XI34/XI1/MM6_d
+ N_XI0/XI34/XI1/NET36_XI0/XI34/XI1/MM6_g N_VSS_XI0/XI34/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM7 N_XI0/XI34/XI1/NET36_XI0/XI34/XI1/MM7_d
+ N_XI0/XI34/XI1/NET35_XI0/XI34/XI1/MM7_g N_VSS_XI0/XI34/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM8 N_XI0/XI34/XI1/NET35_XI0/XI34/XI1/MM8_d
+ N_WL<65>_XI0/XI34/XI1/MM8_g N_BLN<14>_XI0/XI34/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI1/MM5 N_XI0/XI34/XI1/NET34_XI0/XI34/XI1/MM5_d
+ N_XI0/XI34/XI1/NET33_XI0/XI34/XI1/MM5_g N_VDD_XI0/XI34/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI1/MM4 N_XI0/XI34/XI1/NET33_XI0/XI34/XI1/MM4_d
+ N_XI0/XI34/XI1/NET34_XI0/XI34/XI1/MM4_g N_VDD_XI0/XI34/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI1/MM10 N_XI0/XI34/XI1/NET35_XI0/XI34/XI1/MM10_d
+ N_XI0/XI34/XI1/NET36_XI0/XI34/XI1/MM10_g N_VDD_XI0/XI34/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI1/MM11 N_XI0/XI34/XI1/NET36_XI0/XI34/XI1/MM11_d
+ N_XI0/XI34/XI1/NET35_XI0/XI34/XI1/MM11_g N_VDD_XI0/XI34/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI2/MM2 N_XI0/XI34/XI2/NET34_XI0/XI34/XI2/MM2_d
+ N_XI0/XI34/XI2/NET33_XI0/XI34/XI2/MM2_g N_VSS_XI0/XI34/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM3 N_XI0/XI34/XI2/NET33_XI0/XI34/XI2/MM3_d
+ N_WL<64>_XI0/XI34/XI2/MM3_g N_BLN<13>_XI0/XI34/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM0 N_XI0/XI34/XI2/NET34_XI0/XI34/XI2/MM0_d
+ N_WL<64>_XI0/XI34/XI2/MM0_g N_BL<13>_XI0/XI34/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM1 N_XI0/XI34/XI2/NET33_XI0/XI34/XI2/MM1_d
+ N_XI0/XI34/XI2/NET34_XI0/XI34/XI2/MM1_g N_VSS_XI0/XI34/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM9 N_XI0/XI34/XI2/NET36_XI0/XI34/XI2/MM9_d
+ N_WL<65>_XI0/XI34/XI2/MM9_g N_BL<13>_XI0/XI34/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM6 N_XI0/XI34/XI2/NET35_XI0/XI34/XI2/MM6_d
+ N_XI0/XI34/XI2/NET36_XI0/XI34/XI2/MM6_g N_VSS_XI0/XI34/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM7 N_XI0/XI34/XI2/NET36_XI0/XI34/XI2/MM7_d
+ N_XI0/XI34/XI2/NET35_XI0/XI34/XI2/MM7_g N_VSS_XI0/XI34/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM8 N_XI0/XI34/XI2/NET35_XI0/XI34/XI2/MM8_d
+ N_WL<65>_XI0/XI34/XI2/MM8_g N_BLN<13>_XI0/XI34/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI2/MM5 N_XI0/XI34/XI2/NET34_XI0/XI34/XI2/MM5_d
+ N_XI0/XI34/XI2/NET33_XI0/XI34/XI2/MM5_g N_VDD_XI0/XI34/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI2/MM4 N_XI0/XI34/XI2/NET33_XI0/XI34/XI2/MM4_d
+ N_XI0/XI34/XI2/NET34_XI0/XI34/XI2/MM4_g N_VDD_XI0/XI34/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI2/MM10 N_XI0/XI34/XI2/NET35_XI0/XI34/XI2/MM10_d
+ N_XI0/XI34/XI2/NET36_XI0/XI34/XI2/MM10_g N_VDD_XI0/XI34/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI2/MM11 N_XI0/XI34/XI2/NET36_XI0/XI34/XI2/MM11_d
+ N_XI0/XI34/XI2/NET35_XI0/XI34/XI2/MM11_g N_VDD_XI0/XI34/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI3/MM2 N_XI0/XI34/XI3/NET34_XI0/XI34/XI3/MM2_d
+ N_XI0/XI34/XI3/NET33_XI0/XI34/XI3/MM2_g N_VSS_XI0/XI34/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM3 N_XI0/XI34/XI3/NET33_XI0/XI34/XI3/MM3_d
+ N_WL<64>_XI0/XI34/XI3/MM3_g N_BLN<12>_XI0/XI34/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM0 N_XI0/XI34/XI3/NET34_XI0/XI34/XI3/MM0_d
+ N_WL<64>_XI0/XI34/XI3/MM0_g N_BL<12>_XI0/XI34/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM1 N_XI0/XI34/XI3/NET33_XI0/XI34/XI3/MM1_d
+ N_XI0/XI34/XI3/NET34_XI0/XI34/XI3/MM1_g N_VSS_XI0/XI34/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM9 N_XI0/XI34/XI3/NET36_XI0/XI34/XI3/MM9_d
+ N_WL<65>_XI0/XI34/XI3/MM9_g N_BL<12>_XI0/XI34/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM6 N_XI0/XI34/XI3/NET35_XI0/XI34/XI3/MM6_d
+ N_XI0/XI34/XI3/NET36_XI0/XI34/XI3/MM6_g N_VSS_XI0/XI34/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM7 N_XI0/XI34/XI3/NET36_XI0/XI34/XI3/MM7_d
+ N_XI0/XI34/XI3/NET35_XI0/XI34/XI3/MM7_g N_VSS_XI0/XI34/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM8 N_XI0/XI34/XI3/NET35_XI0/XI34/XI3/MM8_d
+ N_WL<65>_XI0/XI34/XI3/MM8_g N_BLN<12>_XI0/XI34/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI3/MM5 N_XI0/XI34/XI3/NET34_XI0/XI34/XI3/MM5_d
+ N_XI0/XI34/XI3/NET33_XI0/XI34/XI3/MM5_g N_VDD_XI0/XI34/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI3/MM4 N_XI0/XI34/XI3/NET33_XI0/XI34/XI3/MM4_d
+ N_XI0/XI34/XI3/NET34_XI0/XI34/XI3/MM4_g N_VDD_XI0/XI34/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI3/MM10 N_XI0/XI34/XI3/NET35_XI0/XI34/XI3/MM10_d
+ N_XI0/XI34/XI3/NET36_XI0/XI34/XI3/MM10_g N_VDD_XI0/XI34/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI3/MM11 N_XI0/XI34/XI3/NET36_XI0/XI34/XI3/MM11_d
+ N_XI0/XI34/XI3/NET35_XI0/XI34/XI3/MM11_g N_VDD_XI0/XI34/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI4/MM2 N_XI0/XI34/XI4/NET34_XI0/XI34/XI4/MM2_d
+ N_XI0/XI34/XI4/NET33_XI0/XI34/XI4/MM2_g N_VSS_XI0/XI34/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM3 N_XI0/XI34/XI4/NET33_XI0/XI34/XI4/MM3_d
+ N_WL<64>_XI0/XI34/XI4/MM3_g N_BLN<11>_XI0/XI34/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM0 N_XI0/XI34/XI4/NET34_XI0/XI34/XI4/MM0_d
+ N_WL<64>_XI0/XI34/XI4/MM0_g N_BL<11>_XI0/XI34/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM1 N_XI0/XI34/XI4/NET33_XI0/XI34/XI4/MM1_d
+ N_XI0/XI34/XI4/NET34_XI0/XI34/XI4/MM1_g N_VSS_XI0/XI34/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM9 N_XI0/XI34/XI4/NET36_XI0/XI34/XI4/MM9_d
+ N_WL<65>_XI0/XI34/XI4/MM9_g N_BL<11>_XI0/XI34/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM6 N_XI0/XI34/XI4/NET35_XI0/XI34/XI4/MM6_d
+ N_XI0/XI34/XI4/NET36_XI0/XI34/XI4/MM6_g N_VSS_XI0/XI34/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM7 N_XI0/XI34/XI4/NET36_XI0/XI34/XI4/MM7_d
+ N_XI0/XI34/XI4/NET35_XI0/XI34/XI4/MM7_g N_VSS_XI0/XI34/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM8 N_XI0/XI34/XI4/NET35_XI0/XI34/XI4/MM8_d
+ N_WL<65>_XI0/XI34/XI4/MM8_g N_BLN<11>_XI0/XI34/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI4/MM5 N_XI0/XI34/XI4/NET34_XI0/XI34/XI4/MM5_d
+ N_XI0/XI34/XI4/NET33_XI0/XI34/XI4/MM5_g N_VDD_XI0/XI34/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI4/MM4 N_XI0/XI34/XI4/NET33_XI0/XI34/XI4/MM4_d
+ N_XI0/XI34/XI4/NET34_XI0/XI34/XI4/MM4_g N_VDD_XI0/XI34/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI4/MM10 N_XI0/XI34/XI4/NET35_XI0/XI34/XI4/MM10_d
+ N_XI0/XI34/XI4/NET36_XI0/XI34/XI4/MM10_g N_VDD_XI0/XI34/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI4/MM11 N_XI0/XI34/XI4/NET36_XI0/XI34/XI4/MM11_d
+ N_XI0/XI34/XI4/NET35_XI0/XI34/XI4/MM11_g N_VDD_XI0/XI34/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI5/MM2 N_XI0/XI34/XI5/NET34_XI0/XI34/XI5/MM2_d
+ N_XI0/XI34/XI5/NET33_XI0/XI34/XI5/MM2_g N_VSS_XI0/XI34/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM3 N_XI0/XI34/XI5/NET33_XI0/XI34/XI5/MM3_d
+ N_WL<64>_XI0/XI34/XI5/MM3_g N_BLN<10>_XI0/XI34/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM0 N_XI0/XI34/XI5/NET34_XI0/XI34/XI5/MM0_d
+ N_WL<64>_XI0/XI34/XI5/MM0_g N_BL<10>_XI0/XI34/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM1 N_XI0/XI34/XI5/NET33_XI0/XI34/XI5/MM1_d
+ N_XI0/XI34/XI5/NET34_XI0/XI34/XI5/MM1_g N_VSS_XI0/XI34/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM9 N_XI0/XI34/XI5/NET36_XI0/XI34/XI5/MM9_d
+ N_WL<65>_XI0/XI34/XI5/MM9_g N_BL<10>_XI0/XI34/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM6 N_XI0/XI34/XI5/NET35_XI0/XI34/XI5/MM6_d
+ N_XI0/XI34/XI5/NET36_XI0/XI34/XI5/MM6_g N_VSS_XI0/XI34/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM7 N_XI0/XI34/XI5/NET36_XI0/XI34/XI5/MM7_d
+ N_XI0/XI34/XI5/NET35_XI0/XI34/XI5/MM7_g N_VSS_XI0/XI34/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM8 N_XI0/XI34/XI5/NET35_XI0/XI34/XI5/MM8_d
+ N_WL<65>_XI0/XI34/XI5/MM8_g N_BLN<10>_XI0/XI34/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI5/MM5 N_XI0/XI34/XI5/NET34_XI0/XI34/XI5/MM5_d
+ N_XI0/XI34/XI5/NET33_XI0/XI34/XI5/MM5_g N_VDD_XI0/XI34/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI5/MM4 N_XI0/XI34/XI5/NET33_XI0/XI34/XI5/MM4_d
+ N_XI0/XI34/XI5/NET34_XI0/XI34/XI5/MM4_g N_VDD_XI0/XI34/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI5/MM10 N_XI0/XI34/XI5/NET35_XI0/XI34/XI5/MM10_d
+ N_XI0/XI34/XI5/NET36_XI0/XI34/XI5/MM10_g N_VDD_XI0/XI34/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI5/MM11 N_XI0/XI34/XI5/NET36_XI0/XI34/XI5/MM11_d
+ N_XI0/XI34/XI5/NET35_XI0/XI34/XI5/MM11_g N_VDD_XI0/XI34/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI6/MM2 N_XI0/XI34/XI6/NET34_XI0/XI34/XI6/MM2_d
+ N_XI0/XI34/XI6/NET33_XI0/XI34/XI6/MM2_g N_VSS_XI0/XI34/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM3 N_XI0/XI34/XI6/NET33_XI0/XI34/XI6/MM3_d
+ N_WL<64>_XI0/XI34/XI6/MM3_g N_BLN<9>_XI0/XI34/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM0 N_XI0/XI34/XI6/NET34_XI0/XI34/XI6/MM0_d
+ N_WL<64>_XI0/XI34/XI6/MM0_g N_BL<9>_XI0/XI34/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM1 N_XI0/XI34/XI6/NET33_XI0/XI34/XI6/MM1_d
+ N_XI0/XI34/XI6/NET34_XI0/XI34/XI6/MM1_g N_VSS_XI0/XI34/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM9 N_XI0/XI34/XI6/NET36_XI0/XI34/XI6/MM9_d
+ N_WL<65>_XI0/XI34/XI6/MM9_g N_BL<9>_XI0/XI34/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM6 N_XI0/XI34/XI6/NET35_XI0/XI34/XI6/MM6_d
+ N_XI0/XI34/XI6/NET36_XI0/XI34/XI6/MM6_g N_VSS_XI0/XI34/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM7 N_XI0/XI34/XI6/NET36_XI0/XI34/XI6/MM7_d
+ N_XI0/XI34/XI6/NET35_XI0/XI34/XI6/MM7_g N_VSS_XI0/XI34/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM8 N_XI0/XI34/XI6/NET35_XI0/XI34/XI6/MM8_d
+ N_WL<65>_XI0/XI34/XI6/MM8_g N_BLN<9>_XI0/XI34/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI6/MM5 N_XI0/XI34/XI6/NET34_XI0/XI34/XI6/MM5_d
+ N_XI0/XI34/XI6/NET33_XI0/XI34/XI6/MM5_g N_VDD_XI0/XI34/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI6/MM4 N_XI0/XI34/XI6/NET33_XI0/XI34/XI6/MM4_d
+ N_XI0/XI34/XI6/NET34_XI0/XI34/XI6/MM4_g N_VDD_XI0/XI34/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI6/MM10 N_XI0/XI34/XI6/NET35_XI0/XI34/XI6/MM10_d
+ N_XI0/XI34/XI6/NET36_XI0/XI34/XI6/MM10_g N_VDD_XI0/XI34/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI6/MM11 N_XI0/XI34/XI6/NET36_XI0/XI34/XI6/MM11_d
+ N_XI0/XI34/XI6/NET35_XI0/XI34/XI6/MM11_g N_VDD_XI0/XI34/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI7/MM2 N_XI0/XI34/XI7/NET34_XI0/XI34/XI7/MM2_d
+ N_XI0/XI34/XI7/NET33_XI0/XI34/XI7/MM2_g N_VSS_XI0/XI34/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM3 N_XI0/XI34/XI7/NET33_XI0/XI34/XI7/MM3_d
+ N_WL<64>_XI0/XI34/XI7/MM3_g N_BLN<8>_XI0/XI34/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM0 N_XI0/XI34/XI7/NET34_XI0/XI34/XI7/MM0_d
+ N_WL<64>_XI0/XI34/XI7/MM0_g N_BL<8>_XI0/XI34/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM1 N_XI0/XI34/XI7/NET33_XI0/XI34/XI7/MM1_d
+ N_XI0/XI34/XI7/NET34_XI0/XI34/XI7/MM1_g N_VSS_XI0/XI34/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM9 N_XI0/XI34/XI7/NET36_XI0/XI34/XI7/MM9_d
+ N_WL<65>_XI0/XI34/XI7/MM9_g N_BL<8>_XI0/XI34/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM6 N_XI0/XI34/XI7/NET35_XI0/XI34/XI7/MM6_d
+ N_XI0/XI34/XI7/NET36_XI0/XI34/XI7/MM6_g N_VSS_XI0/XI34/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM7 N_XI0/XI34/XI7/NET36_XI0/XI34/XI7/MM7_d
+ N_XI0/XI34/XI7/NET35_XI0/XI34/XI7/MM7_g N_VSS_XI0/XI34/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM8 N_XI0/XI34/XI7/NET35_XI0/XI34/XI7/MM8_d
+ N_WL<65>_XI0/XI34/XI7/MM8_g N_BLN<8>_XI0/XI34/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI7/MM5 N_XI0/XI34/XI7/NET34_XI0/XI34/XI7/MM5_d
+ N_XI0/XI34/XI7/NET33_XI0/XI34/XI7/MM5_g N_VDD_XI0/XI34/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI7/MM4 N_XI0/XI34/XI7/NET33_XI0/XI34/XI7/MM4_d
+ N_XI0/XI34/XI7/NET34_XI0/XI34/XI7/MM4_g N_VDD_XI0/XI34/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI7/MM10 N_XI0/XI34/XI7/NET35_XI0/XI34/XI7/MM10_d
+ N_XI0/XI34/XI7/NET36_XI0/XI34/XI7/MM10_g N_VDD_XI0/XI34/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI7/MM11 N_XI0/XI34/XI7/NET36_XI0/XI34/XI7/MM11_d
+ N_XI0/XI34/XI7/NET35_XI0/XI34/XI7/MM11_g N_VDD_XI0/XI34/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI8/MM2 N_XI0/XI34/XI8/NET34_XI0/XI34/XI8/MM2_d
+ N_XI0/XI34/XI8/NET33_XI0/XI34/XI8/MM2_g N_VSS_XI0/XI34/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM3 N_XI0/XI34/XI8/NET33_XI0/XI34/XI8/MM3_d
+ N_WL<64>_XI0/XI34/XI8/MM3_g N_BLN<7>_XI0/XI34/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM0 N_XI0/XI34/XI8/NET34_XI0/XI34/XI8/MM0_d
+ N_WL<64>_XI0/XI34/XI8/MM0_g N_BL<7>_XI0/XI34/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM1 N_XI0/XI34/XI8/NET33_XI0/XI34/XI8/MM1_d
+ N_XI0/XI34/XI8/NET34_XI0/XI34/XI8/MM1_g N_VSS_XI0/XI34/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM9 N_XI0/XI34/XI8/NET36_XI0/XI34/XI8/MM9_d
+ N_WL<65>_XI0/XI34/XI8/MM9_g N_BL<7>_XI0/XI34/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM6 N_XI0/XI34/XI8/NET35_XI0/XI34/XI8/MM6_d
+ N_XI0/XI34/XI8/NET36_XI0/XI34/XI8/MM6_g N_VSS_XI0/XI34/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM7 N_XI0/XI34/XI8/NET36_XI0/XI34/XI8/MM7_d
+ N_XI0/XI34/XI8/NET35_XI0/XI34/XI8/MM7_g N_VSS_XI0/XI34/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM8 N_XI0/XI34/XI8/NET35_XI0/XI34/XI8/MM8_d
+ N_WL<65>_XI0/XI34/XI8/MM8_g N_BLN<7>_XI0/XI34/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI8/MM5 N_XI0/XI34/XI8/NET34_XI0/XI34/XI8/MM5_d
+ N_XI0/XI34/XI8/NET33_XI0/XI34/XI8/MM5_g N_VDD_XI0/XI34/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI8/MM4 N_XI0/XI34/XI8/NET33_XI0/XI34/XI8/MM4_d
+ N_XI0/XI34/XI8/NET34_XI0/XI34/XI8/MM4_g N_VDD_XI0/XI34/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI8/MM10 N_XI0/XI34/XI8/NET35_XI0/XI34/XI8/MM10_d
+ N_XI0/XI34/XI8/NET36_XI0/XI34/XI8/MM10_g N_VDD_XI0/XI34/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI8/MM11 N_XI0/XI34/XI8/NET36_XI0/XI34/XI8/MM11_d
+ N_XI0/XI34/XI8/NET35_XI0/XI34/XI8/MM11_g N_VDD_XI0/XI34/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI9/MM2 N_XI0/XI34/XI9/NET34_XI0/XI34/XI9/MM2_d
+ N_XI0/XI34/XI9/NET33_XI0/XI34/XI9/MM2_g N_VSS_XI0/XI34/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM3 N_XI0/XI34/XI9/NET33_XI0/XI34/XI9/MM3_d
+ N_WL<64>_XI0/XI34/XI9/MM3_g N_BLN<6>_XI0/XI34/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM0 N_XI0/XI34/XI9/NET34_XI0/XI34/XI9/MM0_d
+ N_WL<64>_XI0/XI34/XI9/MM0_g N_BL<6>_XI0/XI34/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM1 N_XI0/XI34/XI9/NET33_XI0/XI34/XI9/MM1_d
+ N_XI0/XI34/XI9/NET34_XI0/XI34/XI9/MM1_g N_VSS_XI0/XI34/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM9 N_XI0/XI34/XI9/NET36_XI0/XI34/XI9/MM9_d
+ N_WL<65>_XI0/XI34/XI9/MM9_g N_BL<6>_XI0/XI34/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM6 N_XI0/XI34/XI9/NET35_XI0/XI34/XI9/MM6_d
+ N_XI0/XI34/XI9/NET36_XI0/XI34/XI9/MM6_g N_VSS_XI0/XI34/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM7 N_XI0/XI34/XI9/NET36_XI0/XI34/XI9/MM7_d
+ N_XI0/XI34/XI9/NET35_XI0/XI34/XI9/MM7_g N_VSS_XI0/XI34/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM8 N_XI0/XI34/XI9/NET35_XI0/XI34/XI9/MM8_d
+ N_WL<65>_XI0/XI34/XI9/MM8_g N_BLN<6>_XI0/XI34/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI9/MM5 N_XI0/XI34/XI9/NET34_XI0/XI34/XI9/MM5_d
+ N_XI0/XI34/XI9/NET33_XI0/XI34/XI9/MM5_g N_VDD_XI0/XI34/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI9/MM4 N_XI0/XI34/XI9/NET33_XI0/XI34/XI9/MM4_d
+ N_XI0/XI34/XI9/NET34_XI0/XI34/XI9/MM4_g N_VDD_XI0/XI34/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI9/MM10 N_XI0/XI34/XI9/NET35_XI0/XI34/XI9/MM10_d
+ N_XI0/XI34/XI9/NET36_XI0/XI34/XI9/MM10_g N_VDD_XI0/XI34/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI9/MM11 N_XI0/XI34/XI9/NET36_XI0/XI34/XI9/MM11_d
+ N_XI0/XI34/XI9/NET35_XI0/XI34/XI9/MM11_g N_VDD_XI0/XI34/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI10/MM2 N_XI0/XI34/XI10/NET34_XI0/XI34/XI10/MM2_d
+ N_XI0/XI34/XI10/NET33_XI0/XI34/XI10/MM2_g N_VSS_XI0/XI34/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM3 N_XI0/XI34/XI10/NET33_XI0/XI34/XI10/MM3_d
+ N_WL<64>_XI0/XI34/XI10/MM3_g N_BLN<5>_XI0/XI34/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM0 N_XI0/XI34/XI10/NET34_XI0/XI34/XI10/MM0_d
+ N_WL<64>_XI0/XI34/XI10/MM0_g N_BL<5>_XI0/XI34/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM1 N_XI0/XI34/XI10/NET33_XI0/XI34/XI10/MM1_d
+ N_XI0/XI34/XI10/NET34_XI0/XI34/XI10/MM1_g N_VSS_XI0/XI34/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM9 N_XI0/XI34/XI10/NET36_XI0/XI34/XI10/MM9_d
+ N_WL<65>_XI0/XI34/XI10/MM9_g N_BL<5>_XI0/XI34/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM6 N_XI0/XI34/XI10/NET35_XI0/XI34/XI10/MM6_d
+ N_XI0/XI34/XI10/NET36_XI0/XI34/XI10/MM6_g N_VSS_XI0/XI34/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM7 N_XI0/XI34/XI10/NET36_XI0/XI34/XI10/MM7_d
+ N_XI0/XI34/XI10/NET35_XI0/XI34/XI10/MM7_g N_VSS_XI0/XI34/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM8 N_XI0/XI34/XI10/NET35_XI0/XI34/XI10/MM8_d
+ N_WL<65>_XI0/XI34/XI10/MM8_g N_BLN<5>_XI0/XI34/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI10/MM5 N_XI0/XI34/XI10/NET34_XI0/XI34/XI10/MM5_d
+ N_XI0/XI34/XI10/NET33_XI0/XI34/XI10/MM5_g N_VDD_XI0/XI34/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI10/MM4 N_XI0/XI34/XI10/NET33_XI0/XI34/XI10/MM4_d
+ N_XI0/XI34/XI10/NET34_XI0/XI34/XI10/MM4_g N_VDD_XI0/XI34/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI10/MM10 N_XI0/XI34/XI10/NET35_XI0/XI34/XI10/MM10_d
+ N_XI0/XI34/XI10/NET36_XI0/XI34/XI10/MM10_g N_VDD_XI0/XI34/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI10/MM11 N_XI0/XI34/XI10/NET36_XI0/XI34/XI10/MM11_d
+ N_XI0/XI34/XI10/NET35_XI0/XI34/XI10/MM11_g N_VDD_XI0/XI34/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI11/MM2 N_XI0/XI34/XI11/NET34_XI0/XI34/XI11/MM2_d
+ N_XI0/XI34/XI11/NET33_XI0/XI34/XI11/MM2_g N_VSS_XI0/XI34/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM3 N_XI0/XI34/XI11/NET33_XI0/XI34/XI11/MM3_d
+ N_WL<64>_XI0/XI34/XI11/MM3_g N_BLN<4>_XI0/XI34/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM0 N_XI0/XI34/XI11/NET34_XI0/XI34/XI11/MM0_d
+ N_WL<64>_XI0/XI34/XI11/MM0_g N_BL<4>_XI0/XI34/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM1 N_XI0/XI34/XI11/NET33_XI0/XI34/XI11/MM1_d
+ N_XI0/XI34/XI11/NET34_XI0/XI34/XI11/MM1_g N_VSS_XI0/XI34/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM9 N_XI0/XI34/XI11/NET36_XI0/XI34/XI11/MM9_d
+ N_WL<65>_XI0/XI34/XI11/MM9_g N_BL<4>_XI0/XI34/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM6 N_XI0/XI34/XI11/NET35_XI0/XI34/XI11/MM6_d
+ N_XI0/XI34/XI11/NET36_XI0/XI34/XI11/MM6_g N_VSS_XI0/XI34/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM7 N_XI0/XI34/XI11/NET36_XI0/XI34/XI11/MM7_d
+ N_XI0/XI34/XI11/NET35_XI0/XI34/XI11/MM7_g N_VSS_XI0/XI34/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM8 N_XI0/XI34/XI11/NET35_XI0/XI34/XI11/MM8_d
+ N_WL<65>_XI0/XI34/XI11/MM8_g N_BLN<4>_XI0/XI34/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI11/MM5 N_XI0/XI34/XI11/NET34_XI0/XI34/XI11/MM5_d
+ N_XI0/XI34/XI11/NET33_XI0/XI34/XI11/MM5_g N_VDD_XI0/XI34/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI11/MM4 N_XI0/XI34/XI11/NET33_XI0/XI34/XI11/MM4_d
+ N_XI0/XI34/XI11/NET34_XI0/XI34/XI11/MM4_g N_VDD_XI0/XI34/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI11/MM10 N_XI0/XI34/XI11/NET35_XI0/XI34/XI11/MM10_d
+ N_XI0/XI34/XI11/NET36_XI0/XI34/XI11/MM10_g N_VDD_XI0/XI34/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI11/MM11 N_XI0/XI34/XI11/NET36_XI0/XI34/XI11/MM11_d
+ N_XI0/XI34/XI11/NET35_XI0/XI34/XI11/MM11_g N_VDD_XI0/XI34/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI12/MM2 N_XI0/XI34/XI12/NET34_XI0/XI34/XI12/MM2_d
+ N_XI0/XI34/XI12/NET33_XI0/XI34/XI12/MM2_g N_VSS_XI0/XI34/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM3 N_XI0/XI34/XI12/NET33_XI0/XI34/XI12/MM3_d
+ N_WL<64>_XI0/XI34/XI12/MM3_g N_BLN<3>_XI0/XI34/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM0 N_XI0/XI34/XI12/NET34_XI0/XI34/XI12/MM0_d
+ N_WL<64>_XI0/XI34/XI12/MM0_g N_BL<3>_XI0/XI34/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM1 N_XI0/XI34/XI12/NET33_XI0/XI34/XI12/MM1_d
+ N_XI0/XI34/XI12/NET34_XI0/XI34/XI12/MM1_g N_VSS_XI0/XI34/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM9 N_XI0/XI34/XI12/NET36_XI0/XI34/XI12/MM9_d
+ N_WL<65>_XI0/XI34/XI12/MM9_g N_BL<3>_XI0/XI34/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM6 N_XI0/XI34/XI12/NET35_XI0/XI34/XI12/MM6_d
+ N_XI0/XI34/XI12/NET36_XI0/XI34/XI12/MM6_g N_VSS_XI0/XI34/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM7 N_XI0/XI34/XI12/NET36_XI0/XI34/XI12/MM7_d
+ N_XI0/XI34/XI12/NET35_XI0/XI34/XI12/MM7_g N_VSS_XI0/XI34/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM8 N_XI0/XI34/XI12/NET35_XI0/XI34/XI12/MM8_d
+ N_WL<65>_XI0/XI34/XI12/MM8_g N_BLN<3>_XI0/XI34/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI12/MM5 N_XI0/XI34/XI12/NET34_XI0/XI34/XI12/MM5_d
+ N_XI0/XI34/XI12/NET33_XI0/XI34/XI12/MM5_g N_VDD_XI0/XI34/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI12/MM4 N_XI0/XI34/XI12/NET33_XI0/XI34/XI12/MM4_d
+ N_XI0/XI34/XI12/NET34_XI0/XI34/XI12/MM4_g N_VDD_XI0/XI34/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI12/MM10 N_XI0/XI34/XI12/NET35_XI0/XI34/XI12/MM10_d
+ N_XI0/XI34/XI12/NET36_XI0/XI34/XI12/MM10_g N_VDD_XI0/XI34/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI12/MM11 N_XI0/XI34/XI12/NET36_XI0/XI34/XI12/MM11_d
+ N_XI0/XI34/XI12/NET35_XI0/XI34/XI12/MM11_g N_VDD_XI0/XI34/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI13/MM2 N_XI0/XI34/XI13/NET34_XI0/XI34/XI13/MM2_d
+ N_XI0/XI34/XI13/NET33_XI0/XI34/XI13/MM2_g N_VSS_XI0/XI34/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM3 N_XI0/XI34/XI13/NET33_XI0/XI34/XI13/MM3_d
+ N_WL<64>_XI0/XI34/XI13/MM3_g N_BLN<2>_XI0/XI34/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM0 N_XI0/XI34/XI13/NET34_XI0/XI34/XI13/MM0_d
+ N_WL<64>_XI0/XI34/XI13/MM0_g N_BL<2>_XI0/XI34/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM1 N_XI0/XI34/XI13/NET33_XI0/XI34/XI13/MM1_d
+ N_XI0/XI34/XI13/NET34_XI0/XI34/XI13/MM1_g N_VSS_XI0/XI34/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM9 N_XI0/XI34/XI13/NET36_XI0/XI34/XI13/MM9_d
+ N_WL<65>_XI0/XI34/XI13/MM9_g N_BL<2>_XI0/XI34/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM6 N_XI0/XI34/XI13/NET35_XI0/XI34/XI13/MM6_d
+ N_XI0/XI34/XI13/NET36_XI0/XI34/XI13/MM6_g N_VSS_XI0/XI34/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM7 N_XI0/XI34/XI13/NET36_XI0/XI34/XI13/MM7_d
+ N_XI0/XI34/XI13/NET35_XI0/XI34/XI13/MM7_g N_VSS_XI0/XI34/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM8 N_XI0/XI34/XI13/NET35_XI0/XI34/XI13/MM8_d
+ N_WL<65>_XI0/XI34/XI13/MM8_g N_BLN<2>_XI0/XI34/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI13/MM5 N_XI0/XI34/XI13/NET34_XI0/XI34/XI13/MM5_d
+ N_XI0/XI34/XI13/NET33_XI0/XI34/XI13/MM5_g N_VDD_XI0/XI34/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI13/MM4 N_XI0/XI34/XI13/NET33_XI0/XI34/XI13/MM4_d
+ N_XI0/XI34/XI13/NET34_XI0/XI34/XI13/MM4_g N_VDD_XI0/XI34/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI13/MM10 N_XI0/XI34/XI13/NET35_XI0/XI34/XI13/MM10_d
+ N_XI0/XI34/XI13/NET36_XI0/XI34/XI13/MM10_g N_VDD_XI0/XI34/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI13/MM11 N_XI0/XI34/XI13/NET36_XI0/XI34/XI13/MM11_d
+ N_XI0/XI34/XI13/NET35_XI0/XI34/XI13/MM11_g N_VDD_XI0/XI34/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI14/MM2 N_XI0/XI34/XI14/NET34_XI0/XI34/XI14/MM2_d
+ N_XI0/XI34/XI14/NET33_XI0/XI34/XI14/MM2_g N_VSS_XI0/XI34/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM3 N_XI0/XI34/XI14/NET33_XI0/XI34/XI14/MM3_d
+ N_WL<64>_XI0/XI34/XI14/MM3_g N_BLN<1>_XI0/XI34/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM0 N_XI0/XI34/XI14/NET34_XI0/XI34/XI14/MM0_d
+ N_WL<64>_XI0/XI34/XI14/MM0_g N_BL<1>_XI0/XI34/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM1 N_XI0/XI34/XI14/NET33_XI0/XI34/XI14/MM1_d
+ N_XI0/XI34/XI14/NET34_XI0/XI34/XI14/MM1_g N_VSS_XI0/XI34/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM9 N_XI0/XI34/XI14/NET36_XI0/XI34/XI14/MM9_d
+ N_WL<65>_XI0/XI34/XI14/MM9_g N_BL<1>_XI0/XI34/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM6 N_XI0/XI34/XI14/NET35_XI0/XI34/XI14/MM6_d
+ N_XI0/XI34/XI14/NET36_XI0/XI34/XI14/MM6_g N_VSS_XI0/XI34/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM7 N_XI0/XI34/XI14/NET36_XI0/XI34/XI14/MM7_d
+ N_XI0/XI34/XI14/NET35_XI0/XI34/XI14/MM7_g N_VSS_XI0/XI34/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM8 N_XI0/XI34/XI14/NET35_XI0/XI34/XI14/MM8_d
+ N_WL<65>_XI0/XI34/XI14/MM8_g N_BLN<1>_XI0/XI34/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI14/MM5 N_XI0/XI34/XI14/NET34_XI0/XI34/XI14/MM5_d
+ N_XI0/XI34/XI14/NET33_XI0/XI34/XI14/MM5_g N_VDD_XI0/XI34/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI14/MM4 N_XI0/XI34/XI14/NET33_XI0/XI34/XI14/MM4_d
+ N_XI0/XI34/XI14/NET34_XI0/XI34/XI14/MM4_g N_VDD_XI0/XI34/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI14/MM10 N_XI0/XI34/XI14/NET35_XI0/XI34/XI14/MM10_d
+ N_XI0/XI34/XI14/NET36_XI0/XI34/XI14/MM10_g N_VDD_XI0/XI34/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI14/MM11 N_XI0/XI34/XI14/NET36_XI0/XI34/XI14/MM11_d
+ N_XI0/XI34/XI14/NET35_XI0/XI34/XI14/MM11_g N_VDD_XI0/XI34/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI15/MM2 N_XI0/XI34/XI15/NET34_XI0/XI34/XI15/MM2_d
+ N_XI0/XI34/XI15/NET33_XI0/XI34/XI15/MM2_g N_VSS_XI0/XI34/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM3 N_XI0/XI34/XI15/NET33_XI0/XI34/XI15/MM3_d
+ N_WL<64>_XI0/XI34/XI15/MM3_g N_BLN<0>_XI0/XI34/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM0 N_XI0/XI34/XI15/NET34_XI0/XI34/XI15/MM0_d
+ N_WL<64>_XI0/XI34/XI15/MM0_g N_BL<0>_XI0/XI34/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM1 N_XI0/XI34/XI15/NET33_XI0/XI34/XI15/MM1_d
+ N_XI0/XI34/XI15/NET34_XI0/XI34/XI15/MM1_g N_VSS_XI0/XI34/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM9 N_XI0/XI34/XI15/NET36_XI0/XI34/XI15/MM9_d
+ N_WL<65>_XI0/XI34/XI15/MM9_g N_BL<0>_XI0/XI34/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM6 N_XI0/XI34/XI15/NET35_XI0/XI34/XI15/MM6_d
+ N_XI0/XI34/XI15/NET36_XI0/XI34/XI15/MM6_g N_VSS_XI0/XI34/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM7 N_XI0/XI34/XI15/NET36_XI0/XI34/XI15/MM7_d
+ N_XI0/XI34/XI15/NET35_XI0/XI34/XI15/MM7_g N_VSS_XI0/XI34/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM8 N_XI0/XI34/XI15/NET35_XI0/XI34/XI15/MM8_d
+ N_WL<65>_XI0/XI34/XI15/MM8_g N_BLN<0>_XI0/XI34/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI34/XI15/MM5 N_XI0/XI34/XI15/NET34_XI0/XI34/XI15/MM5_d
+ N_XI0/XI34/XI15/NET33_XI0/XI34/XI15/MM5_g N_VDD_XI0/XI34/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI15/MM4 N_XI0/XI34/XI15/NET33_XI0/XI34/XI15/MM4_d
+ N_XI0/XI34/XI15/NET34_XI0/XI34/XI15/MM4_g N_VDD_XI0/XI34/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI15/MM10 N_XI0/XI34/XI15/NET35_XI0/XI34/XI15/MM10_d
+ N_XI0/XI34/XI15/NET36_XI0/XI34/XI15/MM10_g N_VDD_XI0/XI34/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI34/XI15/MM11 N_XI0/XI34/XI15/NET36_XI0/XI34/XI15/MM11_d
+ N_XI0/XI34/XI15/NET35_XI0/XI34/XI15/MM11_g N_VDD_XI0/XI34/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI0/MM2 N_XI0/XI35/XI0/NET34_XI0/XI35/XI0/MM2_d
+ N_XI0/XI35/XI0/NET33_XI0/XI35/XI0/MM2_g N_VSS_XI0/XI35/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM3 N_XI0/XI35/XI0/NET33_XI0/XI35/XI0/MM3_d
+ N_WL<66>_XI0/XI35/XI0/MM3_g N_BLN<15>_XI0/XI35/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM0 N_XI0/XI35/XI0/NET34_XI0/XI35/XI0/MM0_d
+ N_WL<66>_XI0/XI35/XI0/MM0_g N_BL<15>_XI0/XI35/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM1 N_XI0/XI35/XI0/NET33_XI0/XI35/XI0/MM1_d
+ N_XI0/XI35/XI0/NET34_XI0/XI35/XI0/MM1_g N_VSS_XI0/XI35/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM9 N_XI0/XI35/XI0/NET36_XI0/XI35/XI0/MM9_d
+ N_WL<67>_XI0/XI35/XI0/MM9_g N_BL<15>_XI0/XI35/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM6 N_XI0/XI35/XI0/NET35_XI0/XI35/XI0/MM6_d
+ N_XI0/XI35/XI0/NET36_XI0/XI35/XI0/MM6_g N_VSS_XI0/XI35/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM7 N_XI0/XI35/XI0/NET36_XI0/XI35/XI0/MM7_d
+ N_XI0/XI35/XI0/NET35_XI0/XI35/XI0/MM7_g N_VSS_XI0/XI35/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM8 N_XI0/XI35/XI0/NET35_XI0/XI35/XI0/MM8_d
+ N_WL<67>_XI0/XI35/XI0/MM8_g N_BLN<15>_XI0/XI35/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI0/MM5 N_XI0/XI35/XI0/NET34_XI0/XI35/XI0/MM5_d
+ N_XI0/XI35/XI0/NET33_XI0/XI35/XI0/MM5_g N_VDD_XI0/XI35/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI0/MM4 N_XI0/XI35/XI0/NET33_XI0/XI35/XI0/MM4_d
+ N_XI0/XI35/XI0/NET34_XI0/XI35/XI0/MM4_g N_VDD_XI0/XI35/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI0/MM10 N_XI0/XI35/XI0/NET35_XI0/XI35/XI0/MM10_d
+ N_XI0/XI35/XI0/NET36_XI0/XI35/XI0/MM10_g N_VDD_XI0/XI35/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI0/MM11 N_XI0/XI35/XI0/NET36_XI0/XI35/XI0/MM11_d
+ N_XI0/XI35/XI0/NET35_XI0/XI35/XI0/MM11_g N_VDD_XI0/XI35/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI1/MM2 N_XI0/XI35/XI1/NET34_XI0/XI35/XI1/MM2_d
+ N_XI0/XI35/XI1/NET33_XI0/XI35/XI1/MM2_g N_VSS_XI0/XI35/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM3 N_XI0/XI35/XI1/NET33_XI0/XI35/XI1/MM3_d
+ N_WL<66>_XI0/XI35/XI1/MM3_g N_BLN<14>_XI0/XI35/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM0 N_XI0/XI35/XI1/NET34_XI0/XI35/XI1/MM0_d
+ N_WL<66>_XI0/XI35/XI1/MM0_g N_BL<14>_XI0/XI35/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM1 N_XI0/XI35/XI1/NET33_XI0/XI35/XI1/MM1_d
+ N_XI0/XI35/XI1/NET34_XI0/XI35/XI1/MM1_g N_VSS_XI0/XI35/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM9 N_XI0/XI35/XI1/NET36_XI0/XI35/XI1/MM9_d
+ N_WL<67>_XI0/XI35/XI1/MM9_g N_BL<14>_XI0/XI35/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM6 N_XI0/XI35/XI1/NET35_XI0/XI35/XI1/MM6_d
+ N_XI0/XI35/XI1/NET36_XI0/XI35/XI1/MM6_g N_VSS_XI0/XI35/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM7 N_XI0/XI35/XI1/NET36_XI0/XI35/XI1/MM7_d
+ N_XI0/XI35/XI1/NET35_XI0/XI35/XI1/MM7_g N_VSS_XI0/XI35/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM8 N_XI0/XI35/XI1/NET35_XI0/XI35/XI1/MM8_d
+ N_WL<67>_XI0/XI35/XI1/MM8_g N_BLN<14>_XI0/XI35/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI1/MM5 N_XI0/XI35/XI1/NET34_XI0/XI35/XI1/MM5_d
+ N_XI0/XI35/XI1/NET33_XI0/XI35/XI1/MM5_g N_VDD_XI0/XI35/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI1/MM4 N_XI0/XI35/XI1/NET33_XI0/XI35/XI1/MM4_d
+ N_XI0/XI35/XI1/NET34_XI0/XI35/XI1/MM4_g N_VDD_XI0/XI35/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI1/MM10 N_XI0/XI35/XI1/NET35_XI0/XI35/XI1/MM10_d
+ N_XI0/XI35/XI1/NET36_XI0/XI35/XI1/MM10_g N_VDD_XI0/XI35/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI1/MM11 N_XI0/XI35/XI1/NET36_XI0/XI35/XI1/MM11_d
+ N_XI0/XI35/XI1/NET35_XI0/XI35/XI1/MM11_g N_VDD_XI0/XI35/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI2/MM2 N_XI0/XI35/XI2/NET34_XI0/XI35/XI2/MM2_d
+ N_XI0/XI35/XI2/NET33_XI0/XI35/XI2/MM2_g N_VSS_XI0/XI35/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM3 N_XI0/XI35/XI2/NET33_XI0/XI35/XI2/MM3_d
+ N_WL<66>_XI0/XI35/XI2/MM3_g N_BLN<13>_XI0/XI35/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM0 N_XI0/XI35/XI2/NET34_XI0/XI35/XI2/MM0_d
+ N_WL<66>_XI0/XI35/XI2/MM0_g N_BL<13>_XI0/XI35/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM1 N_XI0/XI35/XI2/NET33_XI0/XI35/XI2/MM1_d
+ N_XI0/XI35/XI2/NET34_XI0/XI35/XI2/MM1_g N_VSS_XI0/XI35/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM9 N_XI0/XI35/XI2/NET36_XI0/XI35/XI2/MM9_d
+ N_WL<67>_XI0/XI35/XI2/MM9_g N_BL<13>_XI0/XI35/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM6 N_XI0/XI35/XI2/NET35_XI0/XI35/XI2/MM6_d
+ N_XI0/XI35/XI2/NET36_XI0/XI35/XI2/MM6_g N_VSS_XI0/XI35/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM7 N_XI0/XI35/XI2/NET36_XI0/XI35/XI2/MM7_d
+ N_XI0/XI35/XI2/NET35_XI0/XI35/XI2/MM7_g N_VSS_XI0/XI35/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM8 N_XI0/XI35/XI2/NET35_XI0/XI35/XI2/MM8_d
+ N_WL<67>_XI0/XI35/XI2/MM8_g N_BLN<13>_XI0/XI35/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI2/MM5 N_XI0/XI35/XI2/NET34_XI0/XI35/XI2/MM5_d
+ N_XI0/XI35/XI2/NET33_XI0/XI35/XI2/MM5_g N_VDD_XI0/XI35/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI2/MM4 N_XI0/XI35/XI2/NET33_XI0/XI35/XI2/MM4_d
+ N_XI0/XI35/XI2/NET34_XI0/XI35/XI2/MM4_g N_VDD_XI0/XI35/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI2/MM10 N_XI0/XI35/XI2/NET35_XI0/XI35/XI2/MM10_d
+ N_XI0/XI35/XI2/NET36_XI0/XI35/XI2/MM10_g N_VDD_XI0/XI35/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI2/MM11 N_XI0/XI35/XI2/NET36_XI0/XI35/XI2/MM11_d
+ N_XI0/XI35/XI2/NET35_XI0/XI35/XI2/MM11_g N_VDD_XI0/XI35/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI3/MM2 N_XI0/XI35/XI3/NET34_XI0/XI35/XI3/MM2_d
+ N_XI0/XI35/XI3/NET33_XI0/XI35/XI3/MM2_g N_VSS_XI0/XI35/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM3 N_XI0/XI35/XI3/NET33_XI0/XI35/XI3/MM3_d
+ N_WL<66>_XI0/XI35/XI3/MM3_g N_BLN<12>_XI0/XI35/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM0 N_XI0/XI35/XI3/NET34_XI0/XI35/XI3/MM0_d
+ N_WL<66>_XI0/XI35/XI3/MM0_g N_BL<12>_XI0/XI35/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM1 N_XI0/XI35/XI3/NET33_XI0/XI35/XI3/MM1_d
+ N_XI0/XI35/XI3/NET34_XI0/XI35/XI3/MM1_g N_VSS_XI0/XI35/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM9 N_XI0/XI35/XI3/NET36_XI0/XI35/XI3/MM9_d
+ N_WL<67>_XI0/XI35/XI3/MM9_g N_BL<12>_XI0/XI35/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM6 N_XI0/XI35/XI3/NET35_XI0/XI35/XI3/MM6_d
+ N_XI0/XI35/XI3/NET36_XI0/XI35/XI3/MM6_g N_VSS_XI0/XI35/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM7 N_XI0/XI35/XI3/NET36_XI0/XI35/XI3/MM7_d
+ N_XI0/XI35/XI3/NET35_XI0/XI35/XI3/MM7_g N_VSS_XI0/XI35/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM8 N_XI0/XI35/XI3/NET35_XI0/XI35/XI3/MM8_d
+ N_WL<67>_XI0/XI35/XI3/MM8_g N_BLN<12>_XI0/XI35/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI3/MM5 N_XI0/XI35/XI3/NET34_XI0/XI35/XI3/MM5_d
+ N_XI0/XI35/XI3/NET33_XI0/XI35/XI3/MM5_g N_VDD_XI0/XI35/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI3/MM4 N_XI0/XI35/XI3/NET33_XI0/XI35/XI3/MM4_d
+ N_XI0/XI35/XI3/NET34_XI0/XI35/XI3/MM4_g N_VDD_XI0/XI35/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI3/MM10 N_XI0/XI35/XI3/NET35_XI0/XI35/XI3/MM10_d
+ N_XI0/XI35/XI3/NET36_XI0/XI35/XI3/MM10_g N_VDD_XI0/XI35/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI3/MM11 N_XI0/XI35/XI3/NET36_XI0/XI35/XI3/MM11_d
+ N_XI0/XI35/XI3/NET35_XI0/XI35/XI3/MM11_g N_VDD_XI0/XI35/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI4/MM2 N_XI0/XI35/XI4/NET34_XI0/XI35/XI4/MM2_d
+ N_XI0/XI35/XI4/NET33_XI0/XI35/XI4/MM2_g N_VSS_XI0/XI35/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM3 N_XI0/XI35/XI4/NET33_XI0/XI35/XI4/MM3_d
+ N_WL<66>_XI0/XI35/XI4/MM3_g N_BLN<11>_XI0/XI35/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM0 N_XI0/XI35/XI4/NET34_XI0/XI35/XI4/MM0_d
+ N_WL<66>_XI0/XI35/XI4/MM0_g N_BL<11>_XI0/XI35/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM1 N_XI0/XI35/XI4/NET33_XI0/XI35/XI4/MM1_d
+ N_XI0/XI35/XI4/NET34_XI0/XI35/XI4/MM1_g N_VSS_XI0/XI35/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM9 N_XI0/XI35/XI4/NET36_XI0/XI35/XI4/MM9_d
+ N_WL<67>_XI0/XI35/XI4/MM9_g N_BL<11>_XI0/XI35/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM6 N_XI0/XI35/XI4/NET35_XI0/XI35/XI4/MM6_d
+ N_XI0/XI35/XI4/NET36_XI0/XI35/XI4/MM6_g N_VSS_XI0/XI35/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM7 N_XI0/XI35/XI4/NET36_XI0/XI35/XI4/MM7_d
+ N_XI0/XI35/XI4/NET35_XI0/XI35/XI4/MM7_g N_VSS_XI0/XI35/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM8 N_XI0/XI35/XI4/NET35_XI0/XI35/XI4/MM8_d
+ N_WL<67>_XI0/XI35/XI4/MM8_g N_BLN<11>_XI0/XI35/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI4/MM5 N_XI0/XI35/XI4/NET34_XI0/XI35/XI4/MM5_d
+ N_XI0/XI35/XI4/NET33_XI0/XI35/XI4/MM5_g N_VDD_XI0/XI35/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI4/MM4 N_XI0/XI35/XI4/NET33_XI0/XI35/XI4/MM4_d
+ N_XI0/XI35/XI4/NET34_XI0/XI35/XI4/MM4_g N_VDD_XI0/XI35/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI4/MM10 N_XI0/XI35/XI4/NET35_XI0/XI35/XI4/MM10_d
+ N_XI0/XI35/XI4/NET36_XI0/XI35/XI4/MM10_g N_VDD_XI0/XI35/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI4/MM11 N_XI0/XI35/XI4/NET36_XI0/XI35/XI4/MM11_d
+ N_XI0/XI35/XI4/NET35_XI0/XI35/XI4/MM11_g N_VDD_XI0/XI35/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI5/MM2 N_XI0/XI35/XI5/NET34_XI0/XI35/XI5/MM2_d
+ N_XI0/XI35/XI5/NET33_XI0/XI35/XI5/MM2_g N_VSS_XI0/XI35/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM3 N_XI0/XI35/XI5/NET33_XI0/XI35/XI5/MM3_d
+ N_WL<66>_XI0/XI35/XI5/MM3_g N_BLN<10>_XI0/XI35/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM0 N_XI0/XI35/XI5/NET34_XI0/XI35/XI5/MM0_d
+ N_WL<66>_XI0/XI35/XI5/MM0_g N_BL<10>_XI0/XI35/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM1 N_XI0/XI35/XI5/NET33_XI0/XI35/XI5/MM1_d
+ N_XI0/XI35/XI5/NET34_XI0/XI35/XI5/MM1_g N_VSS_XI0/XI35/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM9 N_XI0/XI35/XI5/NET36_XI0/XI35/XI5/MM9_d
+ N_WL<67>_XI0/XI35/XI5/MM9_g N_BL<10>_XI0/XI35/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM6 N_XI0/XI35/XI5/NET35_XI0/XI35/XI5/MM6_d
+ N_XI0/XI35/XI5/NET36_XI0/XI35/XI5/MM6_g N_VSS_XI0/XI35/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM7 N_XI0/XI35/XI5/NET36_XI0/XI35/XI5/MM7_d
+ N_XI0/XI35/XI5/NET35_XI0/XI35/XI5/MM7_g N_VSS_XI0/XI35/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM8 N_XI0/XI35/XI5/NET35_XI0/XI35/XI5/MM8_d
+ N_WL<67>_XI0/XI35/XI5/MM8_g N_BLN<10>_XI0/XI35/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI5/MM5 N_XI0/XI35/XI5/NET34_XI0/XI35/XI5/MM5_d
+ N_XI0/XI35/XI5/NET33_XI0/XI35/XI5/MM5_g N_VDD_XI0/XI35/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI5/MM4 N_XI0/XI35/XI5/NET33_XI0/XI35/XI5/MM4_d
+ N_XI0/XI35/XI5/NET34_XI0/XI35/XI5/MM4_g N_VDD_XI0/XI35/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI5/MM10 N_XI0/XI35/XI5/NET35_XI0/XI35/XI5/MM10_d
+ N_XI0/XI35/XI5/NET36_XI0/XI35/XI5/MM10_g N_VDD_XI0/XI35/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI5/MM11 N_XI0/XI35/XI5/NET36_XI0/XI35/XI5/MM11_d
+ N_XI0/XI35/XI5/NET35_XI0/XI35/XI5/MM11_g N_VDD_XI0/XI35/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI6/MM2 N_XI0/XI35/XI6/NET34_XI0/XI35/XI6/MM2_d
+ N_XI0/XI35/XI6/NET33_XI0/XI35/XI6/MM2_g N_VSS_XI0/XI35/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM3 N_XI0/XI35/XI6/NET33_XI0/XI35/XI6/MM3_d
+ N_WL<66>_XI0/XI35/XI6/MM3_g N_BLN<9>_XI0/XI35/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM0 N_XI0/XI35/XI6/NET34_XI0/XI35/XI6/MM0_d
+ N_WL<66>_XI0/XI35/XI6/MM0_g N_BL<9>_XI0/XI35/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM1 N_XI0/XI35/XI6/NET33_XI0/XI35/XI6/MM1_d
+ N_XI0/XI35/XI6/NET34_XI0/XI35/XI6/MM1_g N_VSS_XI0/XI35/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM9 N_XI0/XI35/XI6/NET36_XI0/XI35/XI6/MM9_d
+ N_WL<67>_XI0/XI35/XI6/MM9_g N_BL<9>_XI0/XI35/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM6 N_XI0/XI35/XI6/NET35_XI0/XI35/XI6/MM6_d
+ N_XI0/XI35/XI6/NET36_XI0/XI35/XI6/MM6_g N_VSS_XI0/XI35/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM7 N_XI0/XI35/XI6/NET36_XI0/XI35/XI6/MM7_d
+ N_XI0/XI35/XI6/NET35_XI0/XI35/XI6/MM7_g N_VSS_XI0/XI35/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM8 N_XI0/XI35/XI6/NET35_XI0/XI35/XI6/MM8_d
+ N_WL<67>_XI0/XI35/XI6/MM8_g N_BLN<9>_XI0/XI35/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI6/MM5 N_XI0/XI35/XI6/NET34_XI0/XI35/XI6/MM5_d
+ N_XI0/XI35/XI6/NET33_XI0/XI35/XI6/MM5_g N_VDD_XI0/XI35/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI6/MM4 N_XI0/XI35/XI6/NET33_XI0/XI35/XI6/MM4_d
+ N_XI0/XI35/XI6/NET34_XI0/XI35/XI6/MM4_g N_VDD_XI0/XI35/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI6/MM10 N_XI0/XI35/XI6/NET35_XI0/XI35/XI6/MM10_d
+ N_XI0/XI35/XI6/NET36_XI0/XI35/XI6/MM10_g N_VDD_XI0/XI35/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI6/MM11 N_XI0/XI35/XI6/NET36_XI0/XI35/XI6/MM11_d
+ N_XI0/XI35/XI6/NET35_XI0/XI35/XI6/MM11_g N_VDD_XI0/XI35/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI7/MM2 N_XI0/XI35/XI7/NET34_XI0/XI35/XI7/MM2_d
+ N_XI0/XI35/XI7/NET33_XI0/XI35/XI7/MM2_g N_VSS_XI0/XI35/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM3 N_XI0/XI35/XI7/NET33_XI0/XI35/XI7/MM3_d
+ N_WL<66>_XI0/XI35/XI7/MM3_g N_BLN<8>_XI0/XI35/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM0 N_XI0/XI35/XI7/NET34_XI0/XI35/XI7/MM0_d
+ N_WL<66>_XI0/XI35/XI7/MM0_g N_BL<8>_XI0/XI35/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM1 N_XI0/XI35/XI7/NET33_XI0/XI35/XI7/MM1_d
+ N_XI0/XI35/XI7/NET34_XI0/XI35/XI7/MM1_g N_VSS_XI0/XI35/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM9 N_XI0/XI35/XI7/NET36_XI0/XI35/XI7/MM9_d
+ N_WL<67>_XI0/XI35/XI7/MM9_g N_BL<8>_XI0/XI35/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM6 N_XI0/XI35/XI7/NET35_XI0/XI35/XI7/MM6_d
+ N_XI0/XI35/XI7/NET36_XI0/XI35/XI7/MM6_g N_VSS_XI0/XI35/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM7 N_XI0/XI35/XI7/NET36_XI0/XI35/XI7/MM7_d
+ N_XI0/XI35/XI7/NET35_XI0/XI35/XI7/MM7_g N_VSS_XI0/XI35/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM8 N_XI0/XI35/XI7/NET35_XI0/XI35/XI7/MM8_d
+ N_WL<67>_XI0/XI35/XI7/MM8_g N_BLN<8>_XI0/XI35/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI7/MM5 N_XI0/XI35/XI7/NET34_XI0/XI35/XI7/MM5_d
+ N_XI0/XI35/XI7/NET33_XI0/XI35/XI7/MM5_g N_VDD_XI0/XI35/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI7/MM4 N_XI0/XI35/XI7/NET33_XI0/XI35/XI7/MM4_d
+ N_XI0/XI35/XI7/NET34_XI0/XI35/XI7/MM4_g N_VDD_XI0/XI35/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI7/MM10 N_XI0/XI35/XI7/NET35_XI0/XI35/XI7/MM10_d
+ N_XI0/XI35/XI7/NET36_XI0/XI35/XI7/MM10_g N_VDD_XI0/XI35/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI7/MM11 N_XI0/XI35/XI7/NET36_XI0/XI35/XI7/MM11_d
+ N_XI0/XI35/XI7/NET35_XI0/XI35/XI7/MM11_g N_VDD_XI0/XI35/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI8/MM2 N_XI0/XI35/XI8/NET34_XI0/XI35/XI8/MM2_d
+ N_XI0/XI35/XI8/NET33_XI0/XI35/XI8/MM2_g N_VSS_XI0/XI35/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM3 N_XI0/XI35/XI8/NET33_XI0/XI35/XI8/MM3_d
+ N_WL<66>_XI0/XI35/XI8/MM3_g N_BLN<7>_XI0/XI35/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM0 N_XI0/XI35/XI8/NET34_XI0/XI35/XI8/MM0_d
+ N_WL<66>_XI0/XI35/XI8/MM0_g N_BL<7>_XI0/XI35/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM1 N_XI0/XI35/XI8/NET33_XI0/XI35/XI8/MM1_d
+ N_XI0/XI35/XI8/NET34_XI0/XI35/XI8/MM1_g N_VSS_XI0/XI35/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM9 N_XI0/XI35/XI8/NET36_XI0/XI35/XI8/MM9_d
+ N_WL<67>_XI0/XI35/XI8/MM9_g N_BL<7>_XI0/XI35/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM6 N_XI0/XI35/XI8/NET35_XI0/XI35/XI8/MM6_d
+ N_XI0/XI35/XI8/NET36_XI0/XI35/XI8/MM6_g N_VSS_XI0/XI35/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM7 N_XI0/XI35/XI8/NET36_XI0/XI35/XI8/MM7_d
+ N_XI0/XI35/XI8/NET35_XI0/XI35/XI8/MM7_g N_VSS_XI0/XI35/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM8 N_XI0/XI35/XI8/NET35_XI0/XI35/XI8/MM8_d
+ N_WL<67>_XI0/XI35/XI8/MM8_g N_BLN<7>_XI0/XI35/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI8/MM5 N_XI0/XI35/XI8/NET34_XI0/XI35/XI8/MM5_d
+ N_XI0/XI35/XI8/NET33_XI0/XI35/XI8/MM5_g N_VDD_XI0/XI35/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI8/MM4 N_XI0/XI35/XI8/NET33_XI0/XI35/XI8/MM4_d
+ N_XI0/XI35/XI8/NET34_XI0/XI35/XI8/MM4_g N_VDD_XI0/XI35/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI8/MM10 N_XI0/XI35/XI8/NET35_XI0/XI35/XI8/MM10_d
+ N_XI0/XI35/XI8/NET36_XI0/XI35/XI8/MM10_g N_VDD_XI0/XI35/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI8/MM11 N_XI0/XI35/XI8/NET36_XI0/XI35/XI8/MM11_d
+ N_XI0/XI35/XI8/NET35_XI0/XI35/XI8/MM11_g N_VDD_XI0/XI35/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI9/MM2 N_XI0/XI35/XI9/NET34_XI0/XI35/XI9/MM2_d
+ N_XI0/XI35/XI9/NET33_XI0/XI35/XI9/MM2_g N_VSS_XI0/XI35/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM3 N_XI0/XI35/XI9/NET33_XI0/XI35/XI9/MM3_d
+ N_WL<66>_XI0/XI35/XI9/MM3_g N_BLN<6>_XI0/XI35/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM0 N_XI0/XI35/XI9/NET34_XI0/XI35/XI9/MM0_d
+ N_WL<66>_XI0/XI35/XI9/MM0_g N_BL<6>_XI0/XI35/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM1 N_XI0/XI35/XI9/NET33_XI0/XI35/XI9/MM1_d
+ N_XI0/XI35/XI9/NET34_XI0/XI35/XI9/MM1_g N_VSS_XI0/XI35/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM9 N_XI0/XI35/XI9/NET36_XI0/XI35/XI9/MM9_d
+ N_WL<67>_XI0/XI35/XI9/MM9_g N_BL<6>_XI0/XI35/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM6 N_XI0/XI35/XI9/NET35_XI0/XI35/XI9/MM6_d
+ N_XI0/XI35/XI9/NET36_XI0/XI35/XI9/MM6_g N_VSS_XI0/XI35/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM7 N_XI0/XI35/XI9/NET36_XI0/XI35/XI9/MM7_d
+ N_XI0/XI35/XI9/NET35_XI0/XI35/XI9/MM7_g N_VSS_XI0/XI35/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM8 N_XI0/XI35/XI9/NET35_XI0/XI35/XI9/MM8_d
+ N_WL<67>_XI0/XI35/XI9/MM8_g N_BLN<6>_XI0/XI35/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI9/MM5 N_XI0/XI35/XI9/NET34_XI0/XI35/XI9/MM5_d
+ N_XI0/XI35/XI9/NET33_XI0/XI35/XI9/MM5_g N_VDD_XI0/XI35/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI9/MM4 N_XI0/XI35/XI9/NET33_XI0/XI35/XI9/MM4_d
+ N_XI0/XI35/XI9/NET34_XI0/XI35/XI9/MM4_g N_VDD_XI0/XI35/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI9/MM10 N_XI0/XI35/XI9/NET35_XI0/XI35/XI9/MM10_d
+ N_XI0/XI35/XI9/NET36_XI0/XI35/XI9/MM10_g N_VDD_XI0/XI35/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI9/MM11 N_XI0/XI35/XI9/NET36_XI0/XI35/XI9/MM11_d
+ N_XI0/XI35/XI9/NET35_XI0/XI35/XI9/MM11_g N_VDD_XI0/XI35/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI10/MM2 N_XI0/XI35/XI10/NET34_XI0/XI35/XI10/MM2_d
+ N_XI0/XI35/XI10/NET33_XI0/XI35/XI10/MM2_g N_VSS_XI0/XI35/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM3 N_XI0/XI35/XI10/NET33_XI0/XI35/XI10/MM3_d
+ N_WL<66>_XI0/XI35/XI10/MM3_g N_BLN<5>_XI0/XI35/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM0 N_XI0/XI35/XI10/NET34_XI0/XI35/XI10/MM0_d
+ N_WL<66>_XI0/XI35/XI10/MM0_g N_BL<5>_XI0/XI35/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM1 N_XI0/XI35/XI10/NET33_XI0/XI35/XI10/MM1_d
+ N_XI0/XI35/XI10/NET34_XI0/XI35/XI10/MM1_g N_VSS_XI0/XI35/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM9 N_XI0/XI35/XI10/NET36_XI0/XI35/XI10/MM9_d
+ N_WL<67>_XI0/XI35/XI10/MM9_g N_BL<5>_XI0/XI35/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM6 N_XI0/XI35/XI10/NET35_XI0/XI35/XI10/MM6_d
+ N_XI0/XI35/XI10/NET36_XI0/XI35/XI10/MM6_g N_VSS_XI0/XI35/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM7 N_XI0/XI35/XI10/NET36_XI0/XI35/XI10/MM7_d
+ N_XI0/XI35/XI10/NET35_XI0/XI35/XI10/MM7_g N_VSS_XI0/XI35/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM8 N_XI0/XI35/XI10/NET35_XI0/XI35/XI10/MM8_d
+ N_WL<67>_XI0/XI35/XI10/MM8_g N_BLN<5>_XI0/XI35/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI10/MM5 N_XI0/XI35/XI10/NET34_XI0/XI35/XI10/MM5_d
+ N_XI0/XI35/XI10/NET33_XI0/XI35/XI10/MM5_g N_VDD_XI0/XI35/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI10/MM4 N_XI0/XI35/XI10/NET33_XI0/XI35/XI10/MM4_d
+ N_XI0/XI35/XI10/NET34_XI0/XI35/XI10/MM4_g N_VDD_XI0/XI35/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI10/MM10 N_XI0/XI35/XI10/NET35_XI0/XI35/XI10/MM10_d
+ N_XI0/XI35/XI10/NET36_XI0/XI35/XI10/MM10_g N_VDD_XI0/XI35/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI10/MM11 N_XI0/XI35/XI10/NET36_XI0/XI35/XI10/MM11_d
+ N_XI0/XI35/XI10/NET35_XI0/XI35/XI10/MM11_g N_VDD_XI0/XI35/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI11/MM2 N_XI0/XI35/XI11/NET34_XI0/XI35/XI11/MM2_d
+ N_XI0/XI35/XI11/NET33_XI0/XI35/XI11/MM2_g N_VSS_XI0/XI35/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM3 N_XI0/XI35/XI11/NET33_XI0/XI35/XI11/MM3_d
+ N_WL<66>_XI0/XI35/XI11/MM3_g N_BLN<4>_XI0/XI35/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM0 N_XI0/XI35/XI11/NET34_XI0/XI35/XI11/MM0_d
+ N_WL<66>_XI0/XI35/XI11/MM0_g N_BL<4>_XI0/XI35/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM1 N_XI0/XI35/XI11/NET33_XI0/XI35/XI11/MM1_d
+ N_XI0/XI35/XI11/NET34_XI0/XI35/XI11/MM1_g N_VSS_XI0/XI35/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM9 N_XI0/XI35/XI11/NET36_XI0/XI35/XI11/MM9_d
+ N_WL<67>_XI0/XI35/XI11/MM9_g N_BL<4>_XI0/XI35/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM6 N_XI0/XI35/XI11/NET35_XI0/XI35/XI11/MM6_d
+ N_XI0/XI35/XI11/NET36_XI0/XI35/XI11/MM6_g N_VSS_XI0/XI35/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM7 N_XI0/XI35/XI11/NET36_XI0/XI35/XI11/MM7_d
+ N_XI0/XI35/XI11/NET35_XI0/XI35/XI11/MM7_g N_VSS_XI0/XI35/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM8 N_XI0/XI35/XI11/NET35_XI0/XI35/XI11/MM8_d
+ N_WL<67>_XI0/XI35/XI11/MM8_g N_BLN<4>_XI0/XI35/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI11/MM5 N_XI0/XI35/XI11/NET34_XI0/XI35/XI11/MM5_d
+ N_XI0/XI35/XI11/NET33_XI0/XI35/XI11/MM5_g N_VDD_XI0/XI35/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI11/MM4 N_XI0/XI35/XI11/NET33_XI0/XI35/XI11/MM4_d
+ N_XI0/XI35/XI11/NET34_XI0/XI35/XI11/MM4_g N_VDD_XI0/XI35/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI11/MM10 N_XI0/XI35/XI11/NET35_XI0/XI35/XI11/MM10_d
+ N_XI0/XI35/XI11/NET36_XI0/XI35/XI11/MM10_g N_VDD_XI0/XI35/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI11/MM11 N_XI0/XI35/XI11/NET36_XI0/XI35/XI11/MM11_d
+ N_XI0/XI35/XI11/NET35_XI0/XI35/XI11/MM11_g N_VDD_XI0/XI35/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI12/MM2 N_XI0/XI35/XI12/NET34_XI0/XI35/XI12/MM2_d
+ N_XI0/XI35/XI12/NET33_XI0/XI35/XI12/MM2_g N_VSS_XI0/XI35/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM3 N_XI0/XI35/XI12/NET33_XI0/XI35/XI12/MM3_d
+ N_WL<66>_XI0/XI35/XI12/MM3_g N_BLN<3>_XI0/XI35/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM0 N_XI0/XI35/XI12/NET34_XI0/XI35/XI12/MM0_d
+ N_WL<66>_XI0/XI35/XI12/MM0_g N_BL<3>_XI0/XI35/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM1 N_XI0/XI35/XI12/NET33_XI0/XI35/XI12/MM1_d
+ N_XI0/XI35/XI12/NET34_XI0/XI35/XI12/MM1_g N_VSS_XI0/XI35/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM9 N_XI0/XI35/XI12/NET36_XI0/XI35/XI12/MM9_d
+ N_WL<67>_XI0/XI35/XI12/MM9_g N_BL<3>_XI0/XI35/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM6 N_XI0/XI35/XI12/NET35_XI0/XI35/XI12/MM6_d
+ N_XI0/XI35/XI12/NET36_XI0/XI35/XI12/MM6_g N_VSS_XI0/XI35/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM7 N_XI0/XI35/XI12/NET36_XI0/XI35/XI12/MM7_d
+ N_XI0/XI35/XI12/NET35_XI0/XI35/XI12/MM7_g N_VSS_XI0/XI35/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM8 N_XI0/XI35/XI12/NET35_XI0/XI35/XI12/MM8_d
+ N_WL<67>_XI0/XI35/XI12/MM8_g N_BLN<3>_XI0/XI35/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI12/MM5 N_XI0/XI35/XI12/NET34_XI0/XI35/XI12/MM5_d
+ N_XI0/XI35/XI12/NET33_XI0/XI35/XI12/MM5_g N_VDD_XI0/XI35/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI12/MM4 N_XI0/XI35/XI12/NET33_XI0/XI35/XI12/MM4_d
+ N_XI0/XI35/XI12/NET34_XI0/XI35/XI12/MM4_g N_VDD_XI0/XI35/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI12/MM10 N_XI0/XI35/XI12/NET35_XI0/XI35/XI12/MM10_d
+ N_XI0/XI35/XI12/NET36_XI0/XI35/XI12/MM10_g N_VDD_XI0/XI35/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI12/MM11 N_XI0/XI35/XI12/NET36_XI0/XI35/XI12/MM11_d
+ N_XI0/XI35/XI12/NET35_XI0/XI35/XI12/MM11_g N_VDD_XI0/XI35/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI13/MM2 N_XI0/XI35/XI13/NET34_XI0/XI35/XI13/MM2_d
+ N_XI0/XI35/XI13/NET33_XI0/XI35/XI13/MM2_g N_VSS_XI0/XI35/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM3 N_XI0/XI35/XI13/NET33_XI0/XI35/XI13/MM3_d
+ N_WL<66>_XI0/XI35/XI13/MM3_g N_BLN<2>_XI0/XI35/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM0 N_XI0/XI35/XI13/NET34_XI0/XI35/XI13/MM0_d
+ N_WL<66>_XI0/XI35/XI13/MM0_g N_BL<2>_XI0/XI35/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM1 N_XI0/XI35/XI13/NET33_XI0/XI35/XI13/MM1_d
+ N_XI0/XI35/XI13/NET34_XI0/XI35/XI13/MM1_g N_VSS_XI0/XI35/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM9 N_XI0/XI35/XI13/NET36_XI0/XI35/XI13/MM9_d
+ N_WL<67>_XI0/XI35/XI13/MM9_g N_BL<2>_XI0/XI35/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM6 N_XI0/XI35/XI13/NET35_XI0/XI35/XI13/MM6_d
+ N_XI0/XI35/XI13/NET36_XI0/XI35/XI13/MM6_g N_VSS_XI0/XI35/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM7 N_XI0/XI35/XI13/NET36_XI0/XI35/XI13/MM7_d
+ N_XI0/XI35/XI13/NET35_XI0/XI35/XI13/MM7_g N_VSS_XI0/XI35/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM8 N_XI0/XI35/XI13/NET35_XI0/XI35/XI13/MM8_d
+ N_WL<67>_XI0/XI35/XI13/MM8_g N_BLN<2>_XI0/XI35/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI13/MM5 N_XI0/XI35/XI13/NET34_XI0/XI35/XI13/MM5_d
+ N_XI0/XI35/XI13/NET33_XI0/XI35/XI13/MM5_g N_VDD_XI0/XI35/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI13/MM4 N_XI0/XI35/XI13/NET33_XI0/XI35/XI13/MM4_d
+ N_XI0/XI35/XI13/NET34_XI0/XI35/XI13/MM4_g N_VDD_XI0/XI35/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI13/MM10 N_XI0/XI35/XI13/NET35_XI0/XI35/XI13/MM10_d
+ N_XI0/XI35/XI13/NET36_XI0/XI35/XI13/MM10_g N_VDD_XI0/XI35/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI13/MM11 N_XI0/XI35/XI13/NET36_XI0/XI35/XI13/MM11_d
+ N_XI0/XI35/XI13/NET35_XI0/XI35/XI13/MM11_g N_VDD_XI0/XI35/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI14/MM2 N_XI0/XI35/XI14/NET34_XI0/XI35/XI14/MM2_d
+ N_XI0/XI35/XI14/NET33_XI0/XI35/XI14/MM2_g N_VSS_XI0/XI35/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM3 N_XI0/XI35/XI14/NET33_XI0/XI35/XI14/MM3_d
+ N_WL<66>_XI0/XI35/XI14/MM3_g N_BLN<1>_XI0/XI35/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM0 N_XI0/XI35/XI14/NET34_XI0/XI35/XI14/MM0_d
+ N_WL<66>_XI0/XI35/XI14/MM0_g N_BL<1>_XI0/XI35/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM1 N_XI0/XI35/XI14/NET33_XI0/XI35/XI14/MM1_d
+ N_XI0/XI35/XI14/NET34_XI0/XI35/XI14/MM1_g N_VSS_XI0/XI35/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM9 N_XI0/XI35/XI14/NET36_XI0/XI35/XI14/MM9_d
+ N_WL<67>_XI0/XI35/XI14/MM9_g N_BL<1>_XI0/XI35/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM6 N_XI0/XI35/XI14/NET35_XI0/XI35/XI14/MM6_d
+ N_XI0/XI35/XI14/NET36_XI0/XI35/XI14/MM6_g N_VSS_XI0/XI35/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM7 N_XI0/XI35/XI14/NET36_XI0/XI35/XI14/MM7_d
+ N_XI0/XI35/XI14/NET35_XI0/XI35/XI14/MM7_g N_VSS_XI0/XI35/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM8 N_XI0/XI35/XI14/NET35_XI0/XI35/XI14/MM8_d
+ N_WL<67>_XI0/XI35/XI14/MM8_g N_BLN<1>_XI0/XI35/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI14/MM5 N_XI0/XI35/XI14/NET34_XI0/XI35/XI14/MM5_d
+ N_XI0/XI35/XI14/NET33_XI0/XI35/XI14/MM5_g N_VDD_XI0/XI35/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI14/MM4 N_XI0/XI35/XI14/NET33_XI0/XI35/XI14/MM4_d
+ N_XI0/XI35/XI14/NET34_XI0/XI35/XI14/MM4_g N_VDD_XI0/XI35/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI14/MM10 N_XI0/XI35/XI14/NET35_XI0/XI35/XI14/MM10_d
+ N_XI0/XI35/XI14/NET36_XI0/XI35/XI14/MM10_g N_VDD_XI0/XI35/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI14/MM11 N_XI0/XI35/XI14/NET36_XI0/XI35/XI14/MM11_d
+ N_XI0/XI35/XI14/NET35_XI0/XI35/XI14/MM11_g N_VDD_XI0/XI35/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI15/MM2 N_XI0/XI35/XI15/NET34_XI0/XI35/XI15/MM2_d
+ N_XI0/XI35/XI15/NET33_XI0/XI35/XI15/MM2_g N_VSS_XI0/XI35/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM3 N_XI0/XI35/XI15/NET33_XI0/XI35/XI15/MM3_d
+ N_WL<66>_XI0/XI35/XI15/MM3_g N_BLN<0>_XI0/XI35/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM0 N_XI0/XI35/XI15/NET34_XI0/XI35/XI15/MM0_d
+ N_WL<66>_XI0/XI35/XI15/MM0_g N_BL<0>_XI0/XI35/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM1 N_XI0/XI35/XI15/NET33_XI0/XI35/XI15/MM1_d
+ N_XI0/XI35/XI15/NET34_XI0/XI35/XI15/MM1_g N_VSS_XI0/XI35/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM9 N_XI0/XI35/XI15/NET36_XI0/XI35/XI15/MM9_d
+ N_WL<67>_XI0/XI35/XI15/MM9_g N_BL<0>_XI0/XI35/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM6 N_XI0/XI35/XI15/NET35_XI0/XI35/XI15/MM6_d
+ N_XI0/XI35/XI15/NET36_XI0/XI35/XI15/MM6_g N_VSS_XI0/XI35/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM7 N_XI0/XI35/XI15/NET36_XI0/XI35/XI15/MM7_d
+ N_XI0/XI35/XI15/NET35_XI0/XI35/XI15/MM7_g N_VSS_XI0/XI35/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM8 N_XI0/XI35/XI15/NET35_XI0/XI35/XI15/MM8_d
+ N_WL<67>_XI0/XI35/XI15/MM8_g N_BLN<0>_XI0/XI35/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI35/XI15/MM5 N_XI0/XI35/XI15/NET34_XI0/XI35/XI15/MM5_d
+ N_XI0/XI35/XI15/NET33_XI0/XI35/XI15/MM5_g N_VDD_XI0/XI35/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI15/MM4 N_XI0/XI35/XI15/NET33_XI0/XI35/XI15/MM4_d
+ N_XI0/XI35/XI15/NET34_XI0/XI35/XI15/MM4_g N_VDD_XI0/XI35/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI15/MM10 N_XI0/XI35/XI15/NET35_XI0/XI35/XI15/MM10_d
+ N_XI0/XI35/XI15/NET36_XI0/XI35/XI15/MM10_g N_VDD_XI0/XI35/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI35/XI15/MM11 N_XI0/XI35/XI15/NET36_XI0/XI35/XI15/MM11_d
+ N_XI0/XI35/XI15/NET35_XI0/XI35/XI15/MM11_g N_VDD_XI0/XI35/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI0/MM2 N_XI0/XI36/XI0/NET34_XI0/XI36/XI0/MM2_d
+ N_XI0/XI36/XI0/NET33_XI0/XI36/XI0/MM2_g N_VSS_XI0/XI36/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM3 N_XI0/XI36/XI0/NET33_XI0/XI36/XI0/MM3_d
+ N_WL<68>_XI0/XI36/XI0/MM3_g N_BLN<15>_XI0/XI36/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM0 N_XI0/XI36/XI0/NET34_XI0/XI36/XI0/MM0_d
+ N_WL<68>_XI0/XI36/XI0/MM0_g N_BL<15>_XI0/XI36/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM1 N_XI0/XI36/XI0/NET33_XI0/XI36/XI0/MM1_d
+ N_XI0/XI36/XI0/NET34_XI0/XI36/XI0/MM1_g N_VSS_XI0/XI36/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM9 N_XI0/XI36/XI0/NET36_XI0/XI36/XI0/MM9_d
+ N_WL<69>_XI0/XI36/XI0/MM9_g N_BL<15>_XI0/XI36/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM6 N_XI0/XI36/XI0/NET35_XI0/XI36/XI0/MM6_d
+ N_XI0/XI36/XI0/NET36_XI0/XI36/XI0/MM6_g N_VSS_XI0/XI36/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM7 N_XI0/XI36/XI0/NET36_XI0/XI36/XI0/MM7_d
+ N_XI0/XI36/XI0/NET35_XI0/XI36/XI0/MM7_g N_VSS_XI0/XI36/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM8 N_XI0/XI36/XI0/NET35_XI0/XI36/XI0/MM8_d
+ N_WL<69>_XI0/XI36/XI0/MM8_g N_BLN<15>_XI0/XI36/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI0/MM5 N_XI0/XI36/XI0/NET34_XI0/XI36/XI0/MM5_d
+ N_XI0/XI36/XI0/NET33_XI0/XI36/XI0/MM5_g N_VDD_XI0/XI36/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI0/MM4 N_XI0/XI36/XI0/NET33_XI0/XI36/XI0/MM4_d
+ N_XI0/XI36/XI0/NET34_XI0/XI36/XI0/MM4_g N_VDD_XI0/XI36/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI0/MM10 N_XI0/XI36/XI0/NET35_XI0/XI36/XI0/MM10_d
+ N_XI0/XI36/XI0/NET36_XI0/XI36/XI0/MM10_g N_VDD_XI0/XI36/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI0/MM11 N_XI0/XI36/XI0/NET36_XI0/XI36/XI0/MM11_d
+ N_XI0/XI36/XI0/NET35_XI0/XI36/XI0/MM11_g N_VDD_XI0/XI36/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI1/MM2 N_XI0/XI36/XI1/NET34_XI0/XI36/XI1/MM2_d
+ N_XI0/XI36/XI1/NET33_XI0/XI36/XI1/MM2_g N_VSS_XI0/XI36/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM3 N_XI0/XI36/XI1/NET33_XI0/XI36/XI1/MM3_d
+ N_WL<68>_XI0/XI36/XI1/MM3_g N_BLN<14>_XI0/XI36/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM0 N_XI0/XI36/XI1/NET34_XI0/XI36/XI1/MM0_d
+ N_WL<68>_XI0/XI36/XI1/MM0_g N_BL<14>_XI0/XI36/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM1 N_XI0/XI36/XI1/NET33_XI0/XI36/XI1/MM1_d
+ N_XI0/XI36/XI1/NET34_XI0/XI36/XI1/MM1_g N_VSS_XI0/XI36/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM9 N_XI0/XI36/XI1/NET36_XI0/XI36/XI1/MM9_d
+ N_WL<69>_XI0/XI36/XI1/MM9_g N_BL<14>_XI0/XI36/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM6 N_XI0/XI36/XI1/NET35_XI0/XI36/XI1/MM6_d
+ N_XI0/XI36/XI1/NET36_XI0/XI36/XI1/MM6_g N_VSS_XI0/XI36/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM7 N_XI0/XI36/XI1/NET36_XI0/XI36/XI1/MM7_d
+ N_XI0/XI36/XI1/NET35_XI0/XI36/XI1/MM7_g N_VSS_XI0/XI36/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM8 N_XI0/XI36/XI1/NET35_XI0/XI36/XI1/MM8_d
+ N_WL<69>_XI0/XI36/XI1/MM8_g N_BLN<14>_XI0/XI36/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI1/MM5 N_XI0/XI36/XI1/NET34_XI0/XI36/XI1/MM5_d
+ N_XI0/XI36/XI1/NET33_XI0/XI36/XI1/MM5_g N_VDD_XI0/XI36/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI1/MM4 N_XI0/XI36/XI1/NET33_XI0/XI36/XI1/MM4_d
+ N_XI0/XI36/XI1/NET34_XI0/XI36/XI1/MM4_g N_VDD_XI0/XI36/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI1/MM10 N_XI0/XI36/XI1/NET35_XI0/XI36/XI1/MM10_d
+ N_XI0/XI36/XI1/NET36_XI0/XI36/XI1/MM10_g N_VDD_XI0/XI36/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI1/MM11 N_XI0/XI36/XI1/NET36_XI0/XI36/XI1/MM11_d
+ N_XI0/XI36/XI1/NET35_XI0/XI36/XI1/MM11_g N_VDD_XI0/XI36/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI2/MM2 N_XI0/XI36/XI2/NET34_XI0/XI36/XI2/MM2_d
+ N_XI0/XI36/XI2/NET33_XI0/XI36/XI2/MM2_g N_VSS_XI0/XI36/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM3 N_XI0/XI36/XI2/NET33_XI0/XI36/XI2/MM3_d
+ N_WL<68>_XI0/XI36/XI2/MM3_g N_BLN<13>_XI0/XI36/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM0 N_XI0/XI36/XI2/NET34_XI0/XI36/XI2/MM0_d
+ N_WL<68>_XI0/XI36/XI2/MM0_g N_BL<13>_XI0/XI36/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM1 N_XI0/XI36/XI2/NET33_XI0/XI36/XI2/MM1_d
+ N_XI0/XI36/XI2/NET34_XI0/XI36/XI2/MM1_g N_VSS_XI0/XI36/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM9 N_XI0/XI36/XI2/NET36_XI0/XI36/XI2/MM9_d
+ N_WL<69>_XI0/XI36/XI2/MM9_g N_BL<13>_XI0/XI36/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM6 N_XI0/XI36/XI2/NET35_XI0/XI36/XI2/MM6_d
+ N_XI0/XI36/XI2/NET36_XI0/XI36/XI2/MM6_g N_VSS_XI0/XI36/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM7 N_XI0/XI36/XI2/NET36_XI0/XI36/XI2/MM7_d
+ N_XI0/XI36/XI2/NET35_XI0/XI36/XI2/MM7_g N_VSS_XI0/XI36/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM8 N_XI0/XI36/XI2/NET35_XI0/XI36/XI2/MM8_d
+ N_WL<69>_XI0/XI36/XI2/MM8_g N_BLN<13>_XI0/XI36/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI2/MM5 N_XI0/XI36/XI2/NET34_XI0/XI36/XI2/MM5_d
+ N_XI0/XI36/XI2/NET33_XI0/XI36/XI2/MM5_g N_VDD_XI0/XI36/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI2/MM4 N_XI0/XI36/XI2/NET33_XI0/XI36/XI2/MM4_d
+ N_XI0/XI36/XI2/NET34_XI0/XI36/XI2/MM4_g N_VDD_XI0/XI36/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI2/MM10 N_XI0/XI36/XI2/NET35_XI0/XI36/XI2/MM10_d
+ N_XI0/XI36/XI2/NET36_XI0/XI36/XI2/MM10_g N_VDD_XI0/XI36/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI2/MM11 N_XI0/XI36/XI2/NET36_XI0/XI36/XI2/MM11_d
+ N_XI0/XI36/XI2/NET35_XI0/XI36/XI2/MM11_g N_VDD_XI0/XI36/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI3/MM2 N_XI0/XI36/XI3/NET34_XI0/XI36/XI3/MM2_d
+ N_XI0/XI36/XI3/NET33_XI0/XI36/XI3/MM2_g N_VSS_XI0/XI36/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM3 N_XI0/XI36/XI3/NET33_XI0/XI36/XI3/MM3_d
+ N_WL<68>_XI0/XI36/XI3/MM3_g N_BLN<12>_XI0/XI36/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM0 N_XI0/XI36/XI3/NET34_XI0/XI36/XI3/MM0_d
+ N_WL<68>_XI0/XI36/XI3/MM0_g N_BL<12>_XI0/XI36/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM1 N_XI0/XI36/XI3/NET33_XI0/XI36/XI3/MM1_d
+ N_XI0/XI36/XI3/NET34_XI0/XI36/XI3/MM1_g N_VSS_XI0/XI36/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM9 N_XI0/XI36/XI3/NET36_XI0/XI36/XI3/MM9_d
+ N_WL<69>_XI0/XI36/XI3/MM9_g N_BL<12>_XI0/XI36/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM6 N_XI0/XI36/XI3/NET35_XI0/XI36/XI3/MM6_d
+ N_XI0/XI36/XI3/NET36_XI0/XI36/XI3/MM6_g N_VSS_XI0/XI36/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM7 N_XI0/XI36/XI3/NET36_XI0/XI36/XI3/MM7_d
+ N_XI0/XI36/XI3/NET35_XI0/XI36/XI3/MM7_g N_VSS_XI0/XI36/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM8 N_XI0/XI36/XI3/NET35_XI0/XI36/XI3/MM8_d
+ N_WL<69>_XI0/XI36/XI3/MM8_g N_BLN<12>_XI0/XI36/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI3/MM5 N_XI0/XI36/XI3/NET34_XI0/XI36/XI3/MM5_d
+ N_XI0/XI36/XI3/NET33_XI0/XI36/XI3/MM5_g N_VDD_XI0/XI36/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI3/MM4 N_XI0/XI36/XI3/NET33_XI0/XI36/XI3/MM4_d
+ N_XI0/XI36/XI3/NET34_XI0/XI36/XI3/MM4_g N_VDD_XI0/XI36/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI3/MM10 N_XI0/XI36/XI3/NET35_XI0/XI36/XI3/MM10_d
+ N_XI0/XI36/XI3/NET36_XI0/XI36/XI3/MM10_g N_VDD_XI0/XI36/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI3/MM11 N_XI0/XI36/XI3/NET36_XI0/XI36/XI3/MM11_d
+ N_XI0/XI36/XI3/NET35_XI0/XI36/XI3/MM11_g N_VDD_XI0/XI36/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI4/MM2 N_XI0/XI36/XI4/NET34_XI0/XI36/XI4/MM2_d
+ N_XI0/XI36/XI4/NET33_XI0/XI36/XI4/MM2_g N_VSS_XI0/XI36/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM3 N_XI0/XI36/XI4/NET33_XI0/XI36/XI4/MM3_d
+ N_WL<68>_XI0/XI36/XI4/MM3_g N_BLN<11>_XI0/XI36/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM0 N_XI0/XI36/XI4/NET34_XI0/XI36/XI4/MM0_d
+ N_WL<68>_XI0/XI36/XI4/MM0_g N_BL<11>_XI0/XI36/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM1 N_XI0/XI36/XI4/NET33_XI0/XI36/XI4/MM1_d
+ N_XI0/XI36/XI4/NET34_XI0/XI36/XI4/MM1_g N_VSS_XI0/XI36/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM9 N_XI0/XI36/XI4/NET36_XI0/XI36/XI4/MM9_d
+ N_WL<69>_XI0/XI36/XI4/MM9_g N_BL<11>_XI0/XI36/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM6 N_XI0/XI36/XI4/NET35_XI0/XI36/XI4/MM6_d
+ N_XI0/XI36/XI4/NET36_XI0/XI36/XI4/MM6_g N_VSS_XI0/XI36/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM7 N_XI0/XI36/XI4/NET36_XI0/XI36/XI4/MM7_d
+ N_XI0/XI36/XI4/NET35_XI0/XI36/XI4/MM7_g N_VSS_XI0/XI36/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM8 N_XI0/XI36/XI4/NET35_XI0/XI36/XI4/MM8_d
+ N_WL<69>_XI0/XI36/XI4/MM8_g N_BLN<11>_XI0/XI36/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI4/MM5 N_XI0/XI36/XI4/NET34_XI0/XI36/XI4/MM5_d
+ N_XI0/XI36/XI4/NET33_XI0/XI36/XI4/MM5_g N_VDD_XI0/XI36/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI4/MM4 N_XI0/XI36/XI4/NET33_XI0/XI36/XI4/MM4_d
+ N_XI0/XI36/XI4/NET34_XI0/XI36/XI4/MM4_g N_VDD_XI0/XI36/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI4/MM10 N_XI0/XI36/XI4/NET35_XI0/XI36/XI4/MM10_d
+ N_XI0/XI36/XI4/NET36_XI0/XI36/XI4/MM10_g N_VDD_XI0/XI36/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI4/MM11 N_XI0/XI36/XI4/NET36_XI0/XI36/XI4/MM11_d
+ N_XI0/XI36/XI4/NET35_XI0/XI36/XI4/MM11_g N_VDD_XI0/XI36/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI5/MM2 N_XI0/XI36/XI5/NET34_XI0/XI36/XI5/MM2_d
+ N_XI0/XI36/XI5/NET33_XI0/XI36/XI5/MM2_g N_VSS_XI0/XI36/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM3 N_XI0/XI36/XI5/NET33_XI0/XI36/XI5/MM3_d
+ N_WL<68>_XI0/XI36/XI5/MM3_g N_BLN<10>_XI0/XI36/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM0 N_XI0/XI36/XI5/NET34_XI0/XI36/XI5/MM0_d
+ N_WL<68>_XI0/XI36/XI5/MM0_g N_BL<10>_XI0/XI36/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM1 N_XI0/XI36/XI5/NET33_XI0/XI36/XI5/MM1_d
+ N_XI0/XI36/XI5/NET34_XI0/XI36/XI5/MM1_g N_VSS_XI0/XI36/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM9 N_XI0/XI36/XI5/NET36_XI0/XI36/XI5/MM9_d
+ N_WL<69>_XI0/XI36/XI5/MM9_g N_BL<10>_XI0/XI36/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM6 N_XI0/XI36/XI5/NET35_XI0/XI36/XI5/MM6_d
+ N_XI0/XI36/XI5/NET36_XI0/XI36/XI5/MM6_g N_VSS_XI0/XI36/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM7 N_XI0/XI36/XI5/NET36_XI0/XI36/XI5/MM7_d
+ N_XI0/XI36/XI5/NET35_XI0/XI36/XI5/MM7_g N_VSS_XI0/XI36/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM8 N_XI0/XI36/XI5/NET35_XI0/XI36/XI5/MM8_d
+ N_WL<69>_XI0/XI36/XI5/MM8_g N_BLN<10>_XI0/XI36/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI5/MM5 N_XI0/XI36/XI5/NET34_XI0/XI36/XI5/MM5_d
+ N_XI0/XI36/XI5/NET33_XI0/XI36/XI5/MM5_g N_VDD_XI0/XI36/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI5/MM4 N_XI0/XI36/XI5/NET33_XI0/XI36/XI5/MM4_d
+ N_XI0/XI36/XI5/NET34_XI0/XI36/XI5/MM4_g N_VDD_XI0/XI36/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI5/MM10 N_XI0/XI36/XI5/NET35_XI0/XI36/XI5/MM10_d
+ N_XI0/XI36/XI5/NET36_XI0/XI36/XI5/MM10_g N_VDD_XI0/XI36/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI5/MM11 N_XI0/XI36/XI5/NET36_XI0/XI36/XI5/MM11_d
+ N_XI0/XI36/XI5/NET35_XI0/XI36/XI5/MM11_g N_VDD_XI0/XI36/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI6/MM2 N_XI0/XI36/XI6/NET34_XI0/XI36/XI6/MM2_d
+ N_XI0/XI36/XI6/NET33_XI0/XI36/XI6/MM2_g N_VSS_XI0/XI36/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM3 N_XI0/XI36/XI6/NET33_XI0/XI36/XI6/MM3_d
+ N_WL<68>_XI0/XI36/XI6/MM3_g N_BLN<9>_XI0/XI36/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM0 N_XI0/XI36/XI6/NET34_XI0/XI36/XI6/MM0_d
+ N_WL<68>_XI0/XI36/XI6/MM0_g N_BL<9>_XI0/XI36/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM1 N_XI0/XI36/XI6/NET33_XI0/XI36/XI6/MM1_d
+ N_XI0/XI36/XI6/NET34_XI0/XI36/XI6/MM1_g N_VSS_XI0/XI36/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM9 N_XI0/XI36/XI6/NET36_XI0/XI36/XI6/MM9_d
+ N_WL<69>_XI0/XI36/XI6/MM9_g N_BL<9>_XI0/XI36/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM6 N_XI0/XI36/XI6/NET35_XI0/XI36/XI6/MM6_d
+ N_XI0/XI36/XI6/NET36_XI0/XI36/XI6/MM6_g N_VSS_XI0/XI36/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM7 N_XI0/XI36/XI6/NET36_XI0/XI36/XI6/MM7_d
+ N_XI0/XI36/XI6/NET35_XI0/XI36/XI6/MM7_g N_VSS_XI0/XI36/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM8 N_XI0/XI36/XI6/NET35_XI0/XI36/XI6/MM8_d
+ N_WL<69>_XI0/XI36/XI6/MM8_g N_BLN<9>_XI0/XI36/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI6/MM5 N_XI0/XI36/XI6/NET34_XI0/XI36/XI6/MM5_d
+ N_XI0/XI36/XI6/NET33_XI0/XI36/XI6/MM5_g N_VDD_XI0/XI36/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI6/MM4 N_XI0/XI36/XI6/NET33_XI0/XI36/XI6/MM4_d
+ N_XI0/XI36/XI6/NET34_XI0/XI36/XI6/MM4_g N_VDD_XI0/XI36/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI6/MM10 N_XI0/XI36/XI6/NET35_XI0/XI36/XI6/MM10_d
+ N_XI0/XI36/XI6/NET36_XI0/XI36/XI6/MM10_g N_VDD_XI0/XI36/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI6/MM11 N_XI0/XI36/XI6/NET36_XI0/XI36/XI6/MM11_d
+ N_XI0/XI36/XI6/NET35_XI0/XI36/XI6/MM11_g N_VDD_XI0/XI36/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI7/MM2 N_XI0/XI36/XI7/NET34_XI0/XI36/XI7/MM2_d
+ N_XI0/XI36/XI7/NET33_XI0/XI36/XI7/MM2_g N_VSS_XI0/XI36/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM3 N_XI0/XI36/XI7/NET33_XI0/XI36/XI7/MM3_d
+ N_WL<68>_XI0/XI36/XI7/MM3_g N_BLN<8>_XI0/XI36/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM0 N_XI0/XI36/XI7/NET34_XI0/XI36/XI7/MM0_d
+ N_WL<68>_XI0/XI36/XI7/MM0_g N_BL<8>_XI0/XI36/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM1 N_XI0/XI36/XI7/NET33_XI0/XI36/XI7/MM1_d
+ N_XI0/XI36/XI7/NET34_XI0/XI36/XI7/MM1_g N_VSS_XI0/XI36/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM9 N_XI0/XI36/XI7/NET36_XI0/XI36/XI7/MM9_d
+ N_WL<69>_XI0/XI36/XI7/MM9_g N_BL<8>_XI0/XI36/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM6 N_XI0/XI36/XI7/NET35_XI0/XI36/XI7/MM6_d
+ N_XI0/XI36/XI7/NET36_XI0/XI36/XI7/MM6_g N_VSS_XI0/XI36/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM7 N_XI0/XI36/XI7/NET36_XI0/XI36/XI7/MM7_d
+ N_XI0/XI36/XI7/NET35_XI0/XI36/XI7/MM7_g N_VSS_XI0/XI36/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM8 N_XI0/XI36/XI7/NET35_XI0/XI36/XI7/MM8_d
+ N_WL<69>_XI0/XI36/XI7/MM8_g N_BLN<8>_XI0/XI36/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI7/MM5 N_XI0/XI36/XI7/NET34_XI0/XI36/XI7/MM5_d
+ N_XI0/XI36/XI7/NET33_XI0/XI36/XI7/MM5_g N_VDD_XI0/XI36/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI7/MM4 N_XI0/XI36/XI7/NET33_XI0/XI36/XI7/MM4_d
+ N_XI0/XI36/XI7/NET34_XI0/XI36/XI7/MM4_g N_VDD_XI0/XI36/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI7/MM10 N_XI0/XI36/XI7/NET35_XI0/XI36/XI7/MM10_d
+ N_XI0/XI36/XI7/NET36_XI0/XI36/XI7/MM10_g N_VDD_XI0/XI36/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI7/MM11 N_XI0/XI36/XI7/NET36_XI0/XI36/XI7/MM11_d
+ N_XI0/XI36/XI7/NET35_XI0/XI36/XI7/MM11_g N_VDD_XI0/XI36/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI8/MM2 N_XI0/XI36/XI8/NET34_XI0/XI36/XI8/MM2_d
+ N_XI0/XI36/XI8/NET33_XI0/XI36/XI8/MM2_g N_VSS_XI0/XI36/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM3 N_XI0/XI36/XI8/NET33_XI0/XI36/XI8/MM3_d
+ N_WL<68>_XI0/XI36/XI8/MM3_g N_BLN<7>_XI0/XI36/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM0 N_XI0/XI36/XI8/NET34_XI0/XI36/XI8/MM0_d
+ N_WL<68>_XI0/XI36/XI8/MM0_g N_BL<7>_XI0/XI36/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM1 N_XI0/XI36/XI8/NET33_XI0/XI36/XI8/MM1_d
+ N_XI0/XI36/XI8/NET34_XI0/XI36/XI8/MM1_g N_VSS_XI0/XI36/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM9 N_XI0/XI36/XI8/NET36_XI0/XI36/XI8/MM9_d
+ N_WL<69>_XI0/XI36/XI8/MM9_g N_BL<7>_XI0/XI36/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM6 N_XI0/XI36/XI8/NET35_XI0/XI36/XI8/MM6_d
+ N_XI0/XI36/XI8/NET36_XI0/XI36/XI8/MM6_g N_VSS_XI0/XI36/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM7 N_XI0/XI36/XI8/NET36_XI0/XI36/XI8/MM7_d
+ N_XI0/XI36/XI8/NET35_XI0/XI36/XI8/MM7_g N_VSS_XI0/XI36/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM8 N_XI0/XI36/XI8/NET35_XI0/XI36/XI8/MM8_d
+ N_WL<69>_XI0/XI36/XI8/MM8_g N_BLN<7>_XI0/XI36/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI8/MM5 N_XI0/XI36/XI8/NET34_XI0/XI36/XI8/MM5_d
+ N_XI0/XI36/XI8/NET33_XI0/XI36/XI8/MM5_g N_VDD_XI0/XI36/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI8/MM4 N_XI0/XI36/XI8/NET33_XI0/XI36/XI8/MM4_d
+ N_XI0/XI36/XI8/NET34_XI0/XI36/XI8/MM4_g N_VDD_XI0/XI36/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI8/MM10 N_XI0/XI36/XI8/NET35_XI0/XI36/XI8/MM10_d
+ N_XI0/XI36/XI8/NET36_XI0/XI36/XI8/MM10_g N_VDD_XI0/XI36/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI8/MM11 N_XI0/XI36/XI8/NET36_XI0/XI36/XI8/MM11_d
+ N_XI0/XI36/XI8/NET35_XI0/XI36/XI8/MM11_g N_VDD_XI0/XI36/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI9/MM2 N_XI0/XI36/XI9/NET34_XI0/XI36/XI9/MM2_d
+ N_XI0/XI36/XI9/NET33_XI0/XI36/XI9/MM2_g N_VSS_XI0/XI36/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM3 N_XI0/XI36/XI9/NET33_XI0/XI36/XI9/MM3_d
+ N_WL<68>_XI0/XI36/XI9/MM3_g N_BLN<6>_XI0/XI36/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM0 N_XI0/XI36/XI9/NET34_XI0/XI36/XI9/MM0_d
+ N_WL<68>_XI0/XI36/XI9/MM0_g N_BL<6>_XI0/XI36/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM1 N_XI0/XI36/XI9/NET33_XI0/XI36/XI9/MM1_d
+ N_XI0/XI36/XI9/NET34_XI0/XI36/XI9/MM1_g N_VSS_XI0/XI36/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM9 N_XI0/XI36/XI9/NET36_XI0/XI36/XI9/MM9_d
+ N_WL<69>_XI0/XI36/XI9/MM9_g N_BL<6>_XI0/XI36/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM6 N_XI0/XI36/XI9/NET35_XI0/XI36/XI9/MM6_d
+ N_XI0/XI36/XI9/NET36_XI0/XI36/XI9/MM6_g N_VSS_XI0/XI36/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM7 N_XI0/XI36/XI9/NET36_XI0/XI36/XI9/MM7_d
+ N_XI0/XI36/XI9/NET35_XI0/XI36/XI9/MM7_g N_VSS_XI0/XI36/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM8 N_XI0/XI36/XI9/NET35_XI0/XI36/XI9/MM8_d
+ N_WL<69>_XI0/XI36/XI9/MM8_g N_BLN<6>_XI0/XI36/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI9/MM5 N_XI0/XI36/XI9/NET34_XI0/XI36/XI9/MM5_d
+ N_XI0/XI36/XI9/NET33_XI0/XI36/XI9/MM5_g N_VDD_XI0/XI36/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI9/MM4 N_XI0/XI36/XI9/NET33_XI0/XI36/XI9/MM4_d
+ N_XI0/XI36/XI9/NET34_XI0/XI36/XI9/MM4_g N_VDD_XI0/XI36/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI9/MM10 N_XI0/XI36/XI9/NET35_XI0/XI36/XI9/MM10_d
+ N_XI0/XI36/XI9/NET36_XI0/XI36/XI9/MM10_g N_VDD_XI0/XI36/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI9/MM11 N_XI0/XI36/XI9/NET36_XI0/XI36/XI9/MM11_d
+ N_XI0/XI36/XI9/NET35_XI0/XI36/XI9/MM11_g N_VDD_XI0/XI36/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI10/MM2 N_XI0/XI36/XI10/NET34_XI0/XI36/XI10/MM2_d
+ N_XI0/XI36/XI10/NET33_XI0/XI36/XI10/MM2_g N_VSS_XI0/XI36/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM3 N_XI0/XI36/XI10/NET33_XI0/XI36/XI10/MM3_d
+ N_WL<68>_XI0/XI36/XI10/MM3_g N_BLN<5>_XI0/XI36/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM0 N_XI0/XI36/XI10/NET34_XI0/XI36/XI10/MM0_d
+ N_WL<68>_XI0/XI36/XI10/MM0_g N_BL<5>_XI0/XI36/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM1 N_XI0/XI36/XI10/NET33_XI0/XI36/XI10/MM1_d
+ N_XI0/XI36/XI10/NET34_XI0/XI36/XI10/MM1_g N_VSS_XI0/XI36/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM9 N_XI0/XI36/XI10/NET36_XI0/XI36/XI10/MM9_d
+ N_WL<69>_XI0/XI36/XI10/MM9_g N_BL<5>_XI0/XI36/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM6 N_XI0/XI36/XI10/NET35_XI0/XI36/XI10/MM6_d
+ N_XI0/XI36/XI10/NET36_XI0/XI36/XI10/MM6_g N_VSS_XI0/XI36/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM7 N_XI0/XI36/XI10/NET36_XI0/XI36/XI10/MM7_d
+ N_XI0/XI36/XI10/NET35_XI0/XI36/XI10/MM7_g N_VSS_XI0/XI36/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM8 N_XI0/XI36/XI10/NET35_XI0/XI36/XI10/MM8_d
+ N_WL<69>_XI0/XI36/XI10/MM8_g N_BLN<5>_XI0/XI36/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI10/MM5 N_XI0/XI36/XI10/NET34_XI0/XI36/XI10/MM5_d
+ N_XI0/XI36/XI10/NET33_XI0/XI36/XI10/MM5_g N_VDD_XI0/XI36/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI10/MM4 N_XI0/XI36/XI10/NET33_XI0/XI36/XI10/MM4_d
+ N_XI0/XI36/XI10/NET34_XI0/XI36/XI10/MM4_g N_VDD_XI0/XI36/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI10/MM10 N_XI0/XI36/XI10/NET35_XI0/XI36/XI10/MM10_d
+ N_XI0/XI36/XI10/NET36_XI0/XI36/XI10/MM10_g N_VDD_XI0/XI36/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI10/MM11 N_XI0/XI36/XI10/NET36_XI0/XI36/XI10/MM11_d
+ N_XI0/XI36/XI10/NET35_XI0/XI36/XI10/MM11_g N_VDD_XI0/XI36/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI11/MM2 N_XI0/XI36/XI11/NET34_XI0/XI36/XI11/MM2_d
+ N_XI0/XI36/XI11/NET33_XI0/XI36/XI11/MM2_g N_VSS_XI0/XI36/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM3 N_XI0/XI36/XI11/NET33_XI0/XI36/XI11/MM3_d
+ N_WL<68>_XI0/XI36/XI11/MM3_g N_BLN<4>_XI0/XI36/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM0 N_XI0/XI36/XI11/NET34_XI0/XI36/XI11/MM0_d
+ N_WL<68>_XI0/XI36/XI11/MM0_g N_BL<4>_XI0/XI36/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM1 N_XI0/XI36/XI11/NET33_XI0/XI36/XI11/MM1_d
+ N_XI0/XI36/XI11/NET34_XI0/XI36/XI11/MM1_g N_VSS_XI0/XI36/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM9 N_XI0/XI36/XI11/NET36_XI0/XI36/XI11/MM9_d
+ N_WL<69>_XI0/XI36/XI11/MM9_g N_BL<4>_XI0/XI36/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM6 N_XI0/XI36/XI11/NET35_XI0/XI36/XI11/MM6_d
+ N_XI0/XI36/XI11/NET36_XI0/XI36/XI11/MM6_g N_VSS_XI0/XI36/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM7 N_XI0/XI36/XI11/NET36_XI0/XI36/XI11/MM7_d
+ N_XI0/XI36/XI11/NET35_XI0/XI36/XI11/MM7_g N_VSS_XI0/XI36/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM8 N_XI0/XI36/XI11/NET35_XI0/XI36/XI11/MM8_d
+ N_WL<69>_XI0/XI36/XI11/MM8_g N_BLN<4>_XI0/XI36/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI11/MM5 N_XI0/XI36/XI11/NET34_XI0/XI36/XI11/MM5_d
+ N_XI0/XI36/XI11/NET33_XI0/XI36/XI11/MM5_g N_VDD_XI0/XI36/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI11/MM4 N_XI0/XI36/XI11/NET33_XI0/XI36/XI11/MM4_d
+ N_XI0/XI36/XI11/NET34_XI0/XI36/XI11/MM4_g N_VDD_XI0/XI36/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI11/MM10 N_XI0/XI36/XI11/NET35_XI0/XI36/XI11/MM10_d
+ N_XI0/XI36/XI11/NET36_XI0/XI36/XI11/MM10_g N_VDD_XI0/XI36/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI11/MM11 N_XI0/XI36/XI11/NET36_XI0/XI36/XI11/MM11_d
+ N_XI0/XI36/XI11/NET35_XI0/XI36/XI11/MM11_g N_VDD_XI0/XI36/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI12/MM2 N_XI0/XI36/XI12/NET34_XI0/XI36/XI12/MM2_d
+ N_XI0/XI36/XI12/NET33_XI0/XI36/XI12/MM2_g N_VSS_XI0/XI36/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM3 N_XI0/XI36/XI12/NET33_XI0/XI36/XI12/MM3_d
+ N_WL<68>_XI0/XI36/XI12/MM3_g N_BLN<3>_XI0/XI36/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM0 N_XI0/XI36/XI12/NET34_XI0/XI36/XI12/MM0_d
+ N_WL<68>_XI0/XI36/XI12/MM0_g N_BL<3>_XI0/XI36/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM1 N_XI0/XI36/XI12/NET33_XI0/XI36/XI12/MM1_d
+ N_XI0/XI36/XI12/NET34_XI0/XI36/XI12/MM1_g N_VSS_XI0/XI36/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM9 N_XI0/XI36/XI12/NET36_XI0/XI36/XI12/MM9_d
+ N_WL<69>_XI0/XI36/XI12/MM9_g N_BL<3>_XI0/XI36/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM6 N_XI0/XI36/XI12/NET35_XI0/XI36/XI12/MM6_d
+ N_XI0/XI36/XI12/NET36_XI0/XI36/XI12/MM6_g N_VSS_XI0/XI36/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM7 N_XI0/XI36/XI12/NET36_XI0/XI36/XI12/MM7_d
+ N_XI0/XI36/XI12/NET35_XI0/XI36/XI12/MM7_g N_VSS_XI0/XI36/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM8 N_XI0/XI36/XI12/NET35_XI0/XI36/XI12/MM8_d
+ N_WL<69>_XI0/XI36/XI12/MM8_g N_BLN<3>_XI0/XI36/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI12/MM5 N_XI0/XI36/XI12/NET34_XI0/XI36/XI12/MM5_d
+ N_XI0/XI36/XI12/NET33_XI0/XI36/XI12/MM5_g N_VDD_XI0/XI36/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI12/MM4 N_XI0/XI36/XI12/NET33_XI0/XI36/XI12/MM4_d
+ N_XI0/XI36/XI12/NET34_XI0/XI36/XI12/MM4_g N_VDD_XI0/XI36/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI12/MM10 N_XI0/XI36/XI12/NET35_XI0/XI36/XI12/MM10_d
+ N_XI0/XI36/XI12/NET36_XI0/XI36/XI12/MM10_g N_VDD_XI0/XI36/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI12/MM11 N_XI0/XI36/XI12/NET36_XI0/XI36/XI12/MM11_d
+ N_XI0/XI36/XI12/NET35_XI0/XI36/XI12/MM11_g N_VDD_XI0/XI36/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI13/MM2 N_XI0/XI36/XI13/NET34_XI0/XI36/XI13/MM2_d
+ N_XI0/XI36/XI13/NET33_XI0/XI36/XI13/MM2_g N_VSS_XI0/XI36/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM3 N_XI0/XI36/XI13/NET33_XI0/XI36/XI13/MM3_d
+ N_WL<68>_XI0/XI36/XI13/MM3_g N_BLN<2>_XI0/XI36/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM0 N_XI0/XI36/XI13/NET34_XI0/XI36/XI13/MM0_d
+ N_WL<68>_XI0/XI36/XI13/MM0_g N_BL<2>_XI0/XI36/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM1 N_XI0/XI36/XI13/NET33_XI0/XI36/XI13/MM1_d
+ N_XI0/XI36/XI13/NET34_XI0/XI36/XI13/MM1_g N_VSS_XI0/XI36/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM9 N_XI0/XI36/XI13/NET36_XI0/XI36/XI13/MM9_d
+ N_WL<69>_XI0/XI36/XI13/MM9_g N_BL<2>_XI0/XI36/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM6 N_XI0/XI36/XI13/NET35_XI0/XI36/XI13/MM6_d
+ N_XI0/XI36/XI13/NET36_XI0/XI36/XI13/MM6_g N_VSS_XI0/XI36/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM7 N_XI0/XI36/XI13/NET36_XI0/XI36/XI13/MM7_d
+ N_XI0/XI36/XI13/NET35_XI0/XI36/XI13/MM7_g N_VSS_XI0/XI36/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM8 N_XI0/XI36/XI13/NET35_XI0/XI36/XI13/MM8_d
+ N_WL<69>_XI0/XI36/XI13/MM8_g N_BLN<2>_XI0/XI36/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI13/MM5 N_XI0/XI36/XI13/NET34_XI0/XI36/XI13/MM5_d
+ N_XI0/XI36/XI13/NET33_XI0/XI36/XI13/MM5_g N_VDD_XI0/XI36/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI13/MM4 N_XI0/XI36/XI13/NET33_XI0/XI36/XI13/MM4_d
+ N_XI0/XI36/XI13/NET34_XI0/XI36/XI13/MM4_g N_VDD_XI0/XI36/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI13/MM10 N_XI0/XI36/XI13/NET35_XI0/XI36/XI13/MM10_d
+ N_XI0/XI36/XI13/NET36_XI0/XI36/XI13/MM10_g N_VDD_XI0/XI36/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI13/MM11 N_XI0/XI36/XI13/NET36_XI0/XI36/XI13/MM11_d
+ N_XI0/XI36/XI13/NET35_XI0/XI36/XI13/MM11_g N_VDD_XI0/XI36/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI14/MM2 N_XI0/XI36/XI14/NET34_XI0/XI36/XI14/MM2_d
+ N_XI0/XI36/XI14/NET33_XI0/XI36/XI14/MM2_g N_VSS_XI0/XI36/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM3 N_XI0/XI36/XI14/NET33_XI0/XI36/XI14/MM3_d
+ N_WL<68>_XI0/XI36/XI14/MM3_g N_BLN<1>_XI0/XI36/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM0 N_XI0/XI36/XI14/NET34_XI0/XI36/XI14/MM0_d
+ N_WL<68>_XI0/XI36/XI14/MM0_g N_BL<1>_XI0/XI36/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM1 N_XI0/XI36/XI14/NET33_XI0/XI36/XI14/MM1_d
+ N_XI0/XI36/XI14/NET34_XI0/XI36/XI14/MM1_g N_VSS_XI0/XI36/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM9 N_XI0/XI36/XI14/NET36_XI0/XI36/XI14/MM9_d
+ N_WL<69>_XI0/XI36/XI14/MM9_g N_BL<1>_XI0/XI36/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM6 N_XI0/XI36/XI14/NET35_XI0/XI36/XI14/MM6_d
+ N_XI0/XI36/XI14/NET36_XI0/XI36/XI14/MM6_g N_VSS_XI0/XI36/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM7 N_XI0/XI36/XI14/NET36_XI0/XI36/XI14/MM7_d
+ N_XI0/XI36/XI14/NET35_XI0/XI36/XI14/MM7_g N_VSS_XI0/XI36/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM8 N_XI0/XI36/XI14/NET35_XI0/XI36/XI14/MM8_d
+ N_WL<69>_XI0/XI36/XI14/MM8_g N_BLN<1>_XI0/XI36/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI14/MM5 N_XI0/XI36/XI14/NET34_XI0/XI36/XI14/MM5_d
+ N_XI0/XI36/XI14/NET33_XI0/XI36/XI14/MM5_g N_VDD_XI0/XI36/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI14/MM4 N_XI0/XI36/XI14/NET33_XI0/XI36/XI14/MM4_d
+ N_XI0/XI36/XI14/NET34_XI0/XI36/XI14/MM4_g N_VDD_XI0/XI36/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI14/MM10 N_XI0/XI36/XI14/NET35_XI0/XI36/XI14/MM10_d
+ N_XI0/XI36/XI14/NET36_XI0/XI36/XI14/MM10_g N_VDD_XI0/XI36/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI14/MM11 N_XI0/XI36/XI14/NET36_XI0/XI36/XI14/MM11_d
+ N_XI0/XI36/XI14/NET35_XI0/XI36/XI14/MM11_g N_VDD_XI0/XI36/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI15/MM2 N_XI0/XI36/XI15/NET34_XI0/XI36/XI15/MM2_d
+ N_XI0/XI36/XI15/NET33_XI0/XI36/XI15/MM2_g N_VSS_XI0/XI36/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM3 N_XI0/XI36/XI15/NET33_XI0/XI36/XI15/MM3_d
+ N_WL<68>_XI0/XI36/XI15/MM3_g N_BLN<0>_XI0/XI36/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM0 N_XI0/XI36/XI15/NET34_XI0/XI36/XI15/MM0_d
+ N_WL<68>_XI0/XI36/XI15/MM0_g N_BL<0>_XI0/XI36/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM1 N_XI0/XI36/XI15/NET33_XI0/XI36/XI15/MM1_d
+ N_XI0/XI36/XI15/NET34_XI0/XI36/XI15/MM1_g N_VSS_XI0/XI36/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM9 N_XI0/XI36/XI15/NET36_XI0/XI36/XI15/MM9_d
+ N_WL<69>_XI0/XI36/XI15/MM9_g N_BL<0>_XI0/XI36/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM6 N_XI0/XI36/XI15/NET35_XI0/XI36/XI15/MM6_d
+ N_XI0/XI36/XI15/NET36_XI0/XI36/XI15/MM6_g N_VSS_XI0/XI36/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM7 N_XI0/XI36/XI15/NET36_XI0/XI36/XI15/MM7_d
+ N_XI0/XI36/XI15/NET35_XI0/XI36/XI15/MM7_g N_VSS_XI0/XI36/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM8 N_XI0/XI36/XI15/NET35_XI0/XI36/XI15/MM8_d
+ N_WL<69>_XI0/XI36/XI15/MM8_g N_BLN<0>_XI0/XI36/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI36/XI15/MM5 N_XI0/XI36/XI15/NET34_XI0/XI36/XI15/MM5_d
+ N_XI0/XI36/XI15/NET33_XI0/XI36/XI15/MM5_g N_VDD_XI0/XI36/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI15/MM4 N_XI0/XI36/XI15/NET33_XI0/XI36/XI15/MM4_d
+ N_XI0/XI36/XI15/NET34_XI0/XI36/XI15/MM4_g N_VDD_XI0/XI36/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI15/MM10 N_XI0/XI36/XI15/NET35_XI0/XI36/XI15/MM10_d
+ N_XI0/XI36/XI15/NET36_XI0/XI36/XI15/MM10_g N_VDD_XI0/XI36/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI36/XI15/MM11 N_XI0/XI36/XI15/NET36_XI0/XI36/XI15/MM11_d
+ N_XI0/XI36/XI15/NET35_XI0/XI36/XI15/MM11_g N_VDD_XI0/XI36/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI0/MM2 N_XI0/XI37/XI0/NET34_XI0/XI37/XI0/MM2_d
+ N_XI0/XI37/XI0/NET33_XI0/XI37/XI0/MM2_g N_VSS_XI0/XI37/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM3 N_XI0/XI37/XI0/NET33_XI0/XI37/XI0/MM3_d
+ N_WL<70>_XI0/XI37/XI0/MM3_g N_BLN<15>_XI0/XI37/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM0 N_XI0/XI37/XI0/NET34_XI0/XI37/XI0/MM0_d
+ N_WL<70>_XI0/XI37/XI0/MM0_g N_BL<15>_XI0/XI37/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM1 N_XI0/XI37/XI0/NET33_XI0/XI37/XI0/MM1_d
+ N_XI0/XI37/XI0/NET34_XI0/XI37/XI0/MM1_g N_VSS_XI0/XI37/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM9 N_XI0/XI37/XI0/NET36_XI0/XI37/XI0/MM9_d
+ N_WL<71>_XI0/XI37/XI0/MM9_g N_BL<15>_XI0/XI37/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM6 N_XI0/XI37/XI0/NET35_XI0/XI37/XI0/MM6_d
+ N_XI0/XI37/XI0/NET36_XI0/XI37/XI0/MM6_g N_VSS_XI0/XI37/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM7 N_XI0/XI37/XI0/NET36_XI0/XI37/XI0/MM7_d
+ N_XI0/XI37/XI0/NET35_XI0/XI37/XI0/MM7_g N_VSS_XI0/XI37/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM8 N_XI0/XI37/XI0/NET35_XI0/XI37/XI0/MM8_d
+ N_WL<71>_XI0/XI37/XI0/MM8_g N_BLN<15>_XI0/XI37/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI0/MM5 N_XI0/XI37/XI0/NET34_XI0/XI37/XI0/MM5_d
+ N_XI0/XI37/XI0/NET33_XI0/XI37/XI0/MM5_g N_VDD_XI0/XI37/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI0/MM4 N_XI0/XI37/XI0/NET33_XI0/XI37/XI0/MM4_d
+ N_XI0/XI37/XI0/NET34_XI0/XI37/XI0/MM4_g N_VDD_XI0/XI37/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI0/MM10 N_XI0/XI37/XI0/NET35_XI0/XI37/XI0/MM10_d
+ N_XI0/XI37/XI0/NET36_XI0/XI37/XI0/MM10_g N_VDD_XI0/XI37/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI0/MM11 N_XI0/XI37/XI0/NET36_XI0/XI37/XI0/MM11_d
+ N_XI0/XI37/XI0/NET35_XI0/XI37/XI0/MM11_g N_VDD_XI0/XI37/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI1/MM2 N_XI0/XI37/XI1/NET34_XI0/XI37/XI1/MM2_d
+ N_XI0/XI37/XI1/NET33_XI0/XI37/XI1/MM2_g N_VSS_XI0/XI37/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM3 N_XI0/XI37/XI1/NET33_XI0/XI37/XI1/MM3_d
+ N_WL<70>_XI0/XI37/XI1/MM3_g N_BLN<14>_XI0/XI37/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM0 N_XI0/XI37/XI1/NET34_XI0/XI37/XI1/MM0_d
+ N_WL<70>_XI0/XI37/XI1/MM0_g N_BL<14>_XI0/XI37/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM1 N_XI0/XI37/XI1/NET33_XI0/XI37/XI1/MM1_d
+ N_XI0/XI37/XI1/NET34_XI0/XI37/XI1/MM1_g N_VSS_XI0/XI37/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM9 N_XI0/XI37/XI1/NET36_XI0/XI37/XI1/MM9_d
+ N_WL<71>_XI0/XI37/XI1/MM9_g N_BL<14>_XI0/XI37/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM6 N_XI0/XI37/XI1/NET35_XI0/XI37/XI1/MM6_d
+ N_XI0/XI37/XI1/NET36_XI0/XI37/XI1/MM6_g N_VSS_XI0/XI37/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM7 N_XI0/XI37/XI1/NET36_XI0/XI37/XI1/MM7_d
+ N_XI0/XI37/XI1/NET35_XI0/XI37/XI1/MM7_g N_VSS_XI0/XI37/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM8 N_XI0/XI37/XI1/NET35_XI0/XI37/XI1/MM8_d
+ N_WL<71>_XI0/XI37/XI1/MM8_g N_BLN<14>_XI0/XI37/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI1/MM5 N_XI0/XI37/XI1/NET34_XI0/XI37/XI1/MM5_d
+ N_XI0/XI37/XI1/NET33_XI0/XI37/XI1/MM5_g N_VDD_XI0/XI37/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI1/MM4 N_XI0/XI37/XI1/NET33_XI0/XI37/XI1/MM4_d
+ N_XI0/XI37/XI1/NET34_XI0/XI37/XI1/MM4_g N_VDD_XI0/XI37/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI1/MM10 N_XI0/XI37/XI1/NET35_XI0/XI37/XI1/MM10_d
+ N_XI0/XI37/XI1/NET36_XI0/XI37/XI1/MM10_g N_VDD_XI0/XI37/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI1/MM11 N_XI0/XI37/XI1/NET36_XI0/XI37/XI1/MM11_d
+ N_XI0/XI37/XI1/NET35_XI0/XI37/XI1/MM11_g N_VDD_XI0/XI37/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI2/MM2 N_XI0/XI37/XI2/NET34_XI0/XI37/XI2/MM2_d
+ N_XI0/XI37/XI2/NET33_XI0/XI37/XI2/MM2_g N_VSS_XI0/XI37/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM3 N_XI0/XI37/XI2/NET33_XI0/XI37/XI2/MM3_d
+ N_WL<70>_XI0/XI37/XI2/MM3_g N_BLN<13>_XI0/XI37/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM0 N_XI0/XI37/XI2/NET34_XI0/XI37/XI2/MM0_d
+ N_WL<70>_XI0/XI37/XI2/MM0_g N_BL<13>_XI0/XI37/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM1 N_XI0/XI37/XI2/NET33_XI0/XI37/XI2/MM1_d
+ N_XI0/XI37/XI2/NET34_XI0/XI37/XI2/MM1_g N_VSS_XI0/XI37/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM9 N_XI0/XI37/XI2/NET36_XI0/XI37/XI2/MM9_d
+ N_WL<71>_XI0/XI37/XI2/MM9_g N_BL<13>_XI0/XI37/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM6 N_XI0/XI37/XI2/NET35_XI0/XI37/XI2/MM6_d
+ N_XI0/XI37/XI2/NET36_XI0/XI37/XI2/MM6_g N_VSS_XI0/XI37/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM7 N_XI0/XI37/XI2/NET36_XI0/XI37/XI2/MM7_d
+ N_XI0/XI37/XI2/NET35_XI0/XI37/XI2/MM7_g N_VSS_XI0/XI37/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM8 N_XI0/XI37/XI2/NET35_XI0/XI37/XI2/MM8_d
+ N_WL<71>_XI0/XI37/XI2/MM8_g N_BLN<13>_XI0/XI37/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI2/MM5 N_XI0/XI37/XI2/NET34_XI0/XI37/XI2/MM5_d
+ N_XI0/XI37/XI2/NET33_XI0/XI37/XI2/MM5_g N_VDD_XI0/XI37/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI2/MM4 N_XI0/XI37/XI2/NET33_XI0/XI37/XI2/MM4_d
+ N_XI0/XI37/XI2/NET34_XI0/XI37/XI2/MM4_g N_VDD_XI0/XI37/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI2/MM10 N_XI0/XI37/XI2/NET35_XI0/XI37/XI2/MM10_d
+ N_XI0/XI37/XI2/NET36_XI0/XI37/XI2/MM10_g N_VDD_XI0/XI37/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI2/MM11 N_XI0/XI37/XI2/NET36_XI0/XI37/XI2/MM11_d
+ N_XI0/XI37/XI2/NET35_XI0/XI37/XI2/MM11_g N_VDD_XI0/XI37/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI3/MM2 N_XI0/XI37/XI3/NET34_XI0/XI37/XI3/MM2_d
+ N_XI0/XI37/XI3/NET33_XI0/XI37/XI3/MM2_g N_VSS_XI0/XI37/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM3 N_XI0/XI37/XI3/NET33_XI0/XI37/XI3/MM3_d
+ N_WL<70>_XI0/XI37/XI3/MM3_g N_BLN<12>_XI0/XI37/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM0 N_XI0/XI37/XI3/NET34_XI0/XI37/XI3/MM0_d
+ N_WL<70>_XI0/XI37/XI3/MM0_g N_BL<12>_XI0/XI37/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM1 N_XI0/XI37/XI3/NET33_XI0/XI37/XI3/MM1_d
+ N_XI0/XI37/XI3/NET34_XI0/XI37/XI3/MM1_g N_VSS_XI0/XI37/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM9 N_XI0/XI37/XI3/NET36_XI0/XI37/XI3/MM9_d
+ N_WL<71>_XI0/XI37/XI3/MM9_g N_BL<12>_XI0/XI37/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM6 N_XI0/XI37/XI3/NET35_XI0/XI37/XI3/MM6_d
+ N_XI0/XI37/XI3/NET36_XI0/XI37/XI3/MM6_g N_VSS_XI0/XI37/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM7 N_XI0/XI37/XI3/NET36_XI0/XI37/XI3/MM7_d
+ N_XI0/XI37/XI3/NET35_XI0/XI37/XI3/MM7_g N_VSS_XI0/XI37/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM8 N_XI0/XI37/XI3/NET35_XI0/XI37/XI3/MM8_d
+ N_WL<71>_XI0/XI37/XI3/MM8_g N_BLN<12>_XI0/XI37/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI3/MM5 N_XI0/XI37/XI3/NET34_XI0/XI37/XI3/MM5_d
+ N_XI0/XI37/XI3/NET33_XI0/XI37/XI3/MM5_g N_VDD_XI0/XI37/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI3/MM4 N_XI0/XI37/XI3/NET33_XI0/XI37/XI3/MM4_d
+ N_XI0/XI37/XI3/NET34_XI0/XI37/XI3/MM4_g N_VDD_XI0/XI37/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI3/MM10 N_XI0/XI37/XI3/NET35_XI0/XI37/XI3/MM10_d
+ N_XI0/XI37/XI3/NET36_XI0/XI37/XI3/MM10_g N_VDD_XI0/XI37/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI3/MM11 N_XI0/XI37/XI3/NET36_XI0/XI37/XI3/MM11_d
+ N_XI0/XI37/XI3/NET35_XI0/XI37/XI3/MM11_g N_VDD_XI0/XI37/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI4/MM2 N_XI0/XI37/XI4/NET34_XI0/XI37/XI4/MM2_d
+ N_XI0/XI37/XI4/NET33_XI0/XI37/XI4/MM2_g N_VSS_XI0/XI37/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM3 N_XI0/XI37/XI4/NET33_XI0/XI37/XI4/MM3_d
+ N_WL<70>_XI0/XI37/XI4/MM3_g N_BLN<11>_XI0/XI37/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM0 N_XI0/XI37/XI4/NET34_XI0/XI37/XI4/MM0_d
+ N_WL<70>_XI0/XI37/XI4/MM0_g N_BL<11>_XI0/XI37/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM1 N_XI0/XI37/XI4/NET33_XI0/XI37/XI4/MM1_d
+ N_XI0/XI37/XI4/NET34_XI0/XI37/XI4/MM1_g N_VSS_XI0/XI37/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM9 N_XI0/XI37/XI4/NET36_XI0/XI37/XI4/MM9_d
+ N_WL<71>_XI0/XI37/XI4/MM9_g N_BL<11>_XI0/XI37/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM6 N_XI0/XI37/XI4/NET35_XI0/XI37/XI4/MM6_d
+ N_XI0/XI37/XI4/NET36_XI0/XI37/XI4/MM6_g N_VSS_XI0/XI37/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM7 N_XI0/XI37/XI4/NET36_XI0/XI37/XI4/MM7_d
+ N_XI0/XI37/XI4/NET35_XI0/XI37/XI4/MM7_g N_VSS_XI0/XI37/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM8 N_XI0/XI37/XI4/NET35_XI0/XI37/XI4/MM8_d
+ N_WL<71>_XI0/XI37/XI4/MM8_g N_BLN<11>_XI0/XI37/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI4/MM5 N_XI0/XI37/XI4/NET34_XI0/XI37/XI4/MM5_d
+ N_XI0/XI37/XI4/NET33_XI0/XI37/XI4/MM5_g N_VDD_XI0/XI37/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI4/MM4 N_XI0/XI37/XI4/NET33_XI0/XI37/XI4/MM4_d
+ N_XI0/XI37/XI4/NET34_XI0/XI37/XI4/MM4_g N_VDD_XI0/XI37/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI4/MM10 N_XI0/XI37/XI4/NET35_XI0/XI37/XI4/MM10_d
+ N_XI0/XI37/XI4/NET36_XI0/XI37/XI4/MM10_g N_VDD_XI0/XI37/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI4/MM11 N_XI0/XI37/XI4/NET36_XI0/XI37/XI4/MM11_d
+ N_XI0/XI37/XI4/NET35_XI0/XI37/XI4/MM11_g N_VDD_XI0/XI37/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI5/MM2 N_XI0/XI37/XI5/NET34_XI0/XI37/XI5/MM2_d
+ N_XI0/XI37/XI5/NET33_XI0/XI37/XI5/MM2_g N_VSS_XI0/XI37/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM3 N_XI0/XI37/XI5/NET33_XI0/XI37/XI5/MM3_d
+ N_WL<70>_XI0/XI37/XI5/MM3_g N_BLN<10>_XI0/XI37/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM0 N_XI0/XI37/XI5/NET34_XI0/XI37/XI5/MM0_d
+ N_WL<70>_XI0/XI37/XI5/MM0_g N_BL<10>_XI0/XI37/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM1 N_XI0/XI37/XI5/NET33_XI0/XI37/XI5/MM1_d
+ N_XI0/XI37/XI5/NET34_XI0/XI37/XI5/MM1_g N_VSS_XI0/XI37/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM9 N_XI0/XI37/XI5/NET36_XI0/XI37/XI5/MM9_d
+ N_WL<71>_XI0/XI37/XI5/MM9_g N_BL<10>_XI0/XI37/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM6 N_XI0/XI37/XI5/NET35_XI0/XI37/XI5/MM6_d
+ N_XI0/XI37/XI5/NET36_XI0/XI37/XI5/MM6_g N_VSS_XI0/XI37/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM7 N_XI0/XI37/XI5/NET36_XI0/XI37/XI5/MM7_d
+ N_XI0/XI37/XI5/NET35_XI0/XI37/XI5/MM7_g N_VSS_XI0/XI37/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM8 N_XI0/XI37/XI5/NET35_XI0/XI37/XI5/MM8_d
+ N_WL<71>_XI0/XI37/XI5/MM8_g N_BLN<10>_XI0/XI37/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI5/MM5 N_XI0/XI37/XI5/NET34_XI0/XI37/XI5/MM5_d
+ N_XI0/XI37/XI5/NET33_XI0/XI37/XI5/MM5_g N_VDD_XI0/XI37/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI5/MM4 N_XI0/XI37/XI5/NET33_XI0/XI37/XI5/MM4_d
+ N_XI0/XI37/XI5/NET34_XI0/XI37/XI5/MM4_g N_VDD_XI0/XI37/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI5/MM10 N_XI0/XI37/XI5/NET35_XI0/XI37/XI5/MM10_d
+ N_XI0/XI37/XI5/NET36_XI0/XI37/XI5/MM10_g N_VDD_XI0/XI37/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI5/MM11 N_XI0/XI37/XI5/NET36_XI0/XI37/XI5/MM11_d
+ N_XI0/XI37/XI5/NET35_XI0/XI37/XI5/MM11_g N_VDD_XI0/XI37/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI6/MM2 N_XI0/XI37/XI6/NET34_XI0/XI37/XI6/MM2_d
+ N_XI0/XI37/XI6/NET33_XI0/XI37/XI6/MM2_g N_VSS_XI0/XI37/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM3 N_XI0/XI37/XI6/NET33_XI0/XI37/XI6/MM3_d
+ N_WL<70>_XI0/XI37/XI6/MM3_g N_BLN<9>_XI0/XI37/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM0 N_XI0/XI37/XI6/NET34_XI0/XI37/XI6/MM0_d
+ N_WL<70>_XI0/XI37/XI6/MM0_g N_BL<9>_XI0/XI37/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM1 N_XI0/XI37/XI6/NET33_XI0/XI37/XI6/MM1_d
+ N_XI0/XI37/XI6/NET34_XI0/XI37/XI6/MM1_g N_VSS_XI0/XI37/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM9 N_XI0/XI37/XI6/NET36_XI0/XI37/XI6/MM9_d
+ N_WL<71>_XI0/XI37/XI6/MM9_g N_BL<9>_XI0/XI37/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM6 N_XI0/XI37/XI6/NET35_XI0/XI37/XI6/MM6_d
+ N_XI0/XI37/XI6/NET36_XI0/XI37/XI6/MM6_g N_VSS_XI0/XI37/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM7 N_XI0/XI37/XI6/NET36_XI0/XI37/XI6/MM7_d
+ N_XI0/XI37/XI6/NET35_XI0/XI37/XI6/MM7_g N_VSS_XI0/XI37/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM8 N_XI0/XI37/XI6/NET35_XI0/XI37/XI6/MM8_d
+ N_WL<71>_XI0/XI37/XI6/MM8_g N_BLN<9>_XI0/XI37/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI6/MM5 N_XI0/XI37/XI6/NET34_XI0/XI37/XI6/MM5_d
+ N_XI0/XI37/XI6/NET33_XI0/XI37/XI6/MM5_g N_VDD_XI0/XI37/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI6/MM4 N_XI0/XI37/XI6/NET33_XI0/XI37/XI6/MM4_d
+ N_XI0/XI37/XI6/NET34_XI0/XI37/XI6/MM4_g N_VDD_XI0/XI37/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI6/MM10 N_XI0/XI37/XI6/NET35_XI0/XI37/XI6/MM10_d
+ N_XI0/XI37/XI6/NET36_XI0/XI37/XI6/MM10_g N_VDD_XI0/XI37/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI6/MM11 N_XI0/XI37/XI6/NET36_XI0/XI37/XI6/MM11_d
+ N_XI0/XI37/XI6/NET35_XI0/XI37/XI6/MM11_g N_VDD_XI0/XI37/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI7/MM2 N_XI0/XI37/XI7/NET34_XI0/XI37/XI7/MM2_d
+ N_XI0/XI37/XI7/NET33_XI0/XI37/XI7/MM2_g N_VSS_XI0/XI37/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM3 N_XI0/XI37/XI7/NET33_XI0/XI37/XI7/MM3_d
+ N_WL<70>_XI0/XI37/XI7/MM3_g N_BLN<8>_XI0/XI37/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM0 N_XI0/XI37/XI7/NET34_XI0/XI37/XI7/MM0_d
+ N_WL<70>_XI0/XI37/XI7/MM0_g N_BL<8>_XI0/XI37/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM1 N_XI0/XI37/XI7/NET33_XI0/XI37/XI7/MM1_d
+ N_XI0/XI37/XI7/NET34_XI0/XI37/XI7/MM1_g N_VSS_XI0/XI37/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM9 N_XI0/XI37/XI7/NET36_XI0/XI37/XI7/MM9_d
+ N_WL<71>_XI0/XI37/XI7/MM9_g N_BL<8>_XI0/XI37/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM6 N_XI0/XI37/XI7/NET35_XI0/XI37/XI7/MM6_d
+ N_XI0/XI37/XI7/NET36_XI0/XI37/XI7/MM6_g N_VSS_XI0/XI37/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM7 N_XI0/XI37/XI7/NET36_XI0/XI37/XI7/MM7_d
+ N_XI0/XI37/XI7/NET35_XI0/XI37/XI7/MM7_g N_VSS_XI0/XI37/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM8 N_XI0/XI37/XI7/NET35_XI0/XI37/XI7/MM8_d
+ N_WL<71>_XI0/XI37/XI7/MM8_g N_BLN<8>_XI0/XI37/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI7/MM5 N_XI0/XI37/XI7/NET34_XI0/XI37/XI7/MM5_d
+ N_XI0/XI37/XI7/NET33_XI0/XI37/XI7/MM5_g N_VDD_XI0/XI37/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI7/MM4 N_XI0/XI37/XI7/NET33_XI0/XI37/XI7/MM4_d
+ N_XI0/XI37/XI7/NET34_XI0/XI37/XI7/MM4_g N_VDD_XI0/XI37/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI7/MM10 N_XI0/XI37/XI7/NET35_XI0/XI37/XI7/MM10_d
+ N_XI0/XI37/XI7/NET36_XI0/XI37/XI7/MM10_g N_VDD_XI0/XI37/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI7/MM11 N_XI0/XI37/XI7/NET36_XI0/XI37/XI7/MM11_d
+ N_XI0/XI37/XI7/NET35_XI0/XI37/XI7/MM11_g N_VDD_XI0/XI37/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI8/MM2 N_XI0/XI37/XI8/NET34_XI0/XI37/XI8/MM2_d
+ N_XI0/XI37/XI8/NET33_XI0/XI37/XI8/MM2_g N_VSS_XI0/XI37/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM3 N_XI0/XI37/XI8/NET33_XI0/XI37/XI8/MM3_d
+ N_WL<70>_XI0/XI37/XI8/MM3_g N_BLN<7>_XI0/XI37/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM0 N_XI0/XI37/XI8/NET34_XI0/XI37/XI8/MM0_d
+ N_WL<70>_XI0/XI37/XI8/MM0_g N_BL<7>_XI0/XI37/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM1 N_XI0/XI37/XI8/NET33_XI0/XI37/XI8/MM1_d
+ N_XI0/XI37/XI8/NET34_XI0/XI37/XI8/MM1_g N_VSS_XI0/XI37/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM9 N_XI0/XI37/XI8/NET36_XI0/XI37/XI8/MM9_d
+ N_WL<71>_XI0/XI37/XI8/MM9_g N_BL<7>_XI0/XI37/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM6 N_XI0/XI37/XI8/NET35_XI0/XI37/XI8/MM6_d
+ N_XI0/XI37/XI8/NET36_XI0/XI37/XI8/MM6_g N_VSS_XI0/XI37/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM7 N_XI0/XI37/XI8/NET36_XI0/XI37/XI8/MM7_d
+ N_XI0/XI37/XI8/NET35_XI0/XI37/XI8/MM7_g N_VSS_XI0/XI37/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM8 N_XI0/XI37/XI8/NET35_XI0/XI37/XI8/MM8_d
+ N_WL<71>_XI0/XI37/XI8/MM8_g N_BLN<7>_XI0/XI37/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI8/MM5 N_XI0/XI37/XI8/NET34_XI0/XI37/XI8/MM5_d
+ N_XI0/XI37/XI8/NET33_XI0/XI37/XI8/MM5_g N_VDD_XI0/XI37/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI8/MM4 N_XI0/XI37/XI8/NET33_XI0/XI37/XI8/MM4_d
+ N_XI0/XI37/XI8/NET34_XI0/XI37/XI8/MM4_g N_VDD_XI0/XI37/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI8/MM10 N_XI0/XI37/XI8/NET35_XI0/XI37/XI8/MM10_d
+ N_XI0/XI37/XI8/NET36_XI0/XI37/XI8/MM10_g N_VDD_XI0/XI37/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI8/MM11 N_XI0/XI37/XI8/NET36_XI0/XI37/XI8/MM11_d
+ N_XI0/XI37/XI8/NET35_XI0/XI37/XI8/MM11_g N_VDD_XI0/XI37/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI9/MM2 N_XI0/XI37/XI9/NET34_XI0/XI37/XI9/MM2_d
+ N_XI0/XI37/XI9/NET33_XI0/XI37/XI9/MM2_g N_VSS_XI0/XI37/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM3 N_XI0/XI37/XI9/NET33_XI0/XI37/XI9/MM3_d
+ N_WL<70>_XI0/XI37/XI9/MM3_g N_BLN<6>_XI0/XI37/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM0 N_XI0/XI37/XI9/NET34_XI0/XI37/XI9/MM0_d
+ N_WL<70>_XI0/XI37/XI9/MM0_g N_BL<6>_XI0/XI37/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM1 N_XI0/XI37/XI9/NET33_XI0/XI37/XI9/MM1_d
+ N_XI0/XI37/XI9/NET34_XI0/XI37/XI9/MM1_g N_VSS_XI0/XI37/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM9 N_XI0/XI37/XI9/NET36_XI0/XI37/XI9/MM9_d
+ N_WL<71>_XI0/XI37/XI9/MM9_g N_BL<6>_XI0/XI37/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM6 N_XI0/XI37/XI9/NET35_XI0/XI37/XI9/MM6_d
+ N_XI0/XI37/XI9/NET36_XI0/XI37/XI9/MM6_g N_VSS_XI0/XI37/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM7 N_XI0/XI37/XI9/NET36_XI0/XI37/XI9/MM7_d
+ N_XI0/XI37/XI9/NET35_XI0/XI37/XI9/MM7_g N_VSS_XI0/XI37/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM8 N_XI0/XI37/XI9/NET35_XI0/XI37/XI9/MM8_d
+ N_WL<71>_XI0/XI37/XI9/MM8_g N_BLN<6>_XI0/XI37/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI9/MM5 N_XI0/XI37/XI9/NET34_XI0/XI37/XI9/MM5_d
+ N_XI0/XI37/XI9/NET33_XI0/XI37/XI9/MM5_g N_VDD_XI0/XI37/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI9/MM4 N_XI0/XI37/XI9/NET33_XI0/XI37/XI9/MM4_d
+ N_XI0/XI37/XI9/NET34_XI0/XI37/XI9/MM4_g N_VDD_XI0/XI37/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI9/MM10 N_XI0/XI37/XI9/NET35_XI0/XI37/XI9/MM10_d
+ N_XI0/XI37/XI9/NET36_XI0/XI37/XI9/MM10_g N_VDD_XI0/XI37/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI9/MM11 N_XI0/XI37/XI9/NET36_XI0/XI37/XI9/MM11_d
+ N_XI0/XI37/XI9/NET35_XI0/XI37/XI9/MM11_g N_VDD_XI0/XI37/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI10/MM2 N_XI0/XI37/XI10/NET34_XI0/XI37/XI10/MM2_d
+ N_XI0/XI37/XI10/NET33_XI0/XI37/XI10/MM2_g N_VSS_XI0/XI37/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM3 N_XI0/XI37/XI10/NET33_XI0/XI37/XI10/MM3_d
+ N_WL<70>_XI0/XI37/XI10/MM3_g N_BLN<5>_XI0/XI37/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM0 N_XI0/XI37/XI10/NET34_XI0/XI37/XI10/MM0_d
+ N_WL<70>_XI0/XI37/XI10/MM0_g N_BL<5>_XI0/XI37/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM1 N_XI0/XI37/XI10/NET33_XI0/XI37/XI10/MM1_d
+ N_XI0/XI37/XI10/NET34_XI0/XI37/XI10/MM1_g N_VSS_XI0/XI37/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM9 N_XI0/XI37/XI10/NET36_XI0/XI37/XI10/MM9_d
+ N_WL<71>_XI0/XI37/XI10/MM9_g N_BL<5>_XI0/XI37/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM6 N_XI0/XI37/XI10/NET35_XI0/XI37/XI10/MM6_d
+ N_XI0/XI37/XI10/NET36_XI0/XI37/XI10/MM6_g N_VSS_XI0/XI37/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM7 N_XI0/XI37/XI10/NET36_XI0/XI37/XI10/MM7_d
+ N_XI0/XI37/XI10/NET35_XI0/XI37/XI10/MM7_g N_VSS_XI0/XI37/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM8 N_XI0/XI37/XI10/NET35_XI0/XI37/XI10/MM8_d
+ N_WL<71>_XI0/XI37/XI10/MM8_g N_BLN<5>_XI0/XI37/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI10/MM5 N_XI0/XI37/XI10/NET34_XI0/XI37/XI10/MM5_d
+ N_XI0/XI37/XI10/NET33_XI0/XI37/XI10/MM5_g N_VDD_XI0/XI37/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI10/MM4 N_XI0/XI37/XI10/NET33_XI0/XI37/XI10/MM4_d
+ N_XI0/XI37/XI10/NET34_XI0/XI37/XI10/MM4_g N_VDD_XI0/XI37/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI10/MM10 N_XI0/XI37/XI10/NET35_XI0/XI37/XI10/MM10_d
+ N_XI0/XI37/XI10/NET36_XI0/XI37/XI10/MM10_g N_VDD_XI0/XI37/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI10/MM11 N_XI0/XI37/XI10/NET36_XI0/XI37/XI10/MM11_d
+ N_XI0/XI37/XI10/NET35_XI0/XI37/XI10/MM11_g N_VDD_XI0/XI37/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI11/MM2 N_XI0/XI37/XI11/NET34_XI0/XI37/XI11/MM2_d
+ N_XI0/XI37/XI11/NET33_XI0/XI37/XI11/MM2_g N_VSS_XI0/XI37/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM3 N_XI0/XI37/XI11/NET33_XI0/XI37/XI11/MM3_d
+ N_WL<70>_XI0/XI37/XI11/MM3_g N_BLN<4>_XI0/XI37/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM0 N_XI0/XI37/XI11/NET34_XI0/XI37/XI11/MM0_d
+ N_WL<70>_XI0/XI37/XI11/MM0_g N_BL<4>_XI0/XI37/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM1 N_XI0/XI37/XI11/NET33_XI0/XI37/XI11/MM1_d
+ N_XI0/XI37/XI11/NET34_XI0/XI37/XI11/MM1_g N_VSS_XI0/XI37/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM9 N_XI0/XI37/XI11/NET36_XI0/XI37/XI11/MM9_d
+ N_WL<71>_XI0/XI37/XI11/MM9_g N_BL<4>_XI0/XI37/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM6 N_XI0/XI37/XI11/NET35_XI0/XI37/XI11/MM6_d
+ N_XI0/XI37/XI11/NET36_XI0/XI37/XI11/MM6_g N_VSS_XI0/XI37/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM7 N_XI0/XI37/XI11/NET36_XI0/XI37/XI11/MM7_d
+ N_XI0/XI37/XI11/NET35_XI0/XI37/XI11/MM7_g N_VSS_XI0/XI37/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM8 N_XI0/XI37/XI11/NET35_XI0/XI37/XI11/MM8_d
+ N_WL<71>_XI0/XI37/XI11/MM8_g N_BLN<4>_XI0/XI37/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI11/MM5 N_XI0/XI37/XI11/NET34_XI0/XI37/XI11/MM5_d
+ N_XI0/XI37/XI11/NET33_XI0/XI37/XI11/MM5_g N_VDD_XI0/XI37/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI11/MM4 N_XI0/XI37/XI11/NET33_XI0/XI37/XI11/MM4_d
+ N_XI0/XI37/XI11/NET34_XI0/XI37/XI11/MM4_g N_VDD_XI0/XI37/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI11/MM10 N_XI0/XI37/XI11/NET35_XI0/XI37/XI11/MM10_d
+ N_XI0/XI37/XI11/NET36_XI0/XI37/XI11/MM10_g N_VDD_XI0/XI37/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI11/MM11 N_XI0/XI37/XI11/NET36_XI0/XI37/XI11/MM11_d
+ N_XI0/XI37/XI11/NET35_XI0/XI37/XI11/MM11_g N_VDD_XI0/XI37/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI12/MM2 N_XI0/XI37/XI12/NET34_XI0/XI37/XI12/MM2_d
+ N_XI0/XI37/XI12/NET33_XI0/XI37/XI12/MM2_g N_VSS_XI0/XI37/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM3 N_XI0/XI37/XI12/NET33_XI0/XI37/XI12/MM3_d
+ N_WL<70>_XI0/XI37/XI12/MM3_g N_BLN<3>_XI0/XI37/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM0 N_XI0/XI37/XI12/NET34_XI0/XI37/XI12/MM0_d
+ N_WL<70>_XI0/XI37/XI12/MM0_g N_BL<3>_XI0/XI37/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM1 N_XI0/XI37/XI12/NET33_XI0/XI37/XI12/MM1_d
+ N_XI0/XI37/XI12/NET34_XI0/XI37/XI12/MM1_g N_VSS_XI0/XI37/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM9 N_XI0/XI37/XI12/NET36_XI0/XI37/XI12/MM9_d
+ N_WL<71>_XI0/XI37/XI12/MM9_g N_BL<3>_XI0/XI37/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM6 N_XI0/XI37/XI12/NET35_XI0/XI37/XI12/MM6_d
+ N_XI0/XI37/XI12/NET36_XI0/XI37/XI12/MM6_g N_VSS_XI0/XI37/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM7 N_XI0/XI37/XI12/NET36_XI0/XI37/XI12/MM7_d
+ N_XI0/XI37/XI12/NET35_XI0/XI37/XI12/MM7_g N_VSS_XI0/XI37/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM8 N_XI0/XI37/XI12/NET35_XI0/XI37/XI12/MM8_d
+ N_WL<71>_XI0/XI37/XI12/MM8_g N_BLN<3>_XI0/XI37/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI12/MM5 N_XI0/XI37/XI12/NET34_XI0/XI37/XI12/MM5_d
+ N_XI0/XI37/XI12/NET33_XI0/XI37/XI12/MM5_g N_VDD_XI0/XI37/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI12/MM4 N_XI0/XI37/XI12/NET33_XI0/XI37/XI12/MM4_d
+ N_XI0/XI37/XI12/NET34_XI0/XI37/XI12/MM4_g N_VDD_XI0/XI37/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI12/MM10 N_XI0/XI37/XI12/NET35_XI0/XI37/XI12/MM10_d
+ N_XI0/XI37/XI12/NET36_XI0/XI37/XI12/MM10_g N_VDD_XI0/XI37/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI12/MM11 N_XI0/XI37/XI12/NET36_XI0/XI37/XI12/MM11_d
+ N_XI0/XI37/XI12/NET35_XI0/XI37/XI12/MM11_g N_VDD_XI0/XI37/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI13/MM2 N_XI0/XI37/XI13/NET34_XI0/XI37/XI13/MM2_d
+ N_XI0/XI37/XI13/NET33_XI0/XI37/XI13/MM2_g N_VSS_XI0/XI37/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM3 N_XI0/XI37/XI13/NET33_XI0/XI37/XI13/MM3_d
+ N_WL<70>_XI0/XI37/XI13/MM3_g N_BLN<2>_XI0/XI37/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM0 N_XI0/XI37/XI13/NET34_XI0/XI37/XI13/MM0_d
+ N_WL<70>_XI0/XI37/XI13/MM0_g N_BL<2>_XI0/XI37/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM1 N_XI0/XI37/XI13/NET33_XI0/XI37/XI13/MM1_d
+ N_XI0/XI37/XI13/NET34_XI0/XI37/XI13/MM1_g N_VSS_XI0/XI37/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM9 N_XI0/XI37/XI13/NET36_XI0/XI37/XI13/MM9_d
+ N_WL<71>_XI0/XI37/XI13/MM9_g N_BL<2>_XI0/XI37/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM6 N_XI0/XI37/XI13/NET35_XI0/XI37/XI13/MM6_d
+ N_XI0/XI37/XI13/NET36_XI0/XI37/XI13/MM6_g N_VSS_XI0/XI37/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM7 N_XI0/XI37/XI13/NET36_XI0/XI37/XI13/MM7_d
+ N_XI0/XI37/XI13/NET35_XI0/XI37/XI13/MM7_g N_VSS_XI0/XI37/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM8 N_XI0/XI37/XI13/NET35_XI0/XI37/XI13/MM8_d
+ N_WL<71>_XI0/XI37/XI13/MM8_g N_BLN<2>_XI0/XI37/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI13/MM5 N_XI0/XI37/XI13/NET34_XI0/XI37/XI13/MM5_d
+ N_XI0/XI37/XI13/NET33_XI0/XI37/XI13/MM5_g N_VDD_XI0/XI37/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI13/MM4 N_XI0/XI37/XI13/NET33_XI0/XI37/XI13/MM4_d
+ N_XI0/XI37/XI13/NET34_XI0/XI37/XI13/MM4_g N_VDD_XI0/XI37/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI13/MM10 N_XI0/XI37/XI13/NET35_XI0/XI37/XI13/MM10_d
+ N_XI0/XI37/XI13/NET36_XI0/XI37/XI13/MM10_g N_VDD_XI0/XI37/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI13/MM11 N_XI0/XI37/XI13/NET36_XI0/XI37/XI13/MM11_d
+ N_XI0/XI37/XI13/NET35_XI0/XI37/XI13/MM11_g N_VDD_XI0/XI37/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI14/MM2 N_XI0/XI37/XI14/NET34_XI0/XI37/XI14/MM2_d
+ N_XI0/XI37/XI14/NET33_XI0/XI37/XI14/MM2_g N_VSS_XI0/XI37/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM3 N_XI0/XI37/XI14/NET33_XI0/XI37/XI14/MM3_d
+ N_WL<70>_XI0/XI37/XI14/MM3_g N_BLN<1>_XI0/XI37/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM0 N_XI0/XI37/XI14/NET34_XI0/XI37/XI14/MM0_d
+ N_WL<70>_XI0/XI37/XI14/MM0_g N_BL<1>_XI0/XI37/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM1 N_XI0/XI37/XI14/NET33_XI0/XI37/XI14/MM1_d
+ N_XI0/XI37/XI14/NET34_XI0/XI37/XI14/MM1_g N_VSS_XI0/XI37/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM9 N_XI0/XI37/XI14/NET36_XI0/XI37/XI14/MM9_d
+ N_WL<71>_XI0/XI37/XI14/MM9_g N_BL<1>_XI0/XI37/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM6 N_XI0/XI37/XI14/NET35_XI0/XI37/XI14/MM6_d
+ N_XI0/XI37/XI14/NET36_XI0/XI37/XI14/MM6_g N_VSS_XI0/XI37/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM7 N_XI0/XI37/XI14/NET36_XI0/XI37/XI14/MM7_d
+ N_XI0/XI37/XI14/NET35_XI0/XI37/XI14/MM7_g N_VSS_XI0/XI37/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM8 N_XI0/XI37/XI14/NET35_XI0/XI37/XI14/MM8_d
+ N_WL<71>_XI0/XI37/XI14/MM8_g N_BLN<1>_XI0/XI37/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI14/MM5 N_XI0/XI37/XI14/NET34_XI0/XI37/XI14/MM5_d
+ N_XI0/XI37/XI14/NET33_XI0/XI37/XI14/MM5_g N_VDD_XI0/XI37/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI14/MM4 N_XI0/XI37/XI14/NET33_XI0/XI37/XI14/MM4_d
+ N_XI0/XI37/XI14/NET34_XI0/XI37/XI14/MM4_g N_VDD_XI0/XI37/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI14/MM10 N_XI0/XI37/XI14/NET35_XI0/XI37/XI14/MM10_d
+ N_XI0/XI37/XI14/NET36_XI0/XI37/XI14/MM10_g N_VDD_XI0/XI37/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI14/MM11 N_XI0/XI37/XI14/NET36_XI0/XI37/XI14/MM11_d
+ N_XI0/XI37/XI14/NET35_XI0/XI37/XI14/MM11_g N_VDD_XI0/XI37/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI15/MM2 N_XI0/XI37/XI15/NET34_XI0/XI37/XI15/MM2_d
+ N_XI0/XI37/XI15/NET33_XI0/XI37/XI15/MM2_g N_VSS_XI0/XI37/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM3 N_XI0/XI37/XI15/NET33_XI0/XI37/XI15/MM3_d
+ N_WL<70>_XI0/XI37/XI15/MM3_g N_BLN<0>_XI0/XI37/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM0 N_XI0/XI37/XI15/NET34_XI0/XI37/XI15/MM0_d
+ N_WL<70>_XI0/XI37/XI15/MM0_g N_BL<0>_XI0/XI37/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM1 N_XI0/XI37/XI15/NET33_XI0/XI37/XI15/MM1_d
+ N_XI0/XI37/XI15/NET34_XI0/XI37/XI15/MM1_g N_VSS_XI0/XI37/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM9 N_XI0/XI37/XI15/NET36_XI0/XI37/XI15/MM9_d
+ N_WL<71>_XI0/XI37/XI15/MM9_g N_BL<0>_XI0/XI37/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM6 N_XI0/XI37/XI15/NET35_XI0/XI37/XI15/MM6_d
+ N_XI0/XI37/XI15/NET36_XI0/XI37/XI15/MM6_g N_VSS_XI0/XI37/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM7 N_XI0/XI37/XI15/NET36_XI0/XI37/XI15/MM7_d
+ N_XI0/XI37/XI15/NET35_XI0/XI37/XI15/MM7_g N_VSS_XI0/XI37/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM8 N_XI0/XI37/XI15/NET35_XI0/XI37/XI15/MM8_d
+ N_WL<71>_XI0/XI37/XI15/MM8_g N_BLN<0>_XI0/XI37/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI37/XI15/MM5 N_XI0/XI37/XI15/NET34_XI0/XI37/XI15/MM5_d
+ N_XI0/XI37/XI15/NET33_XI0/XI37/XI15/MM5_g N_VDD_XI0/XI37/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI15/MM4 N_XI0/XI37/XI15/NET33_XI0/XI37/XI15/MM4_d
+ N_XI0/XI37/XI15/NET34_XI0/XI37/XI15/MM4_g N_VDD_XI0/XI37/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI15/MM10 N_XI0/XI37/XI15/NET35_XI0/XI37/XI15/MM10_d
+ N_XI0/XI37/XI15/NET36_XI0/XI37/XI15/MM10_g N_VDD_XI0/XI37/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI37/XI15/MM11 N_XI0/XI37/XI15/NET36_XI0/XI37/XI15/MM11_d
+ N_XI0/XI37/XI15/NET35_XI0/XI37/XI15/MM11_g N_VDD_XI0/XI37/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI0/MM2 N_XI0/XI38/XI0/NET34_XI0/XI38/XI0/MM2_d
+ N_XI0/XI38/XI0/NET33_XI0/XI38/XI0/MM2_g N_VSS_XI0/XI38/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM3 N_XI0/XI38/XI0/NET33_XI0/XI38/XI0/MM3_d
+ N_WL<72>_XI0/XI38/XI0/MM3_g N_BLN<15>_XI0/XI38/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM0 N_XI0/XI38/XI0/NET34_XI0/XI38/XI0/MM0_d
+ N_WL<72>_XI0/XI38/XI0/MM0_g N_BL<15>_XI0/XI38/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM1 N_XI0/XI38/XI0/NET33_XI0/XI38/XI0/MM1_d
+ N_XI0/XI38/XI0/NET34_XI0/XI38/XI0/MM1_g N_VSS_XI0/XI38/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM9 N_XI0/XI38/XI0/NET36_XI0/XI38/XI0/MM9_d
+ N_WL<73>_XI0/XI38/XI0/MM9_g N_BL<15>_XI0/XI38/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM6 N_XI0/XI38/XI0/NET35_XI0/XI38/XI0/MM6_d
+ N_XI0/XI38/XI0/NET36_XI0/XI38/XI0/MM6_g N_VSS_XI0/XI38/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM7 N_XI0/XI38/XI0/NET36_XI0/XI38/XI0/MM7_d
+ N_XI0/XI38/XI0/NET35_XI0/XI38/XI0/MM7_g N_VSS_XI0/XI38/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM8 N_XI0/XI38/XI0/NET35_XI0/XI38/XI0/MM8_d
+ N_WL<73>_XI0/XI38/XI0/MM8_g N_BLN<15>_XI0/XI38/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI0/MM5 N_XI0/XI38/XI0/NET34_XI0/XI38/XI0/MM5_d
+ N_XI0/XI38/XI0/NET33_XI0/XI38/XI0/MM5_g N_VDD_XI0/XI38/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI0/MM4 N_XI0/XI38/XI0/NET33_XI0/XI38/XI0/MM4_d
+ N_XI0/XI38/XI0/NET34_XI0/XI38/XI0/MM4_g N_VDD_XI0/XI38/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI0/MM10 N_XI0/XI38/XI0/NET35_XI0/XI38/XI0/MM10_d
+ N_XI0/XI38/XI0/NET36_XI0/XI38/XI0/MM10_g N_VDD_XI0/XI38/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI0/MM11 N_XI0/XI38/XI0/NET36_XI0/XI38/XI0/MM11_d
+ N_XI0/XI38/XI0/NET35_XI0/XI38/XI0/MM11_g N_VDD_XI0/XI38/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI1/MM2 N_XI0/XI38/XI1/NET34_XI0/XI38/XI1/MM2_d
+ N_XI0/XI38/XI1/NET33_XI0/XI38/XI1/MM2_g N_VSS_XI0/XI38/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM3 N_XI0/XI38/XI1/NET33_XI0/XI38/XI1/MM3_d
+ N_WL<72>_XI0/XI38/XI1/MM3_g N_BLN<14>_XI0/XI38/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM0 N_XI0/XI38/XI1/NET34_XI0/XI38/XI1/MM0_d
+ N_WL<72>_XI0/XI38/XI1/MM0_g N_BL<14>_XI0/XI38/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM1 N_XI0/XI38/XI1/NET33_XI0/XI38/XI1/MM1_d
+ N_XI0/XI38/XI1/NET34_XI0/XI38/XI1/MM1_g N_VSS_XI0/XI38/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM9 N_XI0/XI38/XI1/NET36_XI0/XI38/XI1/MM9_d
+ N_WL<73>_XI0/XI38/XI1/MM9_g N_BL<14>_XI0/XI38/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM6 N_XI0/XI38/XI1/NET35_XI0/XI38/XI1/MM6_d
+ N_XI0/XI38/XI1/NET36_XI0/XI38/XI1/MM6_g N_VSS_XI0/XI38/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM7 N_XI0/XI38/XI1/NET36_XI0/XI38/XI1/MM7_d
+ N_XI0/XI38/XI1/NET35_XI0/XI38/XI1/MM7_g N_VSS_XI0/XI38/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM8 N_XI0/XI38/XI1/NET35_XI0/XI38/XI1/MM8_d
+ N_WL<73>_XI0/XI38/XI1/MM8_g N_BLN<14>_XI0/XI38/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI1/MM5 N_XI0/XI38/XI1/NET34_XI0/XI38/XI1/MM5_d
+ N_XI0/XI38/XI1/NET33_XI0/XI38/XI1/MM5_g N_VDD_XI0/XI38/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI1/MM4 N_XI0/XI38/XI1/NET33_XI0/XI38/XI1/MM4_d
+ N_XI0/XI38/XI1/NET34_XI0/XI38/XI1/MM4_g N_VDD_XI0/XI38/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI1/MM10 N_XI0/XI38/XI1/NET35_XI0/XI38/XI1/MM10_d
+ N_XI0/XI38/XI1/NET36_XI0/XI38/XI1/MM10_g N_VDD_XI0/XI38/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI1/MM11 N_XI0/XI38/XI1/NET36_XI0/XI38/XI1/MM11_d
+ N_XI0/XI38/XI1/NET35_XI0/XI38/XI1/MM11_g N_VDD_XI0/XI38/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI2/MM2 N_XI0/XI38/XI2/NET34_XI0/XI38/XI2/MM2_d
+ N_XI0/XI38/XI2/NET33_XI0/XI38/XI2/MM2_g N_VSS_XI0/XI38/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM3 N_XI0/XI38/XI2/NET33_XI0/XI38/XI2/MM3_d
+ N_WL<72>_XI0/XI38/XI2/MM3_g N_BLN<13>_XI0/XI38/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM0 N_XI0/XI38/XI2/NET34_XI0/XI38/XI2/MM0_d
+ N_WL<72>_XI0/XI38/XI2/MM0_g N_BL<13>_XI0/XI38/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM1 N_XI0/XI38/XI2/NET33_XI0/XI38/XI2/MM1_d
+ N_XI0/XI38/XI2/NET34_XI0/XI38/XI2/MM1_g N_VSS_XI0/XI38/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM9 N_XI0/XI38/XI2/NET36_XI0/XI38/XI2/MM9_d
+ N_WL<73>_XI0/XI38/XI2/MM9_g N_BL<13>_XI0/XI38/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM6 N_XI0/XI38/XI2/NET35_XI0/XI38/XI2/MM6_d
+ N_XI0/XI38/XI2/NET36_XI0/XI38/XI2/MM6_g N_VSS_XI0/XI38/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM7 N_XI0/XI38/XI2/NET36_XI0/XI38/XI2/MM7_d
+ N_XI0/XI38/XI2/NET35_XI0/XI38/XI2/MM7_g N_VSS_XI0/XI38/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM8 N_XI0/XI38/XI2/NET35_XI0/XI38/XI2/MM8_d
+ N_WL<73>_XI0/XI38/XI2/MM8_g N_BLN<13>_XI0/XI38/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI2/MM5 N_XI0/XI38/XI2/NET34_XI0/XI38/XI2/MM5_d
+ N_XI0/XI38/XI2/NET33_XI0/XI38/XI2/MM5_g N_VDD_XI0/XI38/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI2/MM4 N_XI0/XI38/XI2/NET33_XI0/XI38/XI2/MM4_d
+ N_XI0/XI38/XI2/NET34_XI0/XI38/XI2/MM4_g N_VDD_XI0/XI38/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI2/MM10 N_XI0/XI38/XI2/NET35_XI0/XI38/XI2/MM10_d
+ N_XI0/XI38/XI2/NET36_XI0/XI38/XI2/MM10_g N_VDD_XI0/XI38/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI2/MM11 N_XI0/XI38/XI2/NET36_XI0/XI38/XI2/MM11_d
+ N_XI0/XI38/XI2/NET35_XI0/XI38/XI2/MM11_g N_VDD_XI0/XI38/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI3/MM2 N_XI0/XI38/XI3/NET34_XI0/XI38/XI3/MM2_d
+ N_XI0/XI38/XI3/NET33_XI0/XI38/XI3/MM2_g N_VSS_XI0/XI38/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM3 N_XI0/XI38/XI3/NET33_XI0/XI38/XI3/MM3_d
+ N_WL<72>_XI0/XI38/XI3/MM3_g N_BLN<12>_XI0/XI38/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM0 N_XI0/XI38/XI3/NET34_XI0/XI38/XI3/MM0_d
+ N_WL<72>_XI0/XI38/XI3/MM0_g N_BL<12>_XI0/XI38/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM1 N_XI0/XI38/XI3/NET33_XI0/XI38/XI3/MM1_d
+ N_XI0/XI38/XI3/NET34_XI0/XI38/XI3/MM1_g N_VSS_XI0/XI38/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM9 N_XI0/XI38/XI3/NET36_XI0/XI38/XI3/MM9_d
+ N_WL<73>_XI0/XI38/XI3/MM9_g N_BL<12>_XI0/XI38/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM6 N_XI0/XI38/XI3/NET35_XI0/XI38/XI3/MM6_d
+ N_XI0/XI38/XI3/NET36_XI0/XI38/XI3/MM6_g N_VSS_XI0/XI38/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM7 N_XI0/XI38/XI3/NET36_XI0/XI38/XI3/MM7_d
+ N_XI0/XI38/XI3/NET35_XI0/XI38/XI3/MM7_g N_VSS_XI0/XI38/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM8 N_XI0/XI38/XI3/NET35_XI0/XI38/XI3/MM8_d
+ N_WL<73>_XI0/XI38/XI3/MM8_g N_BLN<12>_XI0/XI38/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI3/MM5 N_XI0/XI38/XI3/NET34_XI0/XI38/XI3/MM5_d
+ N_XI0/XI38/XI3/NET33_XI0/XI38/XI3/MM5_g N_VDD_XI0/XI38/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI3/MM4 N_XI0/XI38/XI3/NET33_XI0/XI38/XI3/MM4_d
+ N_XI0/XI38/XI3/NET34_XI0/XI38/XI3/MM4_g N_VDD_XI0/XI38/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI3/MM10 N_XI0/XI38/XI3/NET35_XI0/XI38/XI3/MM10_d
+ N_XI0/XI38/XI3/NET36_XI0/XI38/XI3/MM10_g N_VDD_XI0/XI38/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI3/MM11 N_XI0/XI38/XI3/NET36_XI0/XI38/XI3/MM11_d
+ N_XI0/XI38/XI3/NET35_XI0/XI38/XI3/MM11_g N_VDD_XI0/XI38/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI4/MM2 N_XI0/XI38/XI4/NET34_XI0/XI38/XI4/MM2_d
+ N_XI0/XI38/XI4/NET33_XI0/XI38/XI4/MM2_g N_VSS_XI0/XI38/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM3 N_XI0/XI38/XI4/NET33_XI0/XI38/XI4/MM3_d
+ N_WL<72>_XI0/XI38/XI4/MM3_g N_BLN<11>_XI0/XI38/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM0 N_XI0/XI38/XI4/NET34_XI0/XI38/XI4/MM0_d
+ N_WL<72>_XI0/XI38/XI4/MM0_g N_BL<11>_XI0/XI38/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM1 N_XI0/XI38/XI4/NET33_XI0/XI38/XI4/MM1_d
+ N_XI0/XI38/XI4/NET34_XI0/XI38/XI4/MM1_g N_VSS_XI0/XI38/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM9 N_XI0/XI38/XI4/NET36_XI0/XI38/XI4/MM9_d
+ N_WL<73>_XI0/XI38/XI4/MM9_g N_BL<11>_XI0/XI38/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM6 N_XI0/XI38/XI4/NET35_XI0/XI38/XI4/MM6_d
+ N_XI0/XI38/XI4/NET36_XI0/XI38/XI4/MM6_g N_VSS_XI0/XI38/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM7 N_XI0/XI38/XI4/NET36_XI0/XI38/XI4/MM7_d
+ N_XI0/XI38/XI4/NET35_XI0/XI38/XI4/MM7_g N_VSS_XI0/XI38/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM8 N_XI0/XI38/XI4/NET35_XI0/XI38/XI4/MM8_d
+ N_WL<73>_XI0/XI38/XI4/MM8_g N_BLN<11>_XI0/XI38/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI4/MM5 N_XI0/XI38/XI4/NET34_XI0/XI38/XI4/MM5_d
+ N_XI0/XI38/XI4/NET33_XI0/XI38/XI4/MM5_g N_VDD_XI0/XI38/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI4/MM4 N_XI0/XI38/XI4/NET33_XI0/XI38/XI4/MM4_d
+ N_XI0/XI38/XI4/NET34_XI0/XI38/XI4/MM4_g N_VDD_XI0/XI38/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI4/MM10 N_XI0/XI38/XI4/NET35_XI0/XI38/XI4/MM10_d
+ N_XI0/XI38/XI4/NET36_XI0/XI38/XI4/MM10_g N_VDD_XI0/XI38/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI4/MM11 N_XI0/XI38/XI4/NET36_XI0/XI38/XI4/MM11_d
+ N_XI0/XI38/XI4/NET35_XI0/XI38/XI4/MM11_g N_VDD_XI0/XI38/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI5/MM2 N_XI0/XI38/XI5/NET34_XI0/XI38/XI5/MM2_d
+ N_XI0/XI38/XI5/NET33_XI0/XI38/XI5/MM2_g N_VSS_XI0/XI38/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM3 N_XI0/XI38/XI5/NET33_XI0/XI38/XI5/MM3_d
+ N_WL<72>_XI0/XI38/XI5/MM3_g N_BLN<10>_XI0/XI38/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM0 N_XI0/XI38/XI5/NET34_XI0/XI38/XI5/MM0_d
+ N_WL<72>_XI0/XI38/XI5/MM0_g N_BL<10>_XI0/XI38/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM1 N_XI0/XI38/XI5/NET33_XI0/XI38/XI5/MM1_d
+ N_XI0/XI38/XI5/NET34_XI0/XI38/XI5/MM1_g N_VSS_XI0/XI38/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM9 N_XI0/XI38/XI5/NET36_XI0/XI38/XI5/MM9_d
+ N_WL<73>_XI0/XI38/XI5/MM9_g N_BL<10>_XI0/XI38/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM6 N_XI0/XI38/XI5/NET35_XI0/XI38/XI5/MM6_d
+ N_XI0/XI38/XI5/NET36_XI0/XI38/XI5/MM6_g N_VSS_XI0/XI38/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM7 N_XI0/XI38/XI5/NET36_XI0/XI38/XI5/MM7_d
+ N_XI0/XI38/XI5/NET35_XI0/XI38/XI5/MM7_g N_VSS_XI0/XI38/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM8 N_XI0/XI38/XI5/NET35_XI0/XI38/XI5/MM8_d
+ N_WL<73>_XI0/XI38/XI5/MM8_g N_BLN<10>_XI0/XI38/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI5/MM5 N_XI0/XI38/XI5/NET34_XI0/XI38/XI5/MM5_d
+ N_XI0/XI38/XI5/NET33_XI0/XI38/XI5/MM5_g N_VDD_XI0/XI38/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI5/MM4 N_XI0/XI38/XI5/NET33_XI0/XI38/XI5/MM4_d
+ N_XI0/XI38/XI5/NET34_XI0/XI38/XI5/MM4_g N_VDD_XI0/XI38/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI5/MM10 N_XI0/XI38/XI5/NET35_XI0/XI38/XI5/MM10_d
+ N_XI0/XI38/XI5/NET36_XI0/XI38/XI5/MM10_g N_VDD_XI0/XI38/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI5/MM11 N_XI0/XI38/XI5/NET36_XI0/XI38/XI5/MM11_d
+ N_XI0/XI38/XI5/NET35_XI0/XI38/XI5/MM11_g N_VDD_XI0/XI38/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI6/MM2 N_XI0/XI38/XI6/NET34_XI0/XI38/XI6/MM2_d
+ N_XI0/XI38/XI6/NET33_XI0/XI38/XI6/MM2_g N_VSS_XI0/XI38/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM3 N_XI0/XI38/XI6/NET33_XI0/XI38/XI6/MM3_d
+ N_WL<72>_XI0/XI38/XI6/MM3_g N_BLN<9>_XI0/XI38/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM0 N_XI0/XI38/XI6/NET34_XI0/XI38/XI6/MM0_d
+ N_WL<72>_XI0/XI38/XI6/MM0_g N_BL<9>_XI0/XI38/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM1 N_XI0/XI38/XI6/NET33_XI0/XI38/XI6/MM1_d
+ N_XI0/XI38/XI6/NET34_XI0/XI38/XI6/MM1_g N_VSS_XI0/XI38/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM9 N_XI0/XI38/XI6/NET36_XI0/XI38/XI6/MM9_d
+ N_WL<73>_XI0/XI38/XI6/MM9_g N_BL<9>_XI0/XI38/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM6 N_XI0/XI38/XI6/NET35_XI0/XI38/XI6/MM6_d
+ N_XI0/XI38/XI6/NET36_XI0/XI38/XI6/MM6_g N_VSS_XI0/XI38/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM7 N_XI0/XI38/XI6/NET36_XI0/XI38/XI6/MM7_d
+ N_XI0/XI38/XI6/NET35_XI0/XI38/XI6/MM7_g N_VSS_XI0/XI38/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM8 N_XI0/XI38/XI6/NET35_XI0/XI38/XI6/MM8_d
+ N_WL<73>_XI0/XI38/XI6/MM8_g N_BLN<9>_XI0/XI38/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI6/MM5 N_XI0/XI38/XI6/NET34_XI0/XI38/XI6/MM5_d
+ N_XI0/XI38/XI6/NET33_XI0/XI38/XI6/MM5_g N_VDD_XI0/XI38/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI6/MM4 N_XI0/XI38/XI6/NET33_XI0/XI38/XI6/MM4_d
+ N_XI0/XI38/XI6/NET34_XI0/XI38/XI6/MM4_g N_VDD_XI0/XI38/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI6/MM10 N_XI0/XI38/XI6/NET35_XI0/XI38/XI6/MM10_d
+ N_XI0/XI38/XI6/NET36_XI0/XI38/XI6/MM10_g N_VDD_XI0/XI38/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI6/MM11 N_XI0/XI38/XI6/NET36_XI0/XI38/XI6/MM11_d
+ N_XI0/XI38/XI6/NET35_XI0/XI38/XI6/MM11_g N_VDD_XI0/XI38/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI7/MM2 N_XI0/XI38/XI7/NET34_XI0/XI38/XI7/MM2_d
+ N_XI0/XI38/XI7/NET33_XI0/XI38/XI7/MM2_g N_VSS_XI0/XI38/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM3 N_XI0/XI38/XI7/NET33_XI0/XI38/XI7/MM3_d
+ N_WL<72>_XI0/XI38/XI7/MM3_g N_BLN<8>_XI0/XI38/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM0 N_XI0/XI38/XI7/NET34_XI0/XI38/XI7/MM0_d
+ N_WL<72>_XI0/XI38/XI7/MM0_g N_BL<8>_XI0/XI38/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM1 N_XI0/XI38/XI7/NET33_XI0/XI38/XI7/MM1_d
+ N_XI0/XI38/XI7/NET34_XI0/XI38/XI7/MM1_g N_VSS_XI0/XI38/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM9 N_XI0/XI38/XI7/NET36_XI0/XI38/XI7/MM9_d
+ N_WL<73>_XI0/XI38/XI7/MM9_g N_BL<8>_XI0/XI38/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM6 N_XI0/XI38/XI7/NET35_XI0/XI38/XI7/MM6_d
+ N_XI0/XI38/XI7/NET36_XI0/XI38/XI7/MM6_g N_VSS_XI0/XI38/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM7 N_XI0/XI38/XI7/NET36_XI0/XI38/XI7/MM7_d
+ N_XI0/XI38/XI7/NET35_XI0/XI38/XI7/MM7_g N_VSS_XI0/XI38/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM8 N_XI0/XI38/XI7/NET35_XI0/XI38/XI7/MM8_d
+ N_WL<73>_XI0/XI38/XI7/MM8_g N_BLN<8>_XI0/XI38/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI7/MM5 N_XI0/XI38/XI7/NET34_XI0/XI38/XI7/MM5_d
+ N_XI0/XI38/XI7/NET33_XI0/XI38/XI7/MM5_g N_VDD_XI0/XI38/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI7/MM4 N_XI0/XI38/XI7/NET33_XI0/XI38/XI7/MM4_d
+ N_XI0/XI38/XI7/NET34_XI0/XI38/XI7/MM4_g N_VDD_XI0/XI38/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI7/MM10 N_XI0/XI38/XI7/NET35_XI0/XI38/XI7/MM10_d
+ N_XI0/XI38/XI7/NET36_XI0/XI38/XI7/MM10_g N_VDD_XI0/XI38/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI7/MM11 N_XI0/XI38/XI7/NET36_XI0/XI38/XI7/MM11_d
+ N_XI0/XI38/XI7/NET35_XI0/XI38/XI7/MM11_g N_VDD_XI0/XI38/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI8/MM2 N_XI0/XI38/XI8/NET34_XI0/XI38/XI8/MM2_d
+ N_XI0/XI38/XI8/NET33_XI0/XI38/XI8/MM2_g N_VSS_XI0/XI38/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM3 N_XI0/XI38/XI8/NET33_XI0/XI38/XI8/MM3_d
+ N_WL<72>_XI0/XI38/XI8/MM3_g N_BLN<7>_XI0/XI38/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM0 N_XI0/XI38/XI8/NET34_XI0/XI38/XI8/MM0_d
+ N_WL<72>_XI0/XI38/XI8/MM0_g N_BL<7>_XI0/XI38/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM1 N_XI0/XI38/XI8/NET33_XI0/XI38/XI8/MM1_d
+ N_XI0/XI38/XI8/NET34_XI0/XI38/XI8/MM1_g N_VSS_XI0/XI38/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM9 N_XI0/XI38/XI8/NET36_XI0/XI38/XI8/MM9_d
+ N_WL<73>_XI0/XI38/XI8/MM9_g N_BL<7>_XI0/XI38/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM6 N_XI0/XI38/XI8/NET35_XI0/XI38/XI8/MM6_d
+ N_XI0/XI38/XI8/NET36_XI0/XI38/XI8/MM6_g N_VSS_XI0/XI38/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM7 N_XI0/XI38/XI8/NET36_XI0/XI38/XI8/MM7_d
+ N_XI0/XI38/XI8/NET35_XI0/XI38/XI8/MM7_g N_VSS_XI0/XI38/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM8 N_XI0/XI38/XI8/NET35_XI0/XI38/XI8/MM8_d
+ N_WL<73>_XI0/XI38/XI8/MM8_g N_BLN<7>_XI0/XI38/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI8/MM5 N_XI0/XI38/XI8/NET34_XI0/XI38/XI8/MM5_d
+ N_XI0/XI38/XI8/NET33_XI0/XI38/XI8/MM5_g N_VDD_XI0/XI38/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI8/MM4 N_XI0/XI38/XI8/NET33_XI0/XI38/XI8/MM4_d
+ N_XI0/XI38/XI8/NET34_XI0/XI38/XI8/MM4_g N_VDD_XI0/XI38/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI8/MM10 N_XI0/XI38/XI8/NET35_XI0/XI38/XI8/MM10_d
+ N_XI0/XI38/XI8/NET36_XI0/XI38/XI8/MM10_g N_VDD_XI0/XI38/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI8/MM11 N_XI0/XI38/XI8/NET36_XI0/XI38/XI8/MM11_d
+ N_XI0/XI38/XI8/NET35_XI0/XI38/XI8/MM11_g N_VDD_XI0/XI38/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI9/MM2 N_XI0/XI38/XI9/NET34_XI0/XI38/XI9/MM2_d
+ N_XI0/XI38/XI9/NET33_XI0/XI38/XI9/MM2_g N_VSS_XI0/XI38/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM3 N_XI0/XI38/XI9/NET33_XI0/XI38/XI9/MM3_d
+ N_WL<72>_XI0/XI38/XI9/MM3_g N_BLN<6>_XI0/XI38/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM0 N_XI0/XI38/XI9/NET34_XI0/XI38/XI9/MM0_d
+ N_WL<72>_XI0/XI38/XI9/MM0_g N_BL<6>_XI0/XI38/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM1 N_XI0/XI38/XI9/NET33_XI0/XI38/XI9/MM1_d
+ N_XI0/XI38/XI9/NET34_XI0/XI38/XI9/MM1_g N_VSS_XI0/XI38/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM9 N_XI0/XI38/XI9/NET36_XI0/XI38/XI9/MM9_d
+ N_WL<73>_XI0/XI38/XI9/MM9_g N_BL<6>_XI0/XI38/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM6 N_XI0/XI38/XI9/NET35_XI0/XI38/XI9/MM6_d
+ N_XI0/XI38/XI9/NET36_XI0/XI38/XI9/MM6_g N_VSS_XI0/XI38/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM7 N_XI0/XI38/XI9/NET36_XI0/XI38/XI9/MM7_d
+ N_XI0/XI38/XI9/NET35_XI0/XI38/XI9/MM7_g N_VSS_XI0/XI38/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM8 N_XI0/XI38/XI9/NET35_XI0/XI38/XI9/MM8_d
+ N_WL<73>_XI0/XI38/XI9/MM8_g N_BLN<6>_XI0/XI38/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI9/MM5 N_XI0/XI38/XI9/NET34_XI0/XI38/XI9/MM5_d
+ N_XI0/XI38/XI9/NET33_XI0/XI38/XI9/MM5_g N_VDD_XI0/XI38/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI9/MM4 N_XI0/XI38/XI9/NET33_XI0/XI38/XI9/MM4_d
+ N_XI0/XI38/XI9/NET34_XI0/XI38/XI9/MM4_g N_VDD_XI0/XI38/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI9/MM10 N_XI0/XI38/XI9/NET35_XI0/XI38/XI9/MM10_d
+ N_XI0/XI38/XI9/NET36_XI0/XI38/XI9/MM10_g N_VDD_XI0/XI38/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI9/MM11 N_XI0/XI38/XI9/NET36_XI0/XI38/XI9/MM11_d
+ N_XI0/XI38/XI9/NET35_XI0/XI38/XI9/MM11_g N_VDD_XI0/XI38/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI10/MM2 N_XI0/XI38/XI10/NET34_XI0/XI38/XI10/MM2_d
+ N_XI0/XI38/XI10/NET33_XI0/XI38/XI10/MM2_g N_VSS_XI0/XI38/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM3 N_XI0/XI38/XI10/NET33_XI0/XI38/XI10/MM3_d
+ N_WL<72>_XI0/XI38/XI10/MM3_g N_BLN<5>_XI0/XI38/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM0 N_XI0/XI38/XI10/NET34_XI0/XI38/XI10/MM0_d
+ N_WL<72>_XI0/XI38/XI10/MM0_g N_BL<5>_XI0/XI38/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM1 N_XI0/XI38/XI10/NET33_XI0/XI38/XI10/MM1_d
+ N_XI0/XI38/XI10/NET34_XI0/XI38/XI10/MM1_g N_VSS_XI0/XI38/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM9 N_XI0/XI38/XI10/NET36_XI0/XI38/XI10/MM9_d
+ N_WL<73>_XI0/XI38/XI10/MM9_g N_BL<5>_XI0/XI38/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM6 N_XI0/XI38/XI10/NET35_XI0/XI38/XI10/MM6_d
+ N_XI0/XI38/XI10/NET36_XI0/XI38/XI10/MM6_g N_VSS_XI0/XI38/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM7 N_XI0/XI38/XI10/NET36_XI0/XI38/XI10/MM7_d
+ N_XI0/XI38/XI10/NET35_XI0/XI38/XI10/MM7_g N_VSS_XI0/XI38/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM8 N_XI0/XI38/XI10/NET35_XI0/XI38/XI10/MM8_d
+ N_WL<73>_XI0/XI38/XI10/MM8_g N_BLN<5>_XI0/XI38/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI10/MM5 N_XI0/XI38/XI10/NET34_XI0/XI38/XI10/MM5_d
+ N_XI0/XI38/XI10/NET33_XI0/XI38/XI10/MM5_g N_VDD_XI0/XI38/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI10/MM4 N_XI0/XI38/XI10/NET33_XI0/XI38/XI10/MM4_d
+ N_XI0/XI38/XI10/NET34_XI0/XI38/XI10/MM4_g N_VDD_XI0/XI38/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI10/MM10 N_XI0/XI38/XI10/NET35_XI0/XI38/XI10/MM10_d
+ N_XI0/XI38/XI10/NET36_XI0/XI38/XI10/MM10_g N_VDD_XI0/XI38/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI10/MM11 N_XI0/XI38/XI10/NET36_XI0/XI38/XI10/MM11_d
+ N_XI0/XI38/XI10/NET35_XI0/XI38/XI10/MM11_g N_VDD_XI0/XI38/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI11/MM2 N_XI0/XI38/XI11/NET34_XI0/XI38/XI11/MM2_d
+ N_XI0/XI38/XI11/NET33_XI0/XI38/XI11/MM2_g N_VSS_XI0/XI38/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM3 N_XI0/XI38/XI11/NET33_XI0/XI38/XI11/MM3_d
+ N_WL<72>_XI0/XI38/XI11/MM3_g N_BLN<4>_XI0/XI38/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM0 N_XI0/XI38/XI11/NET34_XI0/XI38/XI11/MM0_d
+ N_WL<72>_XI0/XI38/XI11/MM0_g N_BL<4>_XI0/XI38/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM1 N_XI0/XI38/XI11/NET33_XI0/XI38/XI11/MM1_d
+ N_XI0/XI38/XI11/NET34_XI0/XI38/XI11/MM1_g N_VSS_XI0/XI38/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM9 N_XI0/XI38/XI11/NET36_XI0/XI38/XI11/MM9_d
+ N_WL<73>_XI0/XI38/XI11/MM9_g N_BL<4>_XI0/XI38/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM6 N_XI0/XI38/XI11/NET35_XI0/XI38/XI11/MM6_d
+ N_XI0/XI38/XI11/NET36_XI0/XI38/XI11/MM6_g N_VSS_XI0/XI38/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM7 N_XI0/XI38/XI11/NET36_XI0/XI38/XI11/MM7_d
+ N_XI0/XI38/XI11/NET35_XI0/XI38/XI11/MM7_g N_VSS_XI0/XI38/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM8 N_XI0/XI38/XI11/NET35_XI0/XI38/XI11/MM8_d
+ N_WL<73>_XI0/XI38/XI11/MM8_g N_BLN<4>_XI0/XI38/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI11/MM5 N_XI0/XI38/XI11/NET34_XI0/XI38/XI11/MM5_d
+ N_XI0/XI38/XI11/NET33_XI0/XI38/XI11/MM5_g N_VDD_XI0/XI38/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI11/MM4 N_XI0/XI38/XI11/NET33_XI0/XI38/XI11/MM4_d
+ N_XI0/XI38/XI11/NET34_XI0/XI38/XI11/MM4_g N_VDD_XI0/XI38/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI11/MM10 N_XI0/XI38/XI11/NET35_XI0/XI38/XI11/MM10_d
+ N_XI0/XI38/XI11/NET36_XI0/XI38/XI11/MM10_g N_VDD_XI0/XI38/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI11/MM11 N_XI0/XI38/XI11/NET36_XI0/XI38/XI11/MM11_d
+ N_XI0/XI38/XI11/NET35_XI0/XI38/XI11/MM11_g N_VDD_XI0/XI38/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI12/MM2 N_XI0/XI38/XI12/NET34_XI0/XI38/XI12/MM2_d
+ N_XI0/XI38/XI12/NET33_XI0/XI38/XI12/MM2_g N_VSS_XI0/XI38/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM3 N_XI0/XI38/XI12/NET33_XI0/XI38/XI12/MM3_d
+ N_WL<72>_XI0/XI38/XI12/MM3_g N_BLN<3>_XI0/XI38/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM0 N_XI0/XI38/XI12/NET34_XI0/XI38/XI12/MM0_d
+ N_WL<72>_XI0/XI38/XI12/MM0_g N_BL<3>_XI0/XI38/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM1 N_XI0/XI38/XI12/NET33_XI0/XI38/XI12/MM1_d
+ N_XI0/XI38/XI12/NET34_XI0/XI38/XI12/MM1_g N_VSS_XI0/XI38/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM9 N_XI0/XI38/XI12/NET36_XI0/XI38/XI12/MM9_d
+ N_WL<73>_XI0/XI38/XI12/MM9_g N_BL<3>_XI0/XI38/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM6 N_XI0/XI38/XI12/NET35_XI0/XI38/XI12/MM6_d
+ N_XI0/XI38/XI12/NET36_XI0/XI38/XI12/MM6_g N_VSS_XI0/XI38/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM7 N_XI0/XI38/XI12/NET36_XI0/XI38/XI12/MM7_d
+ N_XI0/XI38/XI12/NET35_XI0/XI38/XI12/MM7_g N_VSS_XI0/XI38/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM8 N_XI0/XI38/XI12/NET35_XI0/XI38/XI12/MM8_d
+ N_WL<73>_XI0/XI38/XI12/MM8_g N_BLN<3>_XI0/XI38/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI12/MM5 N_XI0/XI38/XI12/NET34_XI0/XI38/XI12/MM5_d
+ N_XI0/XI38/XI12/NET33_XI0/XI38/XI12/MM5_g N_VDD_XI0/XI38/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI12/MM4 N_XI0/XI38/XI12/NET33_XI0/XI38/XI12/MM4_d
+ N_XI0/XI38/XI12/NET34_XI0/XI38/XI12/MM4_g N_VDD_XI0/XI38/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI12/MM10 N_XI0/XI38/XI12/NET35_XI0/XI38/XI12/MM10_d
+ N_XI0/XI38/XI12/NET36_XI0/XI38/XI12/MM10_g N_VDD_XI0/XI38/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI12/MM11 N_XI0/XI38/XI12/NET36_XI0/XI38/XI12/MM11_d
+ N_XI0/XI38/XI12/NET35_XI0/XI38/XI12/MM11_g N_VDD_XI0/XI38/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI13/MM2 N_XI0/XI38/XI13/NET34_XI0/XI38/XI13/MM2_d
+ N_XI0/XI38/XI13/NET33_XI0/XI38/XI13/MM2_g N_VSS_XI0/XI38/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM3 N_XI0/XI38/XI13/NET33_XI0/XI38/XI13/MM3_d
+ N_WL<72>_XI0/XI38/XI13/MM3_g N_BLN<2>_XI0/XI38/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM0 N_XI0/XI38/XI13/NET34_XI0/XI38/XI13/MM0_d
+ N_WL<72>_XI0/XI38/XI13/MM0_g N_BL<2>_XI0/XI38/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM1 N_XI0/XI38/XI13/NET33_XI0/XI38/XI13/MM1_d
+ N_XI0/XI38/XI13/NET34_XI0/XI38/XI13/MM1_g N_VSS_XI0/XI38/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM9 N_XI0/XI38/XI13/NET36_XI0/XI38/XI13/MM9_d
+ N_WL<73>_XI0/XI38/XI13/MM9_g N_BL<2>_XI0/XI38/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM6 N_XI0/XI38/XI13/NET35_XI0/XI38/XI13/MM6_d
+ N_XI0/XI38/XI13/NET36_XI0/XI38/XI13/MM6_g N_VSS_XI0/XI38/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM7 N_XI0/XI38/XI13/NET36_XI0/XI38/XI13/MM7_d
+ N_XI0/XI38/XI13/NET35_XI0/XI38/XI13/MM7_g N_VSS_XI0/XI38/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM8 N_XI0/XI38/XI13/NET35_XI0/XI38/XI13/MM8_d
+ N_WL<73>_XI0/XI38/XI13/MM8_g N_BLN<2>_XI0/XI38/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI13/MM5 N_XI0/XI38/XI13/NET34_XI0/XI38/XI13/MM5_d
+ N_XI0/XI38/XI13/NET33_XI0/XI38/XI13/MM5_g N_VDD_XI0/XI38/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI13/MM4 N_XI0/XI38/XI13/NET33_XI0/XI38/XI13/MM4_d
+ N_XI0/XI38/XI13/NET34_XI0/XI38/XI13/MM4_g N_VDD_XI0/XI38/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI13/MM10 N_XI0/XI38/XI13/NET35_XI0/XI38/XI13/MM10_d
+ N_XI0/XI38/XI13/NET36_XI0/XI38/XI13/MM10_g N_VDD_XI0/XI38/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI13/MM11 N_XI0/XI38/XI13/NET36_XI0/XI38/XI13/MM11_d
+ N_XI0/XI38/XI13/NET35_XI0/XI38/XI13/MM11_g N_VDD_XI0/XI38/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI14/MM2 N_XI0/XI38/XI14/NET34_XI0/XI38/XI14/MM2_d
+ N_XI0/XI38/XI14/NET33_XI0/XI38/XI14/MM2_g N_VSS_XI0/XI38/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM3 N_XI0/XI38/XI14/NET33_XI0/XI38/XI14/MM3_d
+ N_WL<72>_XI0/XI38/XI14/MM3_g N_BLN<1>_XI0/XI38/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM0 N_XI0/XI38/XI14/NET34_XI0/XI38/XI14/MM0_d
+ N_WL<72>_XI0/XI38/XI14/MM0_g N_BL<1>_XI0/XI38/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM1 N_XI0/XI38/XI14/NET33_XI0/XI38/XI14/MM1_d
+ N_XI0/XI38/XI14/NET34_XI0/XI38/XI14/MM1_g N_VSS_XI0/XI38/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM9 N_XI0/XI38/XI14/NET36_XI0/XI38/XI14/MM9_d
+ N_WL<73>_XI0/XI38/XI14/MM9_g N_BL<1>_XI0/XI38/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM6 N_XI0/XI38/XI14/NET35_XI0/XI38/XI14/MM6_d
+ N_XI0/XI38/XI14/NET36_XI0/XI38/XI14/MM6_g N_VSS_XI0/XI38/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM7 N_XI0/XI38/XI14/NET36_XI0/XI38/XI14/MM7_d
+ N_XI0/XI38/XI14/NET35_XI0/XI38/XI14/MM7_g N_VSS_XI0/XI38/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM8 N_XI0/XI38/XI14/NET35_XI0/XI38/XI14/MM8_d
+ N_WL<73>_XI0/XI38/XI14/MM8_g N_BLN<1>_XI0/XI38/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI14/MM5 N_XI0/XI38/XI14/NET34_XI0/XI38/XI14/MM5_d
+ N_XI0/XI38/XI14/NET33_XI0/XI38/XI14/MM5_g N_VDD_XI0/XI38/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI14/MM4 N_XI0/XI38/XI14/NET33_XI0/XI38/XI14/MM4_d
+ N_XI0/XI38/XI14/NET34_XI0/XI38/XI14/MM4_g N_VDD_XI0/XI38/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI14/MM10 N_XI0/XI38/XI14/NET35_XI0/XI38/XI14/MM10_d
+ N_XI0/XI38/XI14/NET36_XI0/XI38/XI14/MM10_g N_VDD_XI0/XI38/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI14/MM11 N_XI0/XI38/XI14/NET36_XI0/XI38/XI14/MM11_d
+ N_XI0/XI38/XI14/NET35_XI0/XI38/XI14/MM11_g N_VDD_XI0/XI38/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI15/MM2 N_XI0/XI38/XI15/NET34_XI0/XI38/XI15/MM2_d
+ N_XI0/XI38/XI15/NET33_XI0/XI38/XI15/MM2_g N_VSS_XI0/XI38/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM3 N_XI0/XI38/XI15/NET33_XI0/XI38/XI15/MM3_d
+ N_WL<72>_XI0/XI38/XI15/MM3_g N_BLN<0>_XI0/XI38/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM0 N_XI0/XI38/XI15/NET34_XI0/XI38/XI15/MM0_d
+ N_WL<72>_XI0/XI38/XI15/MM0_g N_BL<0>_XI0/XI38/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM1 N_XI0/XI38/XI15/NET33_XI0/XI38/XI15/MM1_d
+ N_XI0/XI38/XI15/NET34_XI0/XI38/XI15/MM1_g N_VSS_XI0/XI38/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM9 N_XI0/XI38/XI15/NET36_XI0/XI38/XI15/MM9_d
+ N_WL<73>_XI0/XI38/XI15/MM9_g N_BL<0>_XI0/XI38/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM6 N_XI0/XI38/XI15/NET35_XI0/XI38/XI15/MM6_d
+ N_XI0/XI38/XI15/NET36_XI0/XI38/XI15/MM6_g N_VSS_XI0/XI38/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM7 N_XI0/XI38/XI15/NET36_XI0/XI38/XI15/MM7_d
+ N_XI0/XI38/XI15/NET35_XI0/XI38/XI15/MM7_g N_VSS_XI0/XI38/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM8 N_XI0/XI38/XI15/NET35_XI0/XI38/XI15/MM8_d
+ N_WL<73>_XI0/XI38/XI15/MM8_g N_BLN<0>_XI0/XI38/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI38/XI15/MM5 N_XI0/XI38/XI15/NET34_XI0/XI38/XI15/MM5_d
+ N_XI0/XI38/XI15/NET33_XI0/XI38/XI15/MM5_g N_VDD_XI0/XI38/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI15/MM4 N_XI0/XI38/XI15/NET33_XI0/XI38/XI15/MM4_d
+ N_XI0/XI38/XI15/NET34_XI0/XI38/XI15/MM4_g N_VDD_XI0/XI38/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI15/MM10 N_XI0/XI38/XI15/NET35_XI0/XI38/XI15/MM10_d
+ N_XI0/XI38/XI15/NET36_XI0/XI38/XI15/MM10_g N_VDD_XI0/XI38/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI38/XI15/MM11 N_XI0/XI38/XI15/NET36_XI0/XI38/XI15/MM11_d
+ N_XI0/XI38/XI15/NET35_XI0/XI38/XI15/MM11_g N_VDD_XI0/XI38/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI0/MM2 N_XI0/XI39/XI0/NET34_XI0/XI39/XI0/MM2_d
+ N_XI0/XI39/XI0/NET33_XI0/XI39/XI0/MM2_g N_VSS_XI0/XI39/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM3 N_XI0/XI39/XI0/NET33_XI0/XI39/XI0/MM3_d
+ N_WL<74>_XI0/XI39/XI0/MM3_g N_BLN<15>_XI0/XI39/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM0 N_XI0/XI39/XI0/NET34_XI0/XI39/XI0/MM0_d
+ N_WL<74>_XI0/XI39/XI0/MM0_g N_BL<15>_XI0/XI39/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM1 N_XI0/XI39/XI0/NET33_XI0/XI39/XI0/MM1_d
+ N_XI0/XI39/XI0/NET34_XI0/XI39/XI0/MM1_g N_VSS_XI0/XI39/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM9 N_XI0/XI39/XI0/NET36_XI0/XI39/XI0/MM9_d
+ N_WL<75>_XI0/XI39/XI0/MM9_g N_BL<15>_XI0/XI39/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM6 N_XI0/XI39/XI0/NET35_XI0/XI39/XI0/MM6_d
+ N_XI0/XI39/XI0/NET36_XI0/XI39/XI0/MM6_g N_VSS_XI0/XI39/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM7 N_XI0/XI39/XI0/NET36_XI0/XI39/XI0/MM7_d
+ N_XI0/XI39/XI0/NET35_XI0/XI39/XI0/MM7_g N_VSS_XI0/XI39/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM8 N_XI0/XI39/XI0/NET35_XI0/XI39/XI0/MM8_d
+ N_WL<75>_XI0/XI39/XI0/MM8_g N_BLN<15>_XI0/XI39/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI0/MM5 N_XI0/XI39/XI0/NET34_XI0/XI39/XI0/MM5_d
+ N_XI0/XI39/XI0/NET33_XI0/XI39/XI0/MM5_g N_VDD_XI0/XI39/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI0/MM4 N_XI0/XI39/XI0/NET33_XI0/XI39/XI0/MM4_d
+ N_XI0/XI39/XI0/NET34_XI0/XI39/XI0/MM4_g N_VDD_XI0/XI39/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI0/MM10 N_XI0/XI39/XI0/NET35_XI0/XI39/XI0/MM10_d
+ N_XI0/XI39/XI0/NET36_XI0/XI39/XI0/MM10_g N_VDD_XI0/XI39/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI0/MM11 N_XI0/XI39/XI0/NET36_XI0/XI39/XI0/MM11_d
+ N_XI0/XI39/XI0/NET35_XI0/XI39/XI0/MM11_g N_VDD_XI0/XI39/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI1/MM2 N_XI0/XI39/XI1/NET34_XI0/XI39/XI1/MM2_d
+ N_XI0/XI39/XI1/NET33_XI0/XI39/XI1/MM2_g N_VSS_XI0/XI39/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM3 N_XI0/XI39/XI1/NET33_XI0/XI39/XI1/MM3_d
+ N_WL<74>_XI0/XI39/XI1/MM3_g N_BLN<14>_XI0/XI39/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM0 N_XI0/XI39/XI1/NET34_XI0/XI39/XI1/MM0_d
+ N_WL<74>_XI0/XI39/XI1/MM0_g N_BL<14>_XI0/XI39/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM1 N_XI0/XI39/XI1/NET33_XI0/XI39/XI1/MM1_d
+ N_XI0/XI39/XI1/NET34_XI0/XI39/XI1/MM1_g N_VSS_XI0/XI39/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM9 N_XI0/XI39/XI1/NET36_XI0/XI39/XI1/MM9_d
+ N_WL<75>_XI0/XI39/XI1/MM9_g N_BL<14>_XI0/XI39/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM6 N_XI0/XI39/XI1/NET35_XI0/XI39/XI1/MM6_d
+ N_XI0/XI39/XI1/NET36_XI0/XI39/XI1/MM6_g N_VSS_XI0/XI39/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM7 N_XI0/XI39/XI1/NET36_XI0/XI39/XI1/MM7_d
+ N_XI0/XI39/XI1/NET35_XI0/XI39/XI1/MM7_g N_VSS_XI0/XI39/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM8 N_XI0/XI39/XI1/NET35_XI0/XI39/XI1/MM8_d
+ N_WL<75>_XI0/XI39/XI1/MM8_g N_BLN<14>_XI0/XI39/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI1/MM5 N_XI0/XI39/XI1/NET34_XI0/XI39/XI1/MM5_d
+ N_XI0/XI39/XI1/NET33_XI0/XI39/XI1/MM5_g N_VDD_XI0/XI39/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI1/MM4 N_XI0/XI39/XI1/NET33_XI0/XI39/XI1/MM4_d
+ N_XI0/XI39/XI1/NET34_XI0/XI39/XI1/MM4_g N_VDD_XI0/XI39/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI1/MM10 N_XI0/XI39/XI1/NET35_XI0/XI39/XI1/MM10_d
+ N_XI0/XI39/XI1/NET36_XI0/XI39/XI1/MM10_g N_VDD_XI0/XI39/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI1/MM11 N_XI0/XI39/XI1/NET36_XI0/XI39/XI1/MM11_d
+ N_XI0/XI39/XI1/NET35_XI0/XI39/XI1/MM11_g N_VDD_XI0/XI39/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI2/MM2 N_XI0/XI39/XI2/NET34_XI0/XI39/XI2/MM2_d
+ N_XI0/XI39/XI2/NET33_XI0/XI39/XI2/MM2_g N_VSS_XI0/XI39/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM3 N_XI0/XI39/XI2/NET33_XI0/XI39/XI2/MM3_d
+ N_WL<74>_XI0/XI39/XI2/MM3_g N_BLN<13>_XI0/XI39/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM0 N_XI0/XI39/XI2/NET34_XI0/XI39/XI2/MM0_d
+ N_WL<74>_XI0/XI39/XI2/MM0_g N_BL<13>_XI0/XI39/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM1 N_XI0/XI39/XI2/NET33_XI0/XI39/XI2/MM1_d
+ N_XI0/XI39/XI2/NET34_XI0/XI39/XI2/MM1_g N_VSS_XI0/XI39/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM9 N_XI0/XI39/XI2/NET36_XI0/XI39/XI2/MM9_d
+ N_WL<75>_XI0/XI39/XI2/MM9_g N_BL<13>_XI0/XI39/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM6 N_XI0/XI39/XI2/NET35_XI0/XI39/XI2/MM6_d
+ N_XI0/XI39/XI2/NET36_XI0/XI39/XI2/MM6_g N_VSS_XI0/XI39/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM7 N_XI0/XI39/XI2/NET36_XI0/XI39/XI2/MM7_d
+ N_XI0/XI39/XI2/NET35_XI0/XI39/XI2/MM7_g N_VSS_XI0/XI39/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM8 N_XI0/XI39/XI2/NET35_XI0/XI39/XI2/MM8_d
+ N_WL<75>_XI0/XI39/XI2/MM8_g N_BLN<13>_XI0/XI39/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI2/MM5 N_XI0/XI39/XI2/NET34_XI0/XI39/XI2/MM5_d
+ N_XI0/XI39/XI2/NET33_XI0/XI39/XI2/MM5_g N_VDD_XI0/XI39/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI2/MM4 N_XI0/XI39/XI2/NET33_XI0/XI39/XI2/MM4_d
+ N_XI0/XI39/XI2/NET34_XI0/XI39/XI2/MM4_g N_VDD_XI0/XI39/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI2/MM10 N_XI0/XI39/XI2/NET35_XI0/XI39/XI2/MM10_d
+ N_XI0/XI39/XI2/NET36_XI0/XI39/XI2/MM10_g N_VDD_XI0/XI39/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI2/MM11 N_XI0/XI39/XI2/NET36_XI0/XI39/XI2/MM11_d
+ N_XI0/XI39/XI2/NET35_XI0/XI39/XI2/MM11_g N_VDD_XI0/XI39/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI3/MM2 N_XI0/XI39/XI3/NET34_XI0/XI39/XI3/MM2_d
+ N_XI0/XI39/XI3/NET33_XI0/XI39/XI3/MM2_g N_VSS_XI0/XI39/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM3 N_XI0/XI39/XI3/NET33_XI0/XI39/XI3/MM3_d
+ N_WL<74>_XI0/XI39/XI3/MM3_g N_BLN<12>_XI0/XI39/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM0 N_XI0/XI39/XI3/NET34_XI0/XI39/XI3/MM0_d
+ N_WL<74>_XI0/XI39/XI3/MM0_g N_BL<12>_XI0/XI39/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM1 N_XI0/XI39/XI3/NET33_XI0/XI39/XI3/MM1_d
+ N_XI0/XI39/XI3/NET34_XI0/XI39/XI3/MM1_g N_VSS_XI0/XI39/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM9 N_XI0/XI39/XI3/NET36_XI0/XI39/XI3/MM9_d
+ N_WL<75>_XI0/XI39/XI3/MM9_g N_BL<12>_XI0/XI39/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM6 N_XI0/XI39/XI3/NET35_XI0/XI39/XI3/MM6_d
+ N_XI0/XI39/XI3/NET36_XI0/XI39/XI3/MM6_g N_VSS_XI0/XI39/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM7 N_XI0/XI39/XI3/NET36_XI0/XI39/XI3/MM7_d
+ N_XI0/XI39/XI3/NET35_XI0/XI39/XI3/MM7_g N_VSS_XI0/XI39/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM8 N_XI0/XI39/XI3/NET35_XI0/XI39/XI3/MM8_d
+ N_WL<75>_XI0/XI39/XI3/MM8_g N_BLN<12>_XI0/XI39/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI3/MM5 N_XI0/XI39/XI3/NET34_XI0/XI39/XI3/MM5_d
+ N_XI0/XI39/XI3/NET33_XI0/XI39/XI3/MM5_g N_VDD_XI0/XI39/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI3/MM4 N_XI0/XI39/XI3/NET33_XI0/XI39/XI3/MM4_d
+ N_XI0/XI39/XI3/NET34_XI0/XI39/XI3/MM4_g N_VDD_XI0/XI39/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI3/MM10 N_XI0/XI39/XI3/NET35_XI0/XI39/XI3/MM10_d
+ N_XI0/XI39/XI3/NET36_XI0/XI39/XI3/MM10_g N_VDD_XI0/XI39/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI3/MM11 N_XI0/XI39/XI3/NET36_XI0/XI39/XI3/MM11_d
+ N_XI0/XI39/XI3/NET35_XI0/XI39/XI3/MM11_g N_VDD_XI0/XI39/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI4/MM2 N_XI0/XI39/XI4/NET34_XI0/XI39/XI4/MM2_d
+ N_XI0/XI39/XI4/NET33_XI0/XI39/XI4/MM2_g N_VSS_XI0/XI39/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM3 N_XI0/XI39/XI4/NET33_XI0/XI39/XI4/MM3_d
+ N_WL<74>_XI0/XI39/XI4/MM3_g N_BLN<11>_XI0/XI39/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM0 N_XI0/XI39/XI4/NET34_XI0/XI39/XI4/MM0_d
+ N_WL<74>_XI0/XI39/XI4/MM0_g N_BL<11>_XI0/XI39/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM1 N_XI0/XI39/XI4/NET33_XI0/XI39/XI4/MM1_d
+ N_XI0/XI39/XI4/NET34_XI0/XI39/XI4/MM1_g N_VSS_XI0/XI39/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM9 N_XI0/XI39/XI4/NET36_XI0/XI39/XI4/MM9_d
+ N_WL<75>_XI0/XI39/XI4/MM9_g N_BL<11>_XI0/XI39/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM6 N_XI0/XI39/XI4/NET35_XI0/XI39/XI4/MM6_d
+ N_XI0/XI39/XI4/NET36_XI0/XI39/XI4/MM6_g N_VSS_XI0/XI39/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM7 N_XI0/XI39/XI4/NET36_XI0/XI39/XI4/MM7_d
+ N_XI0/XI39/XI4/NET35_XI0/XI39/XI4/MM7_g N_VSS_XI0/XI39/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM8 N_XI0/XI39/XI4/NET35_XI0/XI39/XI4/MM8_d
+ N_WL<75>_XI0/XI39/XI4/MM8_g N_BLN<11>_XI0/XI39/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI4/MM5 N_XI0/XI39/XI4/NET34_XI0/XI39/XI4/MM5_d
+ N_XI0/XI39/XI4/NET33_XI0/XI39/XI4/MM5_g N_VDD_XI0/XI39/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI4/MM4 N_XI0/XI39/XI4/NET33_XI0/XI39/XI4/MM4_d
+ N_XI0/XI39/XI4/NET34_XI0/XI39/XI4/MM4_g N_VDD_XI0/XI39/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI4/MM10 N_XI0/XI39/XI4/NET35_XI0/XI39/XI4/MM10_d
+ N_XI0/XI39/XI4/NET36_XI0/XI39/XI4/MM10_g N_VDD_XI0/XI39/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI4/MM11 N_XI0/XI39/XI4/NET36_XI0/XI39/XI4/MM11_d
+ N_XI0/XI39/XI4/NET35_XI0/XI39/XI4/MM11_g N_VDD_XI0/XI39/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI5/MM2 N_XI0/XI39/XI5/NET34_XI0/XI39/XI5/MM2_d
+ N_XI0/XI39/XI5/NET33_XI0/XI39/XI5/MM2_g N_VSS_XI0/XI39/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM3 N_XI0/XI39/XI5/NET33_XI0/XI39/XI5/MM3_d
+ N_WL<74>_XI0/XI39/XI5/MM3_g N_BLN<10>_XI0/XI39/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM0 N_XI0/XI39/XI5/NET34_XI0/XI39/XI5/MM0_d
+ N_WL<74>_XI0/XI39/XI5/MM0_g N_BL<10>_XI0/XI39/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM1 N_XI0/XI39/XI5/NET33_XI0/XI39/XI5/MM1_d
+ N_XI0/XI39/XI5/NET34_XI0/XI39/XI5/MM1_g N_VSS_XI0/XI39/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM9 N_XI0/XI39/XI5/NET36_XI0/XI39/XI5/MM9_d
+ N_WL<75>_XI0/XI39/XI5/MM9_g N_BL<10>_XI0/XI39/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM6 N_XI0/XI39/XI5/NET35_XI0/XI39/XI5/MM6_d
+ N_XI0/XI39/XI5/NET36_XI0/XI39/XI5/MM6_g N_VSS_XI0/XI39/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM7 N_XI0/XI39/XI5/NET36_XI0/XI39/XI5/MM7_d
+ N_XI0/XI39/XI5/NET35_XI0/XI39/XI5/MM7_g N_VSS_XI0/XI39/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM8 N_XI0/XI39/XI5/NET35_XI0/XI39/XI5/MM8_d
+ N_WL<75>_XI0/XI39/XI5/MM8_g N_BLN<10>_XI0/XI39/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI5/MM5 N_XI0/XI39/XI5/NET34_XI0/XI39/XI5/MM5_d
+ N_XI0/XI39/XI5/NET33_XI0/XI39/XI5/MM5_g N_VDD_XI0/XI39/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI5/MM4 N_XI0/XI39/XI5/NET33_XI0/XI39/XI5/MM4_d
+ N_XI0/XI39/XI5/NET34_XI0/XI39/XI5/MM4_g N_VDD_XI0/XI39/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI5/MM10 N_XI0/XI39/XI5/NET35_XI0/XI39/XI5/MM10_d
+ N_XI0/XI39/XI5/NET36_XI0/XI39/XI5/MM10_g N_VDD_XI0/XI39/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI5/MM11 N_XI0/XI39/XI5/NET36_XI0/XI39/XI5/MM11_d
+ N_XI0/XI39/XI5/NET35_XI0/XI39/XI5/MM11_g N_VDD_XI0/XI39/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI6/MM2 N_XI0/XI39/XI6/NET34_XI0/XI39/XI6/MM2_d
+ N_XI0/XI39/XI6/NET33_XI0/XI39/XI6/MM2_g N_VSS_XI0/XI39/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM3 N_XI0/XI39/XI6/NET33_XI0/XI39/XI6/MM3_d
+ N_WL<74>_XI0/XI39/XI6/MM3_g N_BLN<9>_XI0/XI39/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM0 N_XI0/XI39/XI6/NET34_XI0/XI39/XI6/MM0_d
+ N_WL<74>_XI0/XI39/XI6/MM0_g N_BL<9>_XI0/XI39/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM1 N_XI0/XI39/XI6/NET33_XI0/XI39/XI6/MM1_d
+ N_XI0/XI39/XI6/NET34_XI0/XI39/XI6/MM1_g N_VSS_XI0/XI39/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM9 N_XI0/XI39/XI6/NET36_XI0/XI39/XI6/MM9_d
+ N_WL<75>_XI0/XI39/XI6/MM9_g N_BL<9>_XI0/XI39/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM6 N_XI0/XI39/XI6/NET35_XI0/XI39/XI6/MM6_d
+ N_XI0/XI39/XI6/NET36_XI0/XI39/XI6/MM6_g N_VSS_XI0/XI39/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM7 N_XI0/XI39/XI6/NET36_XI0/XI39/XI6/MM7_d
+ N_XI0/XI39/XI6/NET35_XI0/XI39/XI6/MM7_g N_VSS_XI0/XI39/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM8 N_XI0/XI39/XI6/NET35_XI0/XI39/XI6/MM8_d
+ N_WL<75>_XI0/XI39/XI6/MM8_g N_BLN<9>_XI0/XI39/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI6/MM5 N_XI0/XI39/XI6/NET34_XI0/XI39/XI6/MM5_d
+ N_XI0/XI39/XI6/NET33_XI0/XI39/XI6/MM5_g N_VDD_XI0/XI39/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI6/MM4 N_XI0/XI39/XI6/NET33_XI0/XI39/XI6/MM4_d
+ N_XI0/XI39/XI6/NET34_XI0/XI39/XI6/MM4_g N_VDD_XI0/XI39/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI6/MM10 N_XI0/XI39/XI6/NET35_XI0/XI39/XI6/MM10_d
+ N_XI0/XI39/XI6/NET36_XI0/XI39/XI6/MM10_g N_VDD_XI0/XI39/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI6/MM11 N_XI0/XI39/XI6/NET36_XI0/XI39/XI6/MM11_d
+ N_XI0/XI39/XI6/NET35_XI0/XI39/XI6/MM11_g N_VDD_XI0/XI39/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI7/MM2 N_XI0/XI39/XI7/NET34_XI0/XI39/XI7/MM2_d
+ N_XI0/XI39/XI7/NET33_XI0/XI39/XI7/MM2_g N_VSS_XI0/XI39/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM3 N_XI0/XI39/XI7/NET33_XI0/XI39/XI7/MM3_d
+ N_WL<74>_XI0/XI39/XI7/MM3_g N_BLN<8>_XI0/XI39/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM0 N_XI0/XI39/XI7/NET34_XI0/XI39/XI7/MM0_d
+ N_WL<74>_XI0/XI39/XI7/MM0_g N_BL<8>_XI0/XI39/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM1 N_XI0/XI39/XI7/NET33_XI0/XI39/XI7/MM1_d
+ N_XI0/XI39/XI7/NET34_XI0/XI39/XI7/MM1_g N_VSS_XI0/XI39/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM9 N_XI0/XI39/XI7/NET36_XI0/XI39/XI7/MM9_d
+ N_WL<75>_XI0/XI39/XI7/MM9_g N_BL<8>_XI0/XI39/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM6 N_XI0/XI39/XI7/NET35_XI0/XI39/XI7/MM6_d
+ N_XI0/XI39/XI7/NET36_XI0/XI39/XI7/MM6_g N_VSS_XI0/XI39/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM7 N_XI0/XI39/XI7/NET36_XI0/XI39/XI7/MM7_d
+ N_XI0/XI39/XI7/NET35_XI0/XI39/XI7/MM7_g N_VSS_XI0/XI39/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM8 N_XI0/XI39/XI7/NET35_XI0/XI39/XI7/MM8_d
+ N_WL<75>_XI0/XI39/XI7/MM8_g N_BLN<8>_XI0/XI39/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI7/MM5 N_XI0/XI39/XI7/NET34_XI0/XI39/XI7/MM5_d
+ N_XI0/XI39/XI7/NET33_XI0/XI39/XI7/MM5_g N_VDD_XI0/XI39/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI7/MM4 N_XI0/XI39/XI7/NET33_XI0/XI39/XI7/MM4_d
+ N_XI0/XI39/XI7/NET34_XI0/XI39/XI7/MM4_g N_VDD_XI0/XI39/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI7/MM10 N_XI0/XI39/XI7/NET35_XI0/XI39/XI7/MM10_d
+ N_XI0/XI39/XI7/NET36_XI0/XI39/XI7/MM10_g N_VDD_XI0/XI39/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI7/MM11 N_XI0/XI39/XI7/NET36_XI0/XI39/XI7/MM11_d
+ N_XI0/XI39/XI7/NET35_XI0/XI39/XI7/MM11_g N_VDD_XI0/XI39/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI8/MM2 N_XI0/XI39/XI8/NET34_XI0/XI39/XI8/MM2_d
+ N_XI0/XI39/XI8/NET33_XI0/XI39/XI8/MM2_g N_VSS_XI0/XI39/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM3 N_XI0/XI39/XI8/NET33_XI0/XI39/XI8/MM3_d
+ N_WL<74>_XI0/XI39/XI8/MM3_g N_BLN<7>_XI0/XI39/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM0 N_XI0/XI39/XI8/NET34_XI0/XI39/XI8/MM0_d
+ N_WL<74>_XI0/XI39/XI8/MM0_g N_BL<7>_XI0/XI39/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM1 N_XI0/XI39/XI8/NET33_XI0/XI39/XI8/MM1_d
+ N_XI0/XI39/XI8/NET34_XI0/XI39/XI8/MM1_g N_VSS_XI0/XI39/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM9 N_XI0/XI39/XI8/NET36_XI0/XI39/XI8/MM9_d
+ N_WL<75>_XI0/XI39/XI8/MM9_g N_BL<7>_XI0/XI39/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM6 N_XI0/XI39/XI8/NET35_XI0/XI39/XI8/MM6_d
+ N_XI0/XI39/XI8/NET36_XI0/XI39/XI8/MM6_g N_VSS_XI0/XI39/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM7 N_XI0/XI39/XI8/NET36_XI0/XI39/XI8/MM7_d
+ N_XI0/XI39/XI8/NET35_XI0/XI39/XI8/MM7_g N_VSS_XI0/XI39/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM8 N_XI0/XI39/XI8/NET35_XI0/XI39/XI8/MM8_d
+ N_WL<75>_XI0/XI39/XI8/MM8_g N_BLN<7>_XI0/XI39/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI8/MM5 N_XI0/XI39/XI8/NET34_XI0/XI39/XI8/MM5_d
+ N_XI0/XI39/XI8/NET33_XI0/XI39/XI8/MM5_g N_VDD_XI0/XI39/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI8/MM4 N_XI0/XI39/XI8/NET33_XI0/XI39/XI8/MM4_d
+ N_XI0/XI39/XI8/NET34_XI0/XI39/XI8/MM4_g N_VDD_XI0/XI39/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI8/MM10 N_XI0/XI39/XI8/NET35_XI0/XI39/XI8/MM10_d
+ N_XI0/XI39/XI8/NET36_XI0/XI39/XI8/MM10_g N_VDD_XI0/XI39/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI8/MM11 N_XI0/XI39/XI8/NET36_XI0/XI39/XI8/MM11_d
+ N_XI0/XI39/XI8/NET35_XI0/XI39/XI8/MM11_g N_VDD_XI0/XI39/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI9/MM2 N_XI0/XI39/XI9/NET34_XI0/XI39/XI9/MM2_d
+ N_XI0/XI39/XI9/NET33_XI0/XI39/XI9/MM2_g N_VSS_XI0/XI39/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM3 N_XI0/XI39/XI9/NET33_XI0/XI39/XI9/MM3_d
+ N_WL<74>_XI0/XI39/XI9/MM3_g N_BLN<6>_XI0/XI39/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM0 N_XI0/XI39/XI9/NET34_XI0/XI39/XI9/MM0_d
+ N_WL<74>_XI0/XI39/XI9/MM0_g N_BL<6>_XI0/XI39/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM1 N_XI0/XI39/XI9/NET33_XI0/XI39/XI9/MM1_d
+ N_XI0/XI39/XI9/NET34_XI0/XI39/XI9/MM1_g N_VSS_XI0/XI39/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM9 N_XI0/XI39/XI9/NET36_XI0/XI39/XI9/MM9_d
+ N_WL<75>_XI0/XI39/XI9/MM9_g N_BL<6>_XI0/XI39/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM6 N_XI0/XI39/XI9/NET35_XI0/XI39/XI9/MM6_d
+ N_XI0/XI39/XI9/NET36_XI0/XI39/XI9/MM6_g N_VSS_XI0/XI39/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM7 N_XI0/XI39/XI9/NET36_XI0/XI39/XI9/MM7_d
+ N_XI0/XI39/XI9/NET35_XI0/XI39/XI9/MM7_g N_VSS_XI0/XI39/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM8 N_XI0/XI39/XI9/NET35_XI0/XI39/XI9/MM8_d
+ N_WL<75>_XI0/XI39/XI9/MM8_g N_BLN<6>_XI0/XI39/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI9/MM5 N_XI0/XI39/XI9/NET34_XI0/XI39/XI9/MM5_d
+ N_XI0/XI39/XI9/NET33_XI0/XI39/XI9/MM5_g N_VDD_XI0/XI39/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI9/MM4 N_XI0/XI39/XI9/NET33_XI0/XI39/XI9/MM4_d
+ N_XI0/XI39/XI9/NET34_XI0/XI39/XI9/MM4_g N_VDD_XI0/XI39/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI9/MM10 N_XI0/XI39/XI9/NET35_XI0/XI39/XI9/MM10_d
+ N_XI0/XI39/XI9/NET36_XI0/XI39/XI9/MM10_g N_VDD_XI0/XI39/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI9/MM11 N_XI0/XI39/XI9/NET36_XI0/XI39/XI9/MM11_d
+ N_XI0/XI39/XI9/NET35_XI0/XI39/XI9/MM11_g N_VDD_XI0/XI39/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI10/MM2 N_XI0/XI39/XI10/NET34_XI0/XI39/XI10/MM2_d
+ N_XI0/XI39/XI10/NET33_XI0/XI39/XI10/MM2_g N_VSS_XI0/XI39/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM3 N_XI0/XI39/XI10/NET33_XI0/XI39/XI10/MM3_d
+ N_WL<74>_XI0/XI39/XI10/MM3_g N_BLN<5>_XI0/XI39/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM0 N_XI0/XI39/XI10/NET34_XI0/XI39/XI10/MM0_d
+ N_WL<74>_XI0/XI39/XI10/MM0_g N_BL<5>_XI0/XI39/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM1 N_XI0/XI39/XI10/NET33_XI0/XI39/XI10/MM1_d
+ N_XI0/XI39/XI10/NET34_XI0/XI39/XI10/MM1_g N_VSS_XI0/XI39/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM9 N_XI0/XI39/XI10/NET36_XI0/XI39/XI10/MM9_d
+ N_WL<75>_XI0/XI39/XI10/MM9_g N_BL<5>_XI0/XI39/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM6 N_XI0/XI39/XI10/NET35_XI0/XI39/XI10/MM6_d
+ N_XI0/XI39/XI10/NET36_XI0/XI39/XI10/MM6_g N_VSS_XI0/XI39/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM7 N_XI0/XI39/XI10/NET36_XI0/XI39/XI10/MM7_d
+ N_XI0/XI39/XI10/NET35_XI0/XI39/XI10/MM7_g N_VSS_XI0/XI39/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM8 N_XI0/XI39/XI10/NET35_XI0/XI39/XI10/MM8_d
+ N_WL<75>_XI0/XI39/XI10/MM8_g N_BLN<5>_XI0/XI39/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI10/MM5 N_XI0/XI39/XI10/NET34_XI0/XI39/XI10/MM5_d
+ N_XI0/XI39/XI10/NET33_XI0/XI39/XI10/MM5_g N_VDD_XI0/XI39/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI10/MM4 N_XI0/XI39/XI10/NET33_XI0/XI39/XI10/MM4_d
+ N_XI0/XI39/XI10/NET34_XI0/XI39/XI10/MM4_g N_VDD_XI0/XI39/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI10/MM10 N_XI0/XI39/XI10/NET35_XI0/XI39/XI10/MM10_d
+ N_XI0/XI39/XI10/NET36_XI0/XI39/XI10/MM10_g N_VDD_XI0/XI39/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI10/MM11 N_XI0/XI39/XI10/NET36_XI0/XI39/XI10/MM11_d
+ N_XI0/XI39/XI10/NET35_XI0/XI39/XI10/MM11_g N_VDD_XI0/XI39/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI11/MM2 N_XI0/XI39/XI11/NET34_XI0/XI39/XI11/MM2_d
+ N_XI0/XI39/XI11/NET33_XI0/XI39/XI11/MM2_g N_VSS_XI0/XI39/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM3 N_XI0/XI39/XI11/NET33_XI0/XI39/XI11/MM3_d
+ N_WL<74>_XI0/XI39/XI11/MM3_g N_BLN<4>_XI0/XI39/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM0 N_XI0/XI39/XI11/NET34_XI0/XI39/XI11/MM0_d
+ N_WL<74>_XI0/XI39/XI11/MM0_g N_BL<4>_XI0/XI39/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM1 N_XI0/XI39/XI11/NET33_XI0/XI39/XI11/MM1_d
+ N_XI0/XI39/XI11/NET34_XI0/XI39/XI11/MM1_g N_VSS_XI0/XI39/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM9 N_XI0/XI39/XI11/NET36_XI0/XI39/XI11/MM9_d
+ N_WL<75>_XI0/XI39/XI11/MM9_g N_BL<4>_XI0/XI39/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM6 N_XI0/XI39/XI11/NET35_XI0/XI39/XI11/MM6_d
+ N_XI0/XI39/XI11/NET36_XI0/XI39/XI11/MM6_g N_VSS_XI0/XI39/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM7 N_XI0/XI39/XI11/NET36_XI0/XI39/XI11/MM7_d
+ N_XI0/XI39/XI11/NET35_XI0/XI39/XI11/MM7_g N_VSS_XI0/XI39/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM8 N_XI0/XI39/XI11/NET35_XI0/XI39/XI11/MM8_d
+ N_WL<75>_XI0/XI39/XI11/MM8_g N_BLN<4>_XI0/XI39/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI11/MM5 N_XI0/XI39/XI11/NET34_XI0/XI39/XI11/MM5_d
+ N_XI0/XI39/XI11/NET33_XI0/XI39/XI11/MM5_g N_VDD_XI0/XI39/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI11/MM4 N_XI0/XI39/XI11/NET33_XI0/XI39/XI11/MM4_d
+ N_XI0/XI39/XI11/NET34_XI0/XI39/XI11/MM4_g N_VDD_XI0/XI39/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI11/MM10 N_XI0/XI39/XI11/NET35_XI0/XI39/XI11/MM10_d
+ N_XI0/XI39/XI11/NET36_XI0/XI39/XI11/MM10_g N_VDD_XI0/XI39/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI11/MM11 N_XI0/XI39/XI11/NET36_XI0/XI39/XI11/MM11_d
+ N_XI0/XI39/XI11/NET35_XI0/XI39/XI11/MM11_g N_VDD_XI0/XI39/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI12/MM2 N_XI0/XI39/XI12/NET34_XI0/XI39/XI12/MM2_d
+ N_XI0/XI39/XI12/NET33_XI0/XI39/XI12/MM2_g N_VSS_XI0/XI39/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM3 N_XI0/XI39/XI12/NET33_XI0/XI39/XI12/MM3_d
+ N_WL<74>_XI0/XI39/XI12/MM3_g N_BLN<3>_XI0/XI39/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM0 N_XI0/XI39/XI12/NET34_XI0/XI39/XI12/MM0_d
+ N_WL<74>_XI0/XI39/XI12/MM0_g N_BL<3>_XI0/XI39/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM1 N_XI0/XI39/XI12/NET33_XI0/XI39/XI12/MM1_d
+ N_XI0/XI39/XI12/NET34_XI0/XI39/XI12/MM1_g N_VSS_XI0/XI39/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM9 N_XI0/XI39/XI12/NET36_XI0/XI39/XI12/MM9_d
+ N_WL<75>_XI0/XI39/XI12/MM9_g N_BL<3>_XI0/XI39/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM6 N_XI0/XI39/XI12/NET35_XI0/XI39/XI12/MM6_d
+ N_XI0/XI39/XI12/NET36_XI0/XI39/XI12/MM6_g N_VSS_XI0/XI39/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM7 N_XI0/XI39/XI12/NET36_XI0/XI39/XI12/MM7_d
+ N_XI0/XI39/XI12/NET35_XI0/XI39/XI12/MM7_g N_VSS_XI0/XI39/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM8 N_XI0/XI39/XI12/NET35_XI0/XI39/XI12/MM8_d
+ N_WL<75>_XI0/XI39/XI12/MM8_g N_BLN<3>_XI0/XI39/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI12/MM5 N_XI0/XI39/XI12/NET34_XI0/XI39/XI12/MM5_d
+ N_XI0/XI39/XI12/NET33_XI0/XI39/XI12/MM5_g N_VDD_XI0/XI39/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI12/MM4 N_XI0/XI39/XI12/NET33_XI0/XI39/XI12/MM4_d
+ N_XI0/XI39/XI12/NET34_XI0/XI39/XI12/MM4_g N_VDD_XI0/XI39/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI12/MM10 N_XI0/XI39/XI12/NET35_XI0/XI39/XI12/MM10_d
+ N_XI0/XI39/XI12/NET36_XI0/XI39/XI12/MM10_g N_VDD_XI0/XI39/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI12/MM11 N_XI0/XI39/XI12/NET36_XI0/XI39/XI12/MM11_d
+ N_XI0/XI39/XI12/NET35_XI0/XI39/XI12/MM11_g N_VDD_XI0/XI39/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI13/MM2 N_XI0/XI39/XI13/NET34_XI0/XI39/XI13/MM2_d
+ N_XI0/XI39/XI13/NET33_XI0/XI39/XI13/MM2_g N_VSS_XI0/XI39/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM3 N_XI0/XI39/XI13/NET33_XI0/XI39/XI13/MM3_d
+ N_WL<74>_XI0/XI39/XI13/MM3_g N_BLN<2>_XI0/XI39/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM0 N_XI0/XI39/XI13/NET34_XI0/XI39/XI13/MM0_d
+ N_WL<74>_XI0/XI39/XI13/MM0_g N_BL<2>_XI0/XI39/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM1 N_XI0/XI39/XI13/NET33_XI0/XI39/XI13/MM1_d
+ N_XI0/XI39/XI13/NET34_XI0/XI39/XI13/MM1_g N_VSS_XI0/XI39/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM9 N_XI0/XI39/XI13/NET36_XI0/XI39/XI13/MM9_d
+ N_WL<75>_XI0/XI39/XI13/MM9_g N_BL<2>_XI0/XI39/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM6 N_XI0/XI39/XI13/NET35_XI0/XI39/XI13/MM6_d
+ N_XI0/XI39/XI13/NET36_XI0/XI39/XI13/MM6_g N_VSS_XI0/XI39/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM7 N_XI0/XI39/XI13/NET36_XI0/XI39/XI13/MM7_d
+ N_XI0/XI39/XI13/NET35_XI0/XI39/XI13/MM7_g N_VSS_XI0/XI39/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM8 N_XI0/XI39/XI13/NET35_XI0/XI39/XI13/MM8_d
+ N_WL<75>_XI0/XI39/XI13/MM8_g N_BLN<2>_XI0/XI39/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI13/MM5 N_XI0/XI39/XI13/NET34_XI0/XI39/XI13/MM5_d
+ N_XI0/XI39/XI13/NET33_XI0/XI39/XI13/MM5_g N_VDD_XI0/XI39/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI13/MM4 N_XI0/XI39/XI13/NET33_XI0/XI39/XI13/MM4_d
+ N_XI0/XI39/XI13/NET34_XI0/XI39/XI13/MM4_g N_VDD_XI0/XI39/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI13/MM10 N_XI0/XI39/XI13/NET35_XI0/XI39/XI13/MM10_d
+ N_XI0/XI39/XI13/NET36_XI0/XI39/XI13/MM10_g N_VDD_XI0/XI39/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI13/MM11 N_XI0/XI39/XI13/NET36_XI0/XI39/XI13/MM11_d
+ N_XI0/XI39/XI13/NET35_XI0/XI39/XI13/MM11_g N_VDD_XI0/XI39/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI14/MM2 N_XI0/XI39/XI14/NET34_XI0/XI39/XI14/MM2_d
+ N_XI0/XI39/XI14/NET33_XI0/XI39/XI14/MM2_g N_VSS_XI0/XI39/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM3 N_XI0/XI39/XI14/NET33_XI0/XI39/XI14/MM3_d
+ N_WL<74>_XI0/XI39/XI14/MM3_g N_BLN<1>_XI0/XI39/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM0 N_XI0/XI39/XI14/NET34_XI0/XI39/XI14/MM0_d
+ N_WL<74>_XI0/XI39/XI14/MM0_g N_BL<1>_XI0/XI39/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM1 N_XI0/XI39/XI14/NET33_XI0/XI39/XI14/MM1_d
+ N_XI0/XI39/XI14/NET34_XI0/XI39/XI14/MM1_g N_VSS_XI0/XI39/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM9 N_XI0/XI39/XI14/NET36_XI0/XI39/XI14/MM9_d
+ N_WL<75>_XI0/XI39/XI14/MM9_g N_BL<1>_XI0/XI39/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM6 N_XI0/XI39/XI14/NET35_XI0/XI39/XI14/MM6_d
+ N_XI0/XI39/XI14/NET36_XI0/XI39/XI14/MM6_g N_VSS_XI0/XI39/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM7 N_XI0/XI39/XI14/NET36_XI0/XI39/XI14/MM7_d
+ N_XI0/XI39/XI14/NET35_XI0/XI39/XI14/MM7_g N_VSS_XI0/XI39/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM8 N_XI0/XI39/XI14/NET35_XI0/XI39/XI14/MM8_d
+ N_WL<75>_XI0/XI39/XI14/MM8_g N_BLN<1>_XI0/XI39/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI14/MM5 N_XI0/XI39/XI14/NET34_XI0/XI39/XI14/MM5_d
+ N_XI0/XI39/XI14/NET33_XI0/XI39/XI14/MM5_g N_VDD_XI0/XI39/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI14/MM4 N_XI0/XI39/XI14/NET33_XI0/XI39/XI14/MM4_d
+ N_XI0/XI39/XI14/NET34_XI0/XI39/XI14/MM4_g N_VDD_XI0/XI39/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI14/MM10 N_XI0/XI39/XI14/NET35_XI0/XI39/XI14/MM10_d
+ N_XI0/XI39/XI14/NET36_XI0/XI39/XI14/MM10_g N_VDD_XI0/XI39/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI14/MM11 N_XI0/XI39/XI14/NET36_XI0/XI39/XI14/MM11_d
+ N_XI0/XI39/XI14/NET35_XI0/XI39/XI14/MM11_g N_VDD_XI0/XI39/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI15/MM2 N_XI0/XI39/XI15/NET34_XI0/XI39/XI15/MM2_d
+ N_XI0/XI39/XI15/NET33_XI0/XI39/XI15/MM2_g N_VSS_XI0/XI39/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM3 N_XI0/XI39/XI15/NET33_XI0/XI39/XI15/MM3_d
+ N_WL<74>_XI0/XI39/XI15/MM3_g N_BLN<0>_XI0/XI39/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM0 N_XI0/XI39/XI15/NET34_XI0/XI39/XI15/MM0_d
+ N_WL<74>_XI0/XI39/XI15/MM0_g N_BL<0>_XI0/XI39/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM1 N_XI0/XI39/XI15/NET33_XI0/XI39/XI15/MM1_d
+ N_XI0/XI39/XI15/NET34_XI0/XI39/XI15/MM1_g N_VSS_XI0/XI39/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM9 N_XI0/XI39/XI15/NET36_XI0/XI39/XI15/MM9_d
+ N_WL<75>_XI0/XI39/XI15/MM9_g N_BL<0>_XI0/XI39/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM6 N_XI0/XI39/XI15/NET35_XI0/XI39/XI15/MM6_d
+ N_XI0/XI39/XI15/NET36_XI0/XI39/XI15/MM6_g N_VSS_XI0/XI39/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM7 N_XI0/XI39/XI15/NET36_XI0/XI39/XI15/MM7_d
+ N_XI0/XI39/XI15/NET35_XI0/XI39/XI15/MM7_g N_VSS_XI0/XI39/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM8 N_XI0/XI39/XI15/NET35_XI0/XI39/XI15/MM8_d
+ N_WL<75>_XI0/XI39/XI15/MM8_g N_BLN<0>_XI0/XI39/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI39/XI15/MM5 N_XI0/XI39/XI15/NET34_XI0/XI39/XI15/MM5_d
+ N_XI0/XI39/XI15/NET33_XI0/XI39/XI15/MM5_g N_VDD_XI0/XI39/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI15/MM4 N_XI0/XI39/XI15/NET33_XI0/XI39/XI15/MM4_d
+ N_XI0/XI39/XI15/NET34_XI0/XI39/XI15/MM4_g N_VDD_XI0/XI39/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI15/MM10 N_XI0/XI39/XI15/NET35_XI0/XI39/XI15/MM10_d
+ N_XI0/XI39/XI15/NET36_XI0/XI39/XI15/MM10_g N_VDD_XI0/XI39/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI39/XI15/MM11 N_XI0/XI39/XI15/NET36_XI0/XI39/XI15/MM11_d
+ N_XI0/XI39/XI15/NET35_XI0/XI39/XI15/MM11_g N_VDD_XI0/XI39/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI0/MM2 N_XI0/XI40/XI0/NET34_XI0/XI40/XI0/MM2_d
+ N_XI0/XI40/XI0/NET33_XI0/XI40/XI0/MM2_g N_VSS_XI0/XI40/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM3 N_XI0/XI40/XI0/NET33_XI0/XI40/XI0/MM3_d
+ N_WL<76>_XI0/XI40/XI0/MM3_g N_BLN<15>_XI0/XI40/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM0 N_XI0/XI40/XI0/NET34_XI0/XI40/XI0/MM0_d
+ N_WL<76>_XI0/XI40/XI0/MM0_g N_BL<15>_XI0/XI40/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM1 N_XI0/XI40/XI0/NET33_XI0/XI40/XI0/MM1_d
+ N_XI0/XI40/XI0/NET34_XI0/XI40/XI0/MM1_g N_VSS_XI0/XI40/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM9 N_XI0/XI40/XI0/NET36_XI0/XI40/XI0/MM9_d
+ N_WL<77>_XI0/XI40/XI0/MM9_g N_BL<15>_XI0/XI40/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM6 N_XI0/XI40/XI0/NET35_XI0/XI40/XI0/MM6_d
+ N_XI0/XI40/XI0/NET36_XI0/XI40/XI0/MM6_g N_VSS_XI0/XI40/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM7 N_XI0/XI40/XI0/NET36_XI0/XI40/XI0/MM7_d
+ N_XI0/XI40/XI0/NET35_XI0/XI40/XI0/MM7_g N_VSS_XI0/XI40/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM8 N_XI0/XI40/XI0/NET35_XI0/XI40/XI0/MM8_d
+ N_WL<77>_XI0/XI40/XI0/MM8_g N_BLN<15>_XI0/XI40/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI0/MM5 N_XI0/XI40/XI0/NET34_XI0/XI40/XI0/MM5_d
+ N_XI0/XI40/XI0/NET33_XI0/XI40/XI0/MM5_g N_VDD_XI0/XI40/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI0/MM4 N_XI0/XI40/XI0/NET33_XI0/XI40/XI0/MM4_d
+ N_XI0/XI40/XI0/NET34_XI0/XI40/XI0/MM4_g N_VDD_XI0/XI40/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI0/MM10 N_XI0/XI40/XI0/NET35_XI0/XI40/XI0/MM10_d
+ N_XI0/XI40/XI0/NET36_XI0/XI40/XI0/MM10_g N_VDD_XI0/XI40/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI0/MM11 N_XI0/XI40/XI0/NET36_XI0/XI40/XI0/MM11_d
+ N_XI0/XI40/XI0/NET35_XI0/XI40/XI0/MM11_g N_VDD_XI0/XI40/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI1/MM2 N_XI0/XI40/XI1/NET34_XI0/XI40/XI1/MM2_d
+ N_XI0/XI40/XI1/NET33_XI0/XI40/XI1/MM2_g N_VSS_XI0/XI40/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM3 N_XI0/XI40/XI1/NET33_XI0/XI40/XI1/MM3_d
+ N_WL<76>_XI0/XI40/XI1/MM3_g N_BLN<14>_XI0/XI40/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM0 N_XI0/XI40/XI1/NET34_XI0/XI40/XI1/MM0_d
+ N_WL<76>_XI0/XI40/XI1/MM0_g N_BL<14>_XI0/XI40/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM1 N_XI0/XI40/XI1/NET33_XI0/XI40/XI1/MM1_d
+ N_XI0/XI40/XI1/NET34_XI0/XI40/XI1/MM1_g N_VSS_XI0/XI40/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM9 N_XI0/XI40/XI1/NET36_XI0/XI40/XI1/MM9_d
+ N_WL<77>_XI0/XI40/XI1/MM9_g N_BL<14>_XI0/XI40/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM6 N_XI0/XI40/XI1/NET35_XI0/XI40/XI1/MM6_d
+ N_XI0/XI40/XI1/NET36_XI0/XI40/XI1/MM6_g N_VSS_XI0/XI40/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM7 N_XI0/XI40/XI1/NET36_XI0/XI40/XI1/MM7_d
+ N_XI0/XI40/XI1/NET35_XI0/XI40/XI1/MM7_g N_VSS_XI0/XI40/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM8 N_XI0/XI40/XI1/NET35_XI0/XI40/XI1/MM8_d
+ N_WL<77>_XI0/XI40/XI1/MM8_g N_BLN<14>_XI0/XI40/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI1/MM5 N_XI0/XI40/XI1/NET34_XI0/XI40/XI1/MM5_d
+ N_XI0/XI40/XI1/NET33_XI0/XI40/XI1/MM5_g N_VDD_XI0/XI40/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI1/MM4 N_XI0/XI40/XI1/NET33_XI0/XI40/XI1/MM4_d
+ N_XI0/XI40/XI1/NET34_XI0/XI40/XI1/MM4_g N_VDD_XI0/XI40/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI1/MM10 N_XI0/XI40/XI1/NET35_XI0/XI40/XI1/MM10_d
+ N_XI0/XI40/XI1/NET36_XI0/XI40/XI1/MM10_g N_VDD_XI0/XI40/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI1/MM11 N_XI0/XI40/XI1/NET36_XI0/XI40/XI1/MM11_d
+ N_XI0/XI40/XI1/NET35_XI0/XI40/XI1/MM11_g N_VDD_XI0/XI40/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI2/MM2 N_XI0/XI40/XI2/NET34_XI0/XI40/XI2/MM2_d
+ N_XI0/XI40/XI2/NET33_XI0/XI40/XI2/MM2_g N_VSS_XI0/XI40/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM3 N_XI0/XI40/XI2/NET33_XI0/XI40/XI2/MM3_d
+ N_WL<76>_XI0/XI40/XI2/MM3_g N_BLN<13>_XI0/XI40/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM0 N_XI0/XI40/XI2/NET34_XI0/XI40/XI2/MM0_d
+ N_WL<76>_XI0/XI40/XI2/MM0_g N_BL<13>_XI0/XI40/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM1 N_XI0/XI40/XI2/NET33_XI0/XI40/XI2/MM1_d
+ N_XI0/XI40/XI2/NET34_XI0/XI40/XI2/MM1_g N_VSS_XI0/XI40/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM9 N_XI0/XI40/XI2/NET36_XI0/XI40/XI2/MM9_d
+ N_WL<77>_XI0/XI40/XI2/MM9_g N_BL<13>_XI0/XI40/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM6 N_XI0/XI40/XI2/NET35_XI0/XI40/XI2/MM6_d
+ N_XI0/XI40/XI2/NET36_XI0/XI40/XI2/MM6_g N_VSS_XI0/XI40/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM7 N_XI0/XI40/XI2/NET36_XI0/XI40/XI2/MM7_d
+ N_XI0/XI40/XI2/NET35_XI0/XI40/XI2/MM7_g N_VSS_XI0/XI40/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM8 N_XI0/XI40/XI2/NET35_XI0/XI40/XI2/MM8_d
+ N_WL<77>_XI0/XI40/XI2/MM8_g N_BLN<13>_XI0/XI40/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI2/MM5 N_XI0/XI40/XI2/NET34_XI0/XI40/XI2/MM5_d
+ N_XI0/XI40/XI2/NET33_XI0/XI40/XI2/MM5_g N_VDD_XI0/XI40/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI2/MM4 N_XI0/XI40/XI2/NET33_XI0/XI40/XI2/MM4_d
+ N_XI0/XI40/XI2/NET34_XI0/XI40/XI2/MM4_g N_VDD_XI0/XI40/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI2/MM10 N_XI0/XI40/XI2/NET35_XI0/XI40/XI2/MM10_d
+ N_XI0/XI40/XI2/NET36_XI0/XI40/XI2/MM10_g N_VDD_XI0/XI40/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI2/MM11 N_XI0/XI40/XI2/NET36_XI0/XI40/XI2/MM11_d
+ N_XI0/XI40/XI2/NET35_XI0/XI40/XI2/MM11_g N_VDD_XI0/XI40/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI3/MM2 N_XI0/XI40/XI3/NET34_XI0/XI40/XI3/MM2_d
+ N_XI0/XI40/XI3/NET33_XI0/XI40/XI3/MM2_g N_VSS_XI0/XI40/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM3 N_XI0/XI40/XI3/NET33_XI0/XI40/XI3/MM3_d
+ N_WL<76>_XI0/XI40/XI3/MM3_g N_BLN<12>_XI0/XI40/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM0 N_XI0/XI40/XI3/NET34_XI0/XI40/XI3/MM0_d
+ N_WL<76>_XI0/XI40/XI3/MM0_g N_BL<12>_XI0/XI40/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM1 N_XI0/XI40/XI3/NET33_XI0/XI40/XI3/MM1_d
+ N_XI0/XI40/XI3/NET34_XI0/XI40/XI3/MM1_g N_VSS_XI0/XI40/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM9 N_XI0/XI40/XI3/NET36_XI0/XI40/XI3/MM9_d
+ N_WL<77>_XI0/XI40/XI3/MM9_g N_BL<12>_XI0/XI40/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM6 N_XI0/XI40/XI3/NET35_XI0/XI40/XI3/MM6_d
+ N_XI0/XI40/XI3/NET36_XI0/XI40/XI3/MM6_g N_VSS_XI0/XI40/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM7 N_XI0/XI40/XI3/NET36_XI0/XI40/XI3/MM7_d
+ N_XI0/XI40/XI3/NET35_XI0/XI40/XI3/MM7_g N_VSS_XI0/XI40/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM8 N_XI0/XI40/XI3/NET35_XI0/XI40/XI3/MM8_d
+ N_WL<77>_XI0/XI40/XI3/MM8_g N_BLN<12>_XI0/XI40/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI3/MM5 N_XI0/XI40/XI3/NET34_XI0/XI40/XI3/MM5_d
+ N_XI0/XI40/XI3/NET33_XI0/XI40/XI3/MM5_g N_VDD_XI0/XI40/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI3/MM4 N_XI0/XI40/XI3/NET33_XI0/XI40/XI3/MM4_d
+ N_XI0/XI40/XI3/NET34_XI0/XI40/XI3/MM4_g N_VDD_XI0/XI40/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI3/MM10 N_XI0/XI40/XI3/NET35_XI0/XI40/XI3/MM10_d
+ N_XI0/XI40/XI3/NET36_XI0/XI40/XI3/MM10_g N_VDD_XI0/XI40/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI3/MM11 N_XI0/XI40/XI3/NET36_XI0/XI40/XI3/MM11_d
+ N_XI0/XI40/XI3/NET35_XI0/XI40/XI3/MM11_g N_VDD_XI0/XI40/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI4/MM2 N_XI0/XI40/XI4/NET34_XI0/XI40/XI4/MM2_d
+ N_XI0/XI40/XI4/NET33_XI0/XI40/XI4/MM2_g N_VSS_XI0/XI40/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM3 N_XI0/XI40/XI4/NET33_XI0/XI40/XI4/MM3_d
+ N_WL<76>_XI0/XI40/XI4/MM3_g N_BLN<11>_XI0/XI40/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM0 N_XI0/XI40/XI4/NET34_XI0/XI40/XI4/MM0_d
+ N_WL<76>_XI0/XI40/XI4/MM0_g N_BL<11>_XI0/XI40/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM1 N_XI0/XI40/XI4/NET33_XI0/XI40/XI4/MM1_d
+ N_XI0/XI40/XI4/NET34_XI0/XI40/XI4/MM1_g N_VSS_XI0/XI40/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM9 N_XI0/XI40/XI4/NET36_XI0/XI40/XI4/MM9_d
+ N_WL<77>_XI0/XI40/XI4/MM9_g N_BL<11>_XI0/XI40/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM6 N_XI0/XI40/XI4/NET35_XI0/XI40/XI4/MM6_d
+ N_XI0/XI40/XI4/NET36_XI0/XI40/XI4/MM6_g N_VSS_XI0/XI40/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM7 N_XI0/XI40/XI4/NET36_XI0/XI40/XI4/MM7_d
+ N_XI0/XI40/XI4/NET35_XI0/XI40/XI4/MM7_g N_VSS_XI0/XI40/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM8 N_XI0/XI40/XI4/NET35_XI0/XI40/XI4/MM8_d
+ N_WL<77>_XI0/XI40/XI4/MM8_g N_BLN<11>_XI0/XI40/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI4/MM5 N_XI0/XI40/XI4/NET34_XI0/XI40/XI4/MM5_d
+ N_XI0/XI40/XI4/NET33_XI0/XI40/XI4/MM5_g N_VDD_XI0/XI40/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI4/MM4 N_XI0/XI40/XI4/NET33_XI0/XI40/XI4/MM4_d
+ N_XI0/XI40/XI4/NET34_XI0/XI40/XI4/MM4_g N_VDD_XI0/XI40/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI4/MM10 N_XI0/XI40/XI4/NET35_XI0/XI40/XI4/MM10_d
+ N_XI0/XI40/XI4/NET36_XI0/XI40/XI4/MM10_g N_VDD_XI0/XI40/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI4/MM11 N_XI0/XI40/XI4/NET36_XI0/XI40/XI4/MM11_d
+ N_XI0/XI40/XI4/NET35_XI0/XI40/XI4/MM11_g N_VDD_XI0/XI40/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI5/MM2 N_XI0/XI40/XI5/NET34_XI0/XI40/XI5/MM2_d
+ N_XI0/XI40/XI5/NET33_XI0/XI40/XI5/MM2_g N_VSS_XI0/XI40/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM3 N_XI0/XI40/XI5/NET33_XI0/XI40/XI5/MM3_d
+ N_WL<76>_XI0/XI40/XI5/MM3_g N_BLN<10>_XI0/XI40/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM0 N_XI0/XI40/XI5/NET34_XI0/XI40/XI5/MM0_d
+ N_WL<76>_XI0/XI40/XI5/MM0_g N_BL<10>_XI0/XI40/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM1 N_XI0/XI40/XI5/NET33_XI0/XI40/XI5/MM1_d
+ N_XI0/XI40/XI5/NET34_XI0/XI40/XI5/MM1_g N_VSS_XI0/XI40/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM9 N_XI0/XI40/XI5/NET36_XI0/XI40/XI5/MM9_d
+ N_WL<77>_XI0/XI40/XI5/MM9_g N_BL<10>_XI0/XI40/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM6 N_XI0/XI40/XI5/NET35_XI0/XI40/XI5/MM6_d
+ N_XI0/XI40/XI5/NET36_XI0/XI40/XI5/MM6_g N_VSS_XI0/XI40/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM7 N_XI0/XI40/XI5/NET36_XI0/XI40/XI5/MM7_d
+ N_XI0/XI40/XI5/NET35_XI0/XI40/XI5/MM7_g N_VSS_XI0/XI40/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM8 N_XI0/XI40/XI5/NET35_XI0/XI40/XI5/MM8_d
+ N_WL<77>_XI0/XI40/XI5/MM8_g N_BLN<10>_XI0/XI40/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI5/MM5 N_XI0/XI40/XI5/NET34_XI0/XI40/XI5/MM5_d
+ N_XI0/XI40/XI5/NET33_XI0/XI40/XI5/MM5_g N_VDD_XI0/XI40/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI5/MM4 N_XI0/XI40/XI5/NET33_XI0/XI40/XI5/MM4_d
+ N_XI0/XI40/XI5/NET34_XI0/XI40/XI5/MM4_g N_VDD_XI0/XI40/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI5/MM10 N_XI0/XI40/XI5/NET35_XI0/XI40/XI5/MM10_d
+ N_XI0/XI40/XI5/NET36_XI0/XI40/XI5/MM10_g N_VDD_XI0/XI40/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI5/MM11 N_XI0/XI40/XI5/NET36_XI0/XI40/XI5/MM11_d
+ N_XI0/XI40/XI5/NET35_XI0/XI40/XI5/MM11_g N_VDD_XI0/XI40/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI6/MM2 N_XI0/XI40/XI6/NET34_XI0/XI40/XI6/MM2_d
+ N_XI0/XI40/XI6/NET33_XI0/XI40/XI6/MM2_g N_VSS_XI0/XI40/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM3 N_XI0/XI40/XI6/NET33_XI0/XI40/XI6/MM3_d
+ N_WL<76>_XI0/XI40/XI6/MM3_g N_BLN<9>_XI0/XI40/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM0 N_XI0/XI40/XI6/NET34_XI0/XI40/XI6/MM0_d
+ N_WL<76>_XI0/XI40/XI6/MM0_g N_BL<9>_XI0/XI40/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM1 N_XI0/XI40/XI6/NET33_XI0/XI40/XI6/MM1_d
+ N_XI0/XI40/XI6/NET34_XI0/XI40/XI6/MM1_g N_VSS_XI0/XI40/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM9 N_XI0/XI40/XI6/NET36_XI0/XI40/XI6/MM9_d
+ N_WL<77>_XI0/XI40/XI6/MM9_g N_BL<9>_XI0/XI40/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM6 N_XI0/XI40/XI6/NET35_XI0/XI40/XI6/MM6_d
+ N_XI0/XI40/XI6/NET36_XI0/XI40/XI6/MM6_g N_VSS_XI0/XI40/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM7 N_XI0/XI40/XI6/NET36_XI0/XI40/XI6/MM7_d
+ N_XI0/XI40/XI6/NET35_XI0/XI40/XI6/MM7_g N_VSS_XI0/XI40/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM8 N_XI0/XI40/XI6/NET35_XI0/XI40/XI6/MM8_d
+ N_WL<77>_XI0/XI40/XI6/MM8_g N_BLN<9>_XI0/XI40/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI6/MM5 N_XI0/XI40/XI6/NET34_XI0/XI40/XI6/MM5_d
+ N_XI0/XI40/XI6/NET33_XI0/XI40/XI6/MM5_g N_VDD_XI0/XI40/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI6/MM4 N_XI0/XI40/XI6/NET33_XI0/XI40/XI6/MM4_d
+ N_XI0/XI40/XI6/NET34_XI0/XI40/XI6/MM4_g N_VDD_XI0/XI40/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI6/MM10 N_XI0/XI40/XI6/NET35_XI0/XI40/XI6/MM10_d
+ N_XI0/XI40/XI6/NET36_XI0/XI40/XI6/MM10_g N_VDD_XI0/XI40/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI6/MM11 N_XI0/XI40/XI6/NET36_XI0/XI40/XI6/MM11_d
+ N_XI0/XI40/XI6/NET35_XI0/XI40/XI6/MM11_g N_VDD_XI0/XI40/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI7/MM2 N_XI0/XI40/XI7/NET34_XI0/XI40/XI7/MM2_d
+ N_XI0/XI40/XI7/NET33_XI0/XI40/XI7/MM2_g N_VSS_XI0/XI40/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM3 N_XI0/XI40/XI7/NET33_XI0/XI40/XI7/MM3_d
+ N_WL<76>_XI0/XI40/XI7/MM3_g N_BLN<8>_XI0/XI40/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM0 N_XI0/XI40/XI7/NET34_XI0/XI40/XI7/MM0_d
+ N_WL<76>_XI0/XI40/XI7/MM0_g N_BL<8>_XI0/XI40/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM1 N_XI0/XI40/XI7/NET33_XI0/XI40/XI7/MM1_d
+ N_XI0/XI40/XI7/NET34_XI0/XI40/XI7/MM1_g N_VSS_XI0/XI40/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM9 N_XI0/XI40/XI7/NET36_XI0/XI40/XI7/MM9_d
+ N_WL<77>_XI0/XI40/XI7/MM9_g N_BL<8>_XI0/XI40/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM6 N_XI0/XI40/XI7/NET35_XI0/XI40/XI7/MM6_d
+ N_XI0/XI40/XI7/NET36_XI0/XI40/XI7/MM6_g N_VSS_XI0/XI40/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM7 N_XI0/XI40/XI7/NET36_XI0/XI40/XI7/MM7_d
+ N_XI0/XI40/XI7/NET35_XI0/XI40/XI7/MM7_g N_VSS_XI0/XI40/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM8 N_XI0/XI40/XI7/NET35_XI0/XI40/XI7/MM8_d
+ N_WL<77>_XI0/XI40/XI7/MM8_g N_BLN<8>_XI0/XI40/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI7/MM5 N_XI0/XI40/XI7/NET34_XI0/XI40/XI7/MM5_d
+ N_XI0/XI40/XI7/NET33_XI0/XI40/XI7/MM5_g N_VDD_XI0/XI40/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI7/MM4 N_XI0/XI40/XI7/NET33_XI0/XI40/XI7/MM4_d
+ N_XI0/XI40/XI7/NET34_XI0/XI40/XI7/MM4_g N_VDD_XI0/XI40/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI7/MM10 N_XI0/XI40/XI7/NET35_XI0/XI40/XI7/MM10_d
+ N_XI0/XI40/XI7/NET36_XI0/XI40/XI7/MM10_g N_VDD_XI0/XI40/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI7/MM11 N_XI0/XI40/XI7/NET36_XI0/XI40/XI7/MM11_d
+ N_XI0/XI40/XI7/NET35_XI0/XI40/XI7/MM11_g N_VDD_XI0/XI40/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI8/MM2 N_XI0/XI40/XI8/NET34_XI0/XI40/XI8/MM2_d
+ N_XI0/XI40/XI8/NET33_XI0/XI40/XI8/MM2_g N_VSS_XI0/XI40/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM3 N_XI0/XI40/XI8/NET33_XI0/XI40/XI8/MM3_d
+ N_WL<76>_XI0/XI40/XI8/MM3_g N_BLN<7>_XI0/XI40/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM0 N_XI0/XI40/XI8/NET34_XI0/XI40/XI8/MM0_d
+ N_WL<76>_XI0/XI40/XI8/MM0_g N_BL<7>_XI0/XI40/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM1 N_XI0/XI40/XI8/NET33_XI0/XI40/XI8/MM1_d
+ N_XI0/XI40/XI8/NET34_XI0/XI40/XI8/MM1_g N_VSS_XI0/XI40/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM9 N_XI0/XI40/XI8/NET36_XI0/XI40/XI8/MM9_d
+ N_WL<77>_XI0/XI40/XI8/MM9_g N_BL<7>_XI0/XI40/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM6 N_XI0/XI40/XI8/NET35_XI0/XI40/XI8/MM6_d
+ N_XI0/XI40/XI8/NET36_XI0/XI40/XI8/MM6_g N_VSS_XI0/XI40/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM7 N_XI0/XI40/XI8/NET36_XI0/XI40/XI8/MM7_d
+ N_XI0/XI40/XI8/NET35_XI0/XI40/XI8/MM7_g N_VSS_XI0/XI40/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM8 N_XI0/XI40/XI8/NET35_XI0/XI40/XI8/MM8_d
+ N_WL<77>_XI0/XI40/XI8/MM8_g N_BLN<7>_XI0/XI40/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI8/MM5 N_XI0/XI40/XI8/NET34_XI0/XI40/XI8/MM5_d
+ N_XI0/XI40/XI8/NET33_XI0/XI40/XI8/MM5_g N_VDD_XI0/XI40/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI8/MM4 N_XI0/XI40/XI8/NET33_XI0/XI40/XI8/MM4_d
+ N_XI0/XI40/XI8/NET34_XI0/XI40/XI8/MM4_g N_VDD_XI0/XI40/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI8/MM10 N_XI0/XI40/XI8/NET35_XI0/XI40/XI8/MM10_d
+ N_XI0/XI40/XI8/NET36_XI0/XI40/XI8/MM10_g N_VDD_XI0/XI40/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI8/MM11 N_XI0/XI40/XI8/NET36_XI0/XI40/XI8/MM11_d
+ N_XI0/XI40/XI8/NET35_XI0/XI40/XI8/MM11_g N_VDD_XI0/XI40/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI9/MM2 N_XI0/XI40/XI9/NET34_XI0/XI40/XI9/MM2_d
+ N_XI0/XI40/XI9/NET33_XI0/XI40/XI9/MM2_g N_VSS_XI0/XI40/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM3 N_XI0/XI40/XI9/NET33_XI0/XI40/XI9/MM3_d
+ N_WL<76>_XI0/XI40/XI9/MM3_g N_BLN<6>_XI0/XI40/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM0 N_XI0/XI40/XI9/NET34_XI0/XI40/XI9/MM0_d
+ N_WL<76>_XI0/XI40/XI9/MM0_g N_BL<6>_XI0/XI40/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM1 N_XI0/XI40/XI9/NET33_XI0/XI40/XI9/MM1_d
+ N_XI0/XI40/XI9/NET34_XI0/XI40/XI9/MM1_g N_VSS_XI0/XI40/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM9 N_XI0/XI40/XI9/NET36_XI0/XI40/XI9/MM9_d
+ N_WL<77>_XI0/XI40/XI9/MM9_g N_BL<6>_XI0/XI40/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM6 N_XI0/XI40/XI9/NET35_XI0/XI40/XI9/MM6_d
+ N_XI0/XI40/XI9/NET36_XI0/XI40/XI9/MM6_g N_VSS_XI0/XI40/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM7 N_XI0/XI40/XI9/NET36_XI0/XI40/XI9/MM7_d
+ N_XI0/XI40/XI9/NET35_XI0/XI40/XI9/MM7_g N_VSS_XI0/XI40/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM8 N_XI0/XI40/XI9/NET35_XI0/XI40/XI9/MM8_d
+ N_WL<77>_XI0/XI40/XI9/MM8_g N_BLN<6>_XI0/XI40/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI9/MM5 N_XI0/XI40/XI9/NET34_XI0/XI40/XI9/MM5_d
+ N_XI0/XI40/XI9/NET33_XI0/XI40/XI9/MM5_g N_VDD_XI0/XI40/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI9/MM4 N_XI0/XI40/XI9/NET33_XI0/XI40/XI9/MM4_d
+ N_XI0/XI40/XI9/NET34_XI0/XI40/XI9/MM4_g N_VDD_XI0/XI40/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI9/MM10 N_XI0/XI40/XI9/NET35_XI0/XI40/XI9/MM10_d
+ N_XI0/XI40/XI9/NET36_XI0/XI40/XI9/MM10_g N_VDD_XI0/XI40/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI9/MM11 N_XI0/XI40/XI9/NET36_XI0/XI40/XI9/MM11_d
+ N_XI0/XI40/XI9/NET35_XI0/XI40/XI9/MM11_g N_VDD_XI0/XI40/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI10/MM2 N_XI0/XI40/XI10/NET34_XI0/XI40/XI10/MM2_d
+ N_XI0/XI40/XI10/NET33_XI0/XI40/XI10/MM2_g N_VSS_XI0/XI40/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM3 N_XI0/XI40/XI10/NET33_XI0/XI40/XI10/MM3_d
+ N_WL<76>_XI0/XI40/XI10/MM3_g N_BLN<5>_XI0/XI40/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM0 N_XI0/XI40/XI10/NET34_XI0/XI40/XI10/MM0_d
+ N_WL<76>_XI0/XI40/XI10/MM0_g N_BL<5>_XI0/XI40/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM1 N_XI0/XI40/XI10/NET33_XI0/XI40/XI10/MM1_d
+ N_XI0/XI40/XI10/NET34_XI0/XI40/XI10/MM1_g N_VSS_XI0/XI40/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM9 N_XI0/XI40/XI10/NET36_XI0/XI40/XI10/MM9_d
+ N_WL<77>_XI0/XI40/XI10/MM9_g N_BL<5>_XI0/XI40/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM6 N_XI0/XI40/XI10/NET35_XI0/XI40/XI10/MM6_d
+ N_XI0/XI40/XI10/NET36_XI0/XI40/XI10/MM6_g N_VSS_XI0/XI40/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM7 N_XI0/XI40/XI10/NET36_XI0/XI40/XI10/MM7_d
+ N_XI0/XI40/XI10/NET35_XI0/XI40/XI10/MM7_g N_VSS_XI0/XI40/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM8 N_XI0/XI40/XI10/NET35_XI0/XI40/XI10/MM8_d
+ N_WL<77>_XI0/XI40/XI10/MM8_g N_BLN<5>_XI0/XI40/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI10/MM5 N_XI0/XI40/XI10/NET34_XI0/XI40/XI10/MM5_d
+ N_XI0/XI40/XI10/NET33_XI0/XI40/XI10/MM5_g N_VDD_XI0/XI40/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI10/MM4 N_XI0/XI40/XI10/NET33_XI0/XI40/XI10/MM4_d
+ N_XI0/XI40/XI10/NET34_XI0/XI40/XI10/MM4_g N_VDD_XI0/XI40/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI10/MM10 N_XI0/XI40/XI10/NET35_XI0/XI40/XI10/MM10_d
+ N_XI0/XI40/XI10/NET36_XI0/XI40/XI10/MM10_g N_VDD_XI0/XI40/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI10/MM11 N_XI0/XI40/XI10/NET36_XI0/XI40/XI10/MM11_d
+ N_XI0/XI40/XI10/NET35_XI0/XI40/XI10/MM11_g N_VDD_XI0/XI40/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI11/MM2 N_XI0/XI40/XI11/NET34_XI0/XI40/XI11/MM2_d
+ N_XI0/XI40/XI11/NET33_XI0/XI40/XI11/MM2_g N_VSS_XI0/XI40/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM3 N_XI0/XI40/XI11/NET33_XI0/XI40/XI11/MM3_d
+ N_WL<76>_XI0/XI40/XI11/MM3_g N_BLN<4>_XI0/XI40/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM0 N_XI0/XI40/XI11/NET34_XI0/XI40/XI11/MM0_d
+ N_WL<76>_XI0/XI40/XI11/MM0_g N_BL<4>_XI0/XI40/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM1 N_XI0/XI40/XI11/NET33_XI0/XI40/XI11/MM1_d
+ N_XI0/XI40/XI11/NET34_XI0/XI40/XI11/MM1_g N_VSS_XI0/XI40/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM9 N_XI0/XI40/XI11/NET36_XI0/XI40/XI11/MM9_d
+ N_WL<77>_XI0/XI40/XI11/MM9_g N_BL<4>_XI0/XI40/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM6 N_XI0/XI40/XI11/NET35_XI0/XI40/XI11/MM6_d
+ N_XI0/XI40/XI11/NET36_XI0/XI40/XI11/MM6_g N_VSS_XI0/XI40/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM7 N_XI0/XI40/XI11/NET36_XI0/XI40/XI11/MM7_d
+ N_XI0/XI40/XI11/NET35_XI0/XI40/XI11/MM7_g N_VSS_XI0/XI40/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM8 N_XI0/XI40/XI11/NET35_XI0/XI40/XI11/MM8_d
+ N_WL<77>_XI0/XI40/XI11/MM8_g N_BLN<4>_XI0/XI40/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI11/MM5 N_XI0/XI40/XI11/NET34_XI0/XI40/XI11/MM5_d
+ N_XI0/XI40/XI11/NET33_XI0/XI40/XI11/MM5_g N_VDD_XI0/XI40/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI11/MM4 N_XI0/XI40/XI11/NET33_XI0/XI40/XI11/MM4_d
+ N_XI0/XI40/XI11/NET34_XI0/XI40/XI11/MM4_g N_VDD_XI0/XI40/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI11/MM10 N_XI0/XI40/XI11/NET35_XI0/XI40/XI11/MM10_d
+ N_XI0/XI40/XI11/NET36_XI0/XI40/XI11/MM10_g N_VDD_XI0/XI40/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI11/MM11 N_XI0/XI40/XI11/NET36_XI0/XI40/XI11/MM11_d
+ N_XI0/XI40/XI11/NET35_XI0/XI40/XI11/MM11_g N_VDD_XI0/XI40/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI12/MM2 N_XI0/XI40/XI12/NET34_XI0/XI40/XI12/MM2_d
+ N_XI0/XI40/XI12/NET33_XI0/XI40/XI12/MM2_g N_VSS_XI0/XI40/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM3 N_XI0/XI40/XI12/NET33_XI0/XI40/XI12/MM3_d
+ N_WL<76>_XI0/XI40/XI12/MM3_g N_BLN<3>_XI0/XI40/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM0 N_XI0/XI40/XI12/NET34_XI0/XI40/XI12/MM0_d
+ N_WL<76>_XI0/XI40/XI12/MM0_g N_BL<3>_XI0/XI40/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM1 N_XI0/XI40/XI12/NET33_XI0/XI40/XI12/MM1_d
+ N_XI0/XI40/XI12/NET34_XI0/XI40/XI12/MM1_g N_VSS_XI0/XI40/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM9 N_XI0/XI40/XI12/NET36_XI0/XI40/XI12/MM9_d
+ N_WL<77>_XI0/XI40/XI12/MM9_g N_BL<3>_XI0/XI40/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM6 N_XI0/XI40/XI12/NET35_XI0/XI40/XI12/MM6_d
+ N_XI0/XI40/XI12/NET36_XI0/XI40/XI12/MM6_g N_VSS_XI0/XI40/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM7 N_XI0/XI40/XI12/NET36_XI0/XI40/XI12/MM7_d
+ N_XI0/XI40/XI12/NET35_XI0/XI40/XI12/MM7_g N_VSS_XI0/XI40/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM8 N_XI0/XI40/XI12/NET35_XI0/XI40/XI12/MM8_d
+ N_WL<77>_XI0/XI40/XI12/MM8_g N_BLN<3>_XI0/XI40/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI12/MM5 N_XI0/XI40/XI12/NET34_XI0/XI40/XI12/MM5_d
+ N_XI0/XI40/XI12/NET33_XI0/XI40/XI12/MM5_g N_VDD_XI0/XI40/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI12/MM4 N_XI0/XI40/XI12/NET33_XI0/XI40/XI12/MM4_d
+ N_XI0/XI40/XI12/NET34_XI0/XI40/XI12/MM4_g N_VDD_XI0/XI40/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI12/MM10 N_XI0/XI40/XI12/NET35_XI0/XI40/XI12/MM10_d
+ N_XI0/XI40/XI12/NET36_XI0/XI40/XI12/MM10_g N_VDD_XI0/XI40/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI12/MM11 N_XI0/XI40/XI12/NET36_XI0/XI40/XI12/MM11_d
+ N_XI0/XI40/XI12/NET35_XI0/XI40/XI12/MM11_g N_VDD_XI0/XI40/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI13/MM2 N_XI0/XI40/XI13/NET34_XI0/XI40/XI13/MM2_d
+ N_XI0/XI40/XI13/NET33_XI0/XI40/XI13/MM2_g N_VSS_XI0/XI40/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM3 N_XI0/XI40/XI13/NET33_XI0/XI40/XI13/MM3_d
+ N_WL<76>_XI0/XI40/XI13/MM3_g N_BLN<2>_XI0/XI40/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM0 N_XI0/XI40/XI13/NET34_XI0/XI40/XI13/MM0_d
+ N_WL<76>_XI0/XI40/XI13/MM0_g N_BL<2>_XI0/XI40/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM1 N_XI0/XI40/XI13/NET33_XI0/XI40/XI13/MM1_d
+ N_XI0/XI40/XI13/NET34_XI0/XI40/XI13/MM1_g N_VSS_XI0/XI40/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM9 N_XI0/XI40/XI13/NET36_XI0/XI40/XI13/MM9_d
+ N_WL<77>_XI0/XI40/XI13/MM9_g N_BL<2>_XI0/XI40/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM6 N_XI0/XI40/XI13/NET35_XI0/XI40/XI13/MM6_d
+ N_XI0/XI40/XI13/NET36_XI0/XI40/XI13/MM6_g N_VSS_XI0/XI40/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM7 N_XI0/XI40/XI13/NET36_XI0/XI40/XI13/MM7_d
+ N_XI0/XI40/XI13/NET35_XI0/XI40/XI13/MM7_g N_VSS_XI0/XI40/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM8 N_XI0/XI40/XI13/NET35_XI0/XI40/XI13/MM8_d
+ N_WL<77>_XI0/XI40/XI13/MM8_g N_BLN<2>_XI0/XI40/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI13/MM5 N_XI0/XI40/XI13/NET34_XI0/XI40/XI13/MM5_d
+ N_XI0/XI40/XI13/NET33_XI0/XI40/XI13/MM5_g N_VDD_XI0/XI40/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI13/MM4 N_XI0/XI40/XI13/NET33_XI0/XI40/XI13/MM4_d
+ N_XI0/XI40/XI13/NET34_XI0/XI40/XI13/MM4_g N_VDD_XI0/XI40/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI13/MM10 N_XI0/XI40/XI13/NET35_XI0/XI40/XI13/MM10_d
+ N_XI0/XI40/XI13/NET36_XI0/XI40/XI13/MM10_g N_VDD_XI0/XI40/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI13/MM11 N_XI0/XI40/XI13/NET36_XI0/XI40/XI13/MM11_d
+ N_XI0/XI40/XI13/NET35_XI0/XI40/XI13/MM11_g N_VDD_XI0/XI40/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI14/MM2 N_XI0/XI40/XI14/NET34_XI0/XI40/XI14/MM2_d
+ N_XI0/XI40/XI14/NET33_XI0/XI40/XI14/MM2_g N_VSS_XI0/XI40/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM3 N_XI0/XI40/XI14/NET33_XI0/XI40/XI14/MM3_d
+ N_WL<76>_XI0/XI40/XI14/MM3_g N_BLN<1>_XI0/XI40/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM0 N_XI0/XI40/XI14/NET34_XI0/XI40/XI14/MM0_d
+ N_WL<76>_XI0/XI40/XI14/MM0_g N_BL<1>_XI0/XI40/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM1 N_XI0/XI40/XI14/NET33_XI0/XI40/XI14/MM1_d
+ N_XI0/XI40/XI14/NET34_XI0/XI40/XI14/MM1_g N_VSS_XI0/XI40/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM9 N_XI0/XI40/XI14/NET36_XI0/XI40/XI14/MM9_d
+ N_WL<77>_XI0/XI40/XI14/MM9_g N_BL<1>_XI0/XI40/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM6 N_XI0/XI40/XI14/NET35_XI0/XI40/XI14/MM6_d
+ N_XI0/XI40/XI14/NET36_XI0/XI40/XI14/MM6_g N_VSS_XI0/XI40/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM7 N_XI0/XI40/XI14/NET36_XI0/XI40/XI14/MM7_d
+ N_XI0/XI40/XI14/NET35_XI0/XI40/XI14/MM7_g N_VSS_XI0/XI40/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM8 N_XI0/XI40/XI14/NET35_XI0/XI40/XI14/MM8_d
+ N_WL<77>_XI0/XI40/XI14/MM8_g N_BLN<1>_XI0/XI40/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI14/MM5 N_XI0/XI40/XI14/NET34_XI0/XI40/XI14/MM5_d
+ N_XI0/XI40/XI14/NET33_XI0/XI40/XI14/MM5_g N_VDD_XI0/XI40/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI14/MM4 N_XI0/XI40/XI14/NET33_XI0/XI40/XI14/MM4_d
+ N_XI0/XI40/XI14/NET34_XI0/XI40/XI14/MM4_g N_VDD_XI0/XI40/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI14/MM10 N_XI0/XI40/XI14/NET35_XI0/XI40/XI14/MM10_d
+ N_XI0/XI40/XI14/NET36_XI0/XI40/XI14/MM10_g N_VDD_XI0/XI40/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI14/MM11 N_XI0/XI40/XI14/NET36_XI0/XI40/XI14/MM11_d
+ N_XI0/XI40/XI14/NET35_XI0/XI40/XI14/MM11_g N_VDD_XI0/XI40/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI15/MM2 N_XI0/XI40/XI15/NET34_XI0/XI40/XI15/MM2_d
+ N_XI0/XI40/XI15/NET33_XI0/XI40/XI15/MM2_g N_VSS_XI0/XI40/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM3 N_XI0/XI40/XI15/NET33_XI0/XI40/XI15/MM3_d
+ N_WL<76>_XI0/XI40/XI15/MM3_g N_BLN<0>_XI0/XI40/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM0 N_XI0/XI40/XI15/NET34_XI0/XI40/XI15/MM0_d
+ N_WL<76>_XI0/XI40/XI15/MM0_g N_BL<0>_XI0/XI40/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM1 N_XI0/XI40/XI15/NET33_XI0/XI40/XI15/MM1_d
+ N_XI0/XI40/XI15/NET34_XI0/XI40/XI15/MM1_g N_VSS_XI0/XI40/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM9 N_XI0/XI40/XI15/NET36_XI0/XI40/XI15/MM9_d
+ N_WL<77>_XI0/XI40/XI15/MM9_g N_BL<0>_XI0/XI40/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM6 N_XI0/XI40/XI15/NET35_XI0/XI40/XI15/MM6_d
+ N_XI0/XI40/XI15/NET36_XI0/XI40/XI15/MM6_g N_VSS_XI0/XI40/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM7 N_XI0/XI40/XI15/NET36_XI0/XI40/XI15/MM7_d
+ N_XI0/XI40/XI15/NET35_XI0/XI40/XI15/MM7_g N_VSS_XI0/XI40/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM8 N_XI0/XI40/XI15/NET35_XI0/XI40/XI15/MM8_d
+ N_WL<77>_XI0/XI40/XI15/MM8_g N_BLN<0>_XI0/XI40/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI40/XI15/MM5 N_XI0/XI40/XI15/NET34_XI0/XI40/XI15/MM5_d
+ N_XI0/XI40/XI15/NET33_XI0/XI40/XI15/MM5_g N_VDD_XI0/XI40/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI15/MM4 N_XI0/XI40/XI15/NET33_XI0/XI40/XI15/MM4_d
+ N_XI0/XI40/XI15/NET34_XI0/XI40/XI15/MM4_g N_VDD_XI0/XI40/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI15/MM10 N_XI0/XI40/XI15/NET35_XI0/XI40/XI15/MM10_d
+ N_XI0/XI40/XI15/NET36_XI0/XI40/XI15/MM10_g N_VDD_XI0/XI40/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI40/XI15/MM11 N_XI0/XI40/XI15/NET36_XI0/XI40/XI15/MM11_d
+ N_XI0/XI40/XI15/NET35_XI0/XI40/XI15/MM11_g N_VDD_XI0/XI40/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI0/MM2 N_XI0/XI41/XI0/NET34_XI0/XI41/XI0/MM2_d
+ N_XI0/XI41/XI0/NET33_XI0/XI41/XI0/MM2_g N_VSS_XI0/XI41/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM3 N_XI0/XI41/XI0/NET33_XI0/XI41/XI0/MM3_d
+ N_WL<78>_XI0/XI41/XI0/MM3_g N_BLN<15>_XI0/XI41/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM0 N_XI0/XI41/XI0/NET34_XI0/XI41/XI0/MM0_d
+ N_WL<78>_XI0/XI41/XI0/MM0_g N_BL<15>_XI0/XI41/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM1 N_XI0/XI41/XI0/NET33_XI0/XI41/XI0/MM1_d
+ N_XI0/XI41/XI0/NET34_XI0/XI41/XI0/MM1_g N_VSS_XI0/XI41/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM9 N_XI0/XI41/XI0/NET36_XI0/XI41/XI0/MM9_d
+ N_WL<79>_XI0/XI41/XI0/MM9_g N_BL<15>_XI0/XI41/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM6 N_XI0/XI41/XI0/NET35_XI0/XI41/XI0/MM6_d
+ N_XI0/XI41/XI0/NET36_XI0/XI41/XI0/MM6_g N_VSS_XI0/XI41/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM7 N_XI0/XI41/XI0/NET36_XI0/XI41/XI0/MM7_d
+ N_XI0/XI41/XI0/NET35_XI0/XI41/XI0/MM7_g N_VSS_XI0/XI41/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM8 N_XI0/XI41/XI0/NET35_XI0/XI41/XI0/MM8_d
+ N_WL<79>_XI0/XI41/XI0/MM8_g N_BLN<15>_XI0/XI41/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI0/MM5 N_XI0/XI41/XI0/NET34_XI0/XI41/XI0/MM5_d
+ N_XI0/XI41/XI0/NET33_XI0/XI41/XI0/MM5_g N_VDD_XI0/XI41/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI0/MM4 N_XI0/XI41/XI0/NET33_XI0/XI41/XI0/MM4_d
+ N_XI0/XI41/XI0/NET34_XI0/XI41/XI0/MM4_g N_VDD_XI0/XI41/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI0/MM10 N_XI0/XI41/XI0/NET35_XI0/XI41/XI0/MM10_d
+ N_XI0/XI41/XI0/NET36_XI0/XI41/XI0/MM10_g N_VDD_XI0/XI41/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI0/MM11 N_XI0/XI41/XI0/NET36_XI0/XI41/XI0/MM11_d
+ N_XI0/XI41/XI0/NET35_XI0/XI41/XI0/MM11_g N_VDD_XI0/XI41/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI1/MM2 N_XI0/XI41/XI1/NET34_XI0/XI41/XI1/MM2_d
+ N_XI0/XI41/XI1/NET33_XI0/XI41/XI1/MM2_g N_VSS_XI0/XI41/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM3 N_XI0/XI41/XI1/NET33_XI0/XI41/XI1/MM3_d
+ N_WL<78>_XI0/XI41/XI1/MM3_g N_BLN<14>_XI0/XI41/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM0 N_XI0/XI41/XI1/NET34_XI0/XI41/XI1/MM0_d
+ N_WL<78>_XI0/XI41/XI1/MM0_g N_BL<14>_XI0/XI41/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM1 N_XI0/XI41/XI1/NET33_XI0/XI41/XI1/MM1_d
+ N_XI0/XI41/XI1/NET34_XI0/XI41/XI1/MM1_g N_VSS_XI0/XI41/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM9 N_XI0/XI41/XI1/NET36_XI0/XI41/XI1/MM9_d
+ N_WL<79>_XI0/XI41/XI1/MM9_g N_BL<14>_XI0/XI41/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM6 N_XI0/XI41/XI1/NET35_XI0/XI41/XI1/MM6_d
+ N_XI0/XI41/XI1/NET36_XI0/XI41/XI1/MM6_g N_VSS_XI0/XI41/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM7 N_XI0/XI41/XI1/NET36_XI0/XI41/XI1/MM7_d
+ N_XI0/XI41/XI1/NET35_XI0/XI41/XI1/MM7_g N_VSS_XI0/XI41/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM8 N_XI0/XI41/XI1/NET35_XI0/XI41/XI1/MM8_d
+ N_WL<79>_XI0/XI41/XI1/MM8_g N_BLN<14>_XI0/XI41/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI1/MM5 N_XI0/XI41/XI1/NET34_XI0/XI41/XI1/MM5_d
+ N_XI0/XI41/XI1/NET33_XI0/XI41/XI1/MM5_g N_VDD_XI0/XI41/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI1/MM4 N_XI0/XI41/XI1/NET33_XI0/XI41/XI1/MM4_d
+ N_XI0/XI41/XI1/NET34_XI0/XI41/XI1/MM4_g N_VDD_XI0/XI41/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI1/MM10 N_XI0/XI41/XI1/NET35_XI0/XI41/XI1/MM10_d
+ N_XI0/XI41/XI1/NET36_XI0/XI41/XI1/MM10_g N_VDD_XI0/XI41/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI1/MM11 N_XI0/XI41/XI1/NET36_XI0/XI41/XI1/MM11_d
+ N_XI0/XI41/XI1/NET35_XI0/XI41/XI1/MM11_g N_VDD_XI0/XI41/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI2/MM2 N_XI0/XI41/XI2/NET34_XI0/XI41/XI2/MM2_d
+ N_XI0/XI41/XI2/NET33_XI0/XI41/XI2/MM2_g N_VSS_XI0/XI41/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM3 N_XI0/XI41/XI2/NET33_XI0/XI41/XI2/MM3_d
+ N_WL<78>_XI0/XI41/XI2/MM3_g N_BLN<13>_XI0/XI41/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM0 N_XI0/XI41/XI2/NET34_XI0/XI41/XI2/MM0_d
+ N_WL<78>_XI0/XI41/XI2/MM0_g N_BL<13>_XI0/XI41/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM1 N_XI0/XI41/XI2/NET33_XI0/XI41/XI2/MM1_d
+ N_XI0/XI41/XI2/NET34_XI0/XI41/XI2/MM1_g N_VSS_XI0/XI41/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM9 N_XI0/XI41/XI2/NET36_XI0/XI41/XI2/MM9_d
+ N_WL<79>_XI0/XI41/XI2/MM9_g N_BL<13>_XI0/XI41/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM6 N_XI0/XI41/XI2/NET35_XI0/XI41/XI2/MM6_d
+ N_XI0/XI41/XI2/NET36_XI0/XI41/XI2/MM6_g N_VSS_XI0/XI41/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM7 N_XI0/XI41/XI2/NET36_XI0/XI41/XI2/MM7_d
+ N_XI0/XI41/XI2/NET35_XI0/XI41/XI2/MM7_g N_VSS_XI0/XI41/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM8 N_XI0/XI41/XI2/NET35_XI0/XI41/XI2/MM8_d
+ N_WL<79>_XI0/XI41/XI2/MM8_g N_BLN<13>_XI0/XI41/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI2/MM5 N_XI0/XI41/XI2/NET34_XI0/XI41/XI2/MM5_d
+ N_XI0/XI41/XI2/NET33_XI0/XI41/XI2/MM5_g N_VDD_XI0/XI41/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI2/MM4 N_XI0/XI41/XI2/NET33_XI0/XI41/XI2/MM4_d
+ N_XI0/XI41/XI2/NET34_XI0/XI41/XI2/MM4_g N_VDD_XI0/XI41/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI2/MM10 N_XI0/XI41/XI2/NET35_XI0/XI41/XI2/MM10_d
+ N_XI0/XI41/XI2/NET36_XI0/XI41/XI2/MM10_g N_VDD_XI0/XI41/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI2/MM11 N_XI0/XI41/XI2/NET36_XI0/XI41/XI2/MM11_d
+ N_XI0/XI41/XI2/NET35_XI0/XI41/XI2/MM11_g N_VDD_XI0/XI41/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI3/MM2 N_XI0/XI41/XI3/NET34_XI0/XI41/XI3/MM2_d
+ N_XI0/XI41/XI3/NET33_XI0/XI41/XI3/MM2_g N_VSS_XI0/XI41/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM3 N_XI0/XI41/XI3/NET33_XI0/XI41/XI3/MM3_d
+ N_WL<78>_XI0/XI41/XI3/MM3_g N_BLN<12>_XI0/XI41/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM0 N_XI0/XI41/XI3/NET34_XI0/XI41/XI3/MM0_d
+ N_WL<78>_XI0/XI41/XI3/MM0_g N_BL<12>_XI0/XI41/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM1 N_XI0/XI41/XI3/NET33_XI0/XI41/XI3/MM1_d
+ N_XI0/XI41/XI3/NET34_XI0/XI41/XI3/MM1_g N_VSS_XI0/XI41/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM9 N_XI0/XI41/XI3/NET36_XI0/XI41/XI3/MM9_d
+ N_WL<79>_XI0/XI41/XI3/MM9_g N_BL<12>_XI0/XI41/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM6 N_XI0/XI41/XI3/NET35_XI0/XI41/XI3/MM6_d
+ N_XI0/XI41/XI3/NET36_XI0/XI41/XI3/MM6_g N_VSS_XI0/XI41/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM7 N_XI0/XI41/XI3/NET36_XI0/XI41/XI3/MM7_d
+ N_XI0/XI41/XI3/NET35_XI0/XI41/XI3/MM7_g N_VSS_XI0/XI41/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM8 N_XI0/XI41/XI3/NET35_XI0/XI41/XI3/MM8_d
+ N_WL<79>_XI0/XI41/XI3/MM8_g N_BLN<12>_XI0/XI41/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI3/MM5 N_XI0/XI41/XI3/NET34_XI0/XI41/XI3/MM5_d
+ N_XI0/XI41/XI3/NET33_XI0/XI41/XI3/MM5_g N_VDD_XI0/XI41/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI3/MM4 N_XI0/XI41/XI3/NET33_XI0/XI41/XI3/MM4_d
+ N_XI0/XI41/XI3/NET34_XI0/XI41/XI3/MM4_g N_VDD_XI0/XI41/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI3/MM10 N_XI0/XI41/XI3/NET35_XI0/XI41/XI3/MM10_d
+ N_XI0/XI41/XI3/NET36_XI0/XI41/XI3/MM10_g N_VDD_XI0/XI41/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI3/MM11 N_XI0/XI41/XI3/NET36_XI0/XI41/XI3/MM11_d
+ N_XI0/XI41/XI3/NET35_XI0/XI41/XI3/MM11_g N_VDD_XI0/XI41/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI4/MM2 N_XI0/XI41/XI4/NET34_XI0/XI41/XI4/MM2_d
+ N_XI0/XI41/XI4/NET33_XI0/XI41/XI4/MM2_g N_VSS_XI0/XI41/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM3 N_XI0/XI41/XI4/NET33_XI0/XI41/XI4/MM3_d
+ N_WL<78>_XI0/XI41/XI4/MM3_g N_BLN<11>_XI0/XI41/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM0 N_XI0/XI41/XI4/NET34_XI0/XI41/XI4/MM0_d
+ N_WL<78>_XI0/XI41/XI4/MM0_g N_BL<11>_XI0/XI41/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM1 N_XI0/XI41/XI4/NET33_XI0/XI41/XI4/MM1_d
+ N_XI0/XI41/XI4/NET34_XI0/XI41/XI4/MM1_g N_VSS_XI0/XI41/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM9 N_XI0/XI41/XI4/NET36_XI0/XI41/XI4/MM9_d
+ N_WL<79>_XI0/XI41/XI4/MM9_g N_BL<11>_XI0/XI41/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM6 N_XI0/XI41/XI4/NET35_XI0/XI41/XI4/MM6_d
+ N_XI0/XI41/XI4/NET36_XI0/XI41/XI4/MM6_g N_VSS_XI0/XI41/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM7 N_XI0/XI41/XI4/NET36_XI0/XI41/XI4/MM7_d
+ N_XI0/XI41/XI4/NET35_XI0/XI41/XI4/MM7_g N_VSS_XI0/XI41/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM8 N_XI0/XI41/XI4/NET35_XI0/XI41/XI4/MM8_d
+ N_WL<79>_XI0/XI41/XI4/MM8_g N_BLN<11>_XI0/XI41/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI4/MM5 N_XI0/XI41/XI4/NET34_XI0/XI41/XI4/MM5_d
+ N_XI0/XI41/XI4/NET33_XI0/XI41/XI4/MM5_g N_VDD_XI0/XI41/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI4/MM4 N_XI0/XI41/XI4/NET33_XI0/XI41/XI4/MM4_d
+ N_XI0/XI41/XI4/NET34_XI0/XI41/XI4/MM4_g N_VDD_XI0/XI41/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI4/MM10 N_XI0/XI41/XI4/NET35_XI0/XI41/XI4/MM10_d
+ N_XI0/XI41/XI4/NET36_XI0/XI41/XI4/MM10_g N_VDD_XI0/XI41/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI4/MM11 N_XI0/XI41/XI4/NET36_XI0/XI41/XI4/MM11_d
+ N_XI0/XI41/XI4/NET35_XI0/XI41/XI4/MM11_g N_VDD_XI0/XI41/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI5/MM2 N_XI0/XI41/XI5/NET34_XI0/XI41/XI5/MM2_d
+ N_XI0/XI41/XI5/NET33_XI0/XI41/XI5/MM2_g N_VSS_XI0/XI41/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM3 N_XI0/XI41/XI5/NET33_XI0/XI41/XI5/MM3_d
+ N_WL<78>_XI0/XI41/XI5/MM3_g N_BLN<10>_XI0/XI41/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM0 N_XI0/XI41/XI5/NET34_XI0/XI41/XI5/MM0_d
+ N_WL<78>_XI0/XI41/XI5/MM0_g N_BL<10>_XI0/XI41/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM1 N_XI0/XI41/XI5/NET33_XI0/XI41/XI5/MM1_d
+ N_XI0/XI41/XI5/NET34_XI0/XI41/XI5/MM1_g N_VSS_XI0/XI41/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM9 N_XI0/XI41/XI5/NET36_XI0/XI41/XI5/MM9_d
+ N_WL<79>_XI0/XI41/XI5/MM9_g N_BL<10>_XI0/XI41/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM6 N_XI0/XI41/XI5/NET35_XI0/XI41/XI5/MM6_d
+ N_XI0/XI41/XI5/NET36_XI0/XI41/XI5/MM6_g N_VSS_XI0/XI41/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM7 N_XI0/XI41/XI5/NET36_XI0/XI41/XI5/MM7_d
+ N_XI0/XI41/XI5/NET35_XI0/XI41/XI5/MM7_g N_VSS_XI0/XI41/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM8 N_XI0/XI41/XI5/NET35_XI0/XI41/XI5/MM8_d
+ N_WL<79>_XI0/XI41/XI5/MM8_g N_BLN<10>_XI0/XI41/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI5/MM5 N_XI0/XI41/XI5/NET34_XI0/XI41/XI5/MM5_d
+ N_XI0/XI41/XI5/NET33_XI0/XI41/XI5/MM5_g N_VDD_XI0/XI41/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI5/MM4 N_XI0/XI41/XI5/NET33_XI0/XI41/XI5/MM4_d
+ N_XI0/XI41/XI5/NET34_XI0/XI41/XI5/MM4_g N_VDD_XI0/XI41/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI5/MM10 N_XI0/XI41/XI5/NET35_XI0/XI41/XI5/MM10_d
+ N_XI0/XI41/XI5/NET36_XI0/XI41/XI5/MM10_g N_VDD_XI0/XI41/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI5/MM11 N_XI0/XI41/XI5/NET36_XI0/XI41/XI5/MM11_d
+ N_XI0/XI41/XI5/NET35_XI0/XI41/XI5/MM11_g N_VDD_XI0/XI41/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI6/MM2 N_XI0/XI41/XI6/NET34_XI0/XI41/XI6/MM2_d
+ N_XI0/XI41/XI6/NET33_XI0/XI41/XI6/MM2_g N_VSS_XI0/XI41/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM3 N_XI0/XI41/XI6/NET33_XI0/XI41/XI6/MM3_d
+ N_WL<78>_XI0/XI41/XI6/MM3_g N_BLN<9>_XI0/XI41/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM0 N_XI0/XI41/XI6/NET34_XI0/XI41/XI6/MM0_d
+ N_WL<78>_XI0/XI41/XI6/MM0_g N_BL<9>_XI0/XI41/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM1 N_XI0/XI41/XI6/NET33_XI0/XI41/XI6/MM1_d
+ N_XI0/XI41/XI6/NET34_XI0/XI41/XI6/MM1_g N_VSS_XI0/XI41/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM9 N_XI0/XI41/XI6/NET36_XI0/XI41/XI6/MM9_d
+ N_WL<79>_XI0/XI41/XI6/MM9_g N_BL<9>_XI0/XI41/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM6 N_XI0/XI41/XI6/NET35_XI0/XI41/XI6/MM6_d
+ N_XI0/XI41/XI6/NET36_XI0/XI41/XI6/MM6_g N_VSS_XI0/XI41/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM7 N_XI0/XI41/XI6/NET36_XI0/XI41/XI6/MM7_d
+ N_XI0/XI41/XI6/NET35_XI0/XI41/XI6/MM7_g N_VSS_XI0/XI41/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM8 N_XI0/XI41/XI6/NET35_XI0/XI41/XI6/MM8_d
+ N_WL<79>_XI0/XI41/XI6/MM8_g N_BLN<9>_XI0/XI41/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI6/MM5 N_XI0/XI41/XI6/NET34_XI0/XI41/XI6/MM5_d
+ N_XI0/XI41/XI6/NET33_XI0/XI41/XI6/MM5_g N_VDD_XI0/XI41/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI6/MM4 N_XI0/XI41/XI6/NET33_XI0/XI41/XI6/MM4_d
+ N_XI0/XI41/XI6/NET34_XI0/XI41/XI6/MM4_g N_VDD_XI0/XI41/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI6/MM10 N_XI0/XI41/XI6/NET35_XI0/XI41/XI6/MM10_d
+ N_XI0/XI41/XI6/NET36_XI0/XI41/XI6/MM10_g N_VDD_XI0/XI41/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI6/MM11 N_XI0/XI41/XI6/NET36_XI0/XI41/XI6/MM11_d
+ N_XI0/XI41/XI6/NET35_XI0/XI41/XI6/MM11_g N_VDD_XI0/XI41/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI7/MM2 N_XI0/XI41/XI7/NET34_XI0/XI41/XI7/MM2_d
+ N_XI0/XI41/XI7/NET33_XI0/XI41/XI7/MM2_g N_VSS_XI0/XI41/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM3 N_XI0/XI41/XI7/NET33_XI0/XI41/XI7/MM3_d
+ N_WL<78>_XI0/XI41/XI7/MM3_g N_BLN<8>_XI0/XI41/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM0 N_XI0/XI41/XI7/NET34_XI0/XI41/XI7/MM0_d
+ N_WL<78>_XI0/XI41/XI7/MM0_g N_BL<8>_XI0/XI41/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM1 N_XI0/XI41/XI7/NET33_XI0/XI41/XI7/MM1_d
+ N_XI0/XI41/XI7/NET34_XI0/XI41/XI7/MM1_g N_VSS_XI0/XI41/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM9 N_XI0/XI41/XI7/NET36_XI0/XI41/XI7/MM9_d
+ N_WL<79>_XI0/XI41/XI7/MM9_g N_BL<8>_XI0/XI41/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM6 N_XI0/XI41/XI7/NET35_XI0/XI41/XI7/MM6_d
+ N_XI0/XI41/XI7/NET36_XI0/XI41/XI7/MM6_g N_VSS_XI0/XI41/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM7 N_XI0/XI41/XI7/NET36_XI0/XI41/XI7/MM7_d
+ N_XI0/XI41/XI7/NET35_XI0/XI41/XI7/MM7_g N_VSS_XI0/XI41/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM8 N_XI0/XI41/XI7/NET35_XI0/XI41/XI7/MM8_d
+ N_WL<79>_XI0/XI41/XI7/MM8_g N_BLN<8>_XI0/XI41/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI7/MM5 N_XI0/XI41/XI7/NET34_XI0/XI41/XI7/MM5_d
+ N_XI0/XI41/XI7/NET33_XI0/XI41/XI7/MM5_g N_VDD_XI0/XI41/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI7/MM4 N_XI0/XI41/XI7/NET33_XI0/XI41/XI7/MM4_d
+ N_XI0/XI41/XI7/NET34_XI0/XI41/XI7/MM4_g N_VDD_XI0/XI41/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI7/MM10 N_XI0/XI41/XI7/NET35_XI0/XI41/XI7/MM10_d
+ N_XI0/XI41/XI7/NET36_XI0/XI41/XI7/MM10_g N_VDD_XI0/XI41/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI7/MM11 N_XI0/XI41/XI7/NET36_XI0/XI41/XI7/MM11_d
+ N_XI0/XI41/XI7/NET35_XI0/XI41/XI7/MM11_g N_VDD_XI0/XI41/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI8/MM2 N_XI0/XI41/XI8/NET34_XI0/XI41/XI8/MM2_d
+ N_XI0/XI41/XI8/NET33_XI0/XI41/XI8/MM2_g N_VSS_XI0/XI41/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM3 N_XI0/XI41/XI8/NET33_XI0/XI41/XI8/MM3_d
+ N_WL<78>_XI0/XI41/XI8/MM3_g N_BLN<7>_XI0/XI41/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM0 N_XI0/XI41/XI8/NET34_XI0/XI41/XI8/MM0_d
+ N_WL<78>_XI0/XI41/XI8/MM0_g N_BL<7>_XI0/XI41/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM1 N_XI0/XI41/XI8/NET33_XI0/XI41/XI8/MM1_d
+ N_XI0/XI41/XI8/NET34_XI0/XI41/XI8/MM1_g N_VSS_XI0/XI41/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM9 N_XI0/XI41/XI8/NET36_XI0/XI41/XI8/MM9_d
+ N_WL<79>_XI0/XI41/XI8/MM9_g N_BL<7>_XI0/XI41/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM6 N_XI0/XI41/XI8/NET35_XI0/XI41/XI8/MM6_d
+ N_XI0/XI41/XI8/NET36_XI0/XI41/XI8/MM6_g N_VSS_XI0/XI41/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM7 N_XI0/XI41/XI8/NET36_XI0/XI41/XI8/MM7_d
+ N_XI0/XI41/XI8/NET35_XI0/XI41/XI8/MM7_g N_VSS_XI0/XI41/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM8 N_XI0/XI41/XI8/NET35_XI0/XI41/XI8/MM8_d
+ N_WL<79>_XI0/XI41/XI8/MM8_g N_BLN<7>_XI0/XI41/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI8/MM5 N_XI0/XI41/XI8/NET34_XI0/XI41/XI8/MM5_d
+ N_XI0/XI41/XI8/NET33_XI0/XI41/XI8/MM5_g N_VDD_XI0/XI41/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI8/MM4 N_XI0/XI41/XI8/NET33_XI0/XI41/XI8/MM4_d
+ N_XI0/XI41/XI8/NET34_XI0/XI41/XI8/MM4_g N_VDD_XI0/XI41/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI8/MM10 N_XI0/XI41/XI8/NET35_XI0/XI41/XI8/MM10_d
+ N_XI0/XI41/XI8/NET36_XI0/XI41/XI8/MM10_g N_VDD_XI0/XI41/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI8/MM11 N_XI0/XI41/XI8/NET36_XI0/XI41/XI8/MM11_d
+ N_XI0/XI41/XI8/NET35_XI0/XI41/XI8/MM11_g N_VDD_XI0/XI41/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI9/MM2 N_XI0/XI41/XI9/NET34_XI0/XI41/XI9/MM2_d
+ N_XI0/XI41/XI9/NET33_XI0/XI41/XI9/MM2_g N_VSS_XI0/XI41/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM3 N_XI0/XI41/XI9/NET33_XI0/XI41/XI9/MM3_d
+ N_WL<78>_XI0/XI41/XI9/MM3_g N_BLN<6>_XI0/XI41/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM0 N_XI0/XI41/XI9/NET34_XI0/XI41/XI9/MM0_d
+ N_WL<78>_XI0/XI41/XI9/MM0_g N_BL<6>_XI0/XI41/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM1 N_XI0/XI41/XI9/NET33_XI0/XI41/XI9/MM1_d
+ N_XI0/XI41/XI9/NET34_XI0/XI41/XI9/MM1_g N_VSS_XI0/XI41/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM9 N_XI0/XI41/XI9/NET36_XI0/XI41/XI9/MM9_d
+ N_WL<79>_XI0/XI41/XI9/MM9_g N_BL<6>_XI0/XI41/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM6 N_XI0/XI41/XI9/NET35_XI0/XI41/XI9/MM6_d
+ N_XI0/XI41/XI9/NET36_XI0/XI41/XI9/MM6_g N_VSS_XI0/XI41/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM7 N_XI0/XI41/XI9/NET36_XI0/XI41/XI9/MM7_d
+ N_XI0/XI41/XI9/NET35_XI0/XI41/XI9/MM7_g N_VSS_XI0/XI41/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM8 N_XI0/XI41/XI9/NET35_XI0/XI41/XI9/MM8_d
+ N_WL<79>_XI0/XI41/XI9/MM8_g N_BLN<6>_XI0/XI41/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI9/MM5 N_XI0/XI41/XI9/NET34_XI0/XI41/XI9/MM5_d
+ N_XI0/XI41/XI9/NET33_XI0/XI41/XI9/MM5_g N_VDD_XI0/XI41/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI9/MM4 N_XI0/XI41/XI9/NET33_XI0/XI41/XI9/MM4_d
+ N_XI0/XI41/XI9/NET34_XI0/XI41/XI9/MM4_g N_VDD_XI0/XI41/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI9/MM10 N_XI0/XI41/XI9/NET35_XI0/XI41/XI9/MM10_d
+ N_XI0/XI41/XI9/NET36_XI0/XI41/XI9/MM10_g N_VDD_XI0/XI41/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI9/MM11 N_XI0/XI41/XI9/NET36_XI0/XI41/XI9/MM11_d
+ N_XI0/XI41/XI9/NET35_XI0/XI41/XI9/MM11_g N_VDD_XI0/XI41/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI10/MM2 N_XI0/XI41/XI10/NET34_XI0/XI41/XI10/MM2_d
+ N_XI0/XI41/XI10/NET33_XI0/XI41/XI10/MM2_g N_VSS_XI0/XI41/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM3 N_XI0/XI41/XI10/NET33_XI0/XI41/XI10/MM3_d
+ N_WL<78>_XI0/XI41/XI10/MM3_g N_BLN<5>_XI0/XI41/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM0 N_XI0/XI41/XI10/NET34_XI0/XI41/XI10/MM0_d
+ N_WL<78>_XI0/XI41/XI10/MM0_g N_BL<5>_XI0/XI41/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM1 N_XI0/XI41/XI10/NET33_XI0/XI41/XI10/MM1_d
+ N_XI0/XI41/XI10/NET34_XI0/XI41/XI10/MM1_g N_VSS_XI0/XI41/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM9 N_XI0/XI41/XI10/NET36_XI0/XI41/XI10/MM9_d
+ N_WL<79>_XI0/XI41/XI10/MM9_g N_BL<5>_XI0/XI41/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM6 N_XI0/XI41/XI10/NET35_XI0/XI41/XI10/MM6_d
+ N_XI0/XI41/XI10/NET36_XI0/XI41/XI10/MM6_g N_VSS_XI0/XI41/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM7 N_XI0/XI41/XI10/NET36_XI0/XI41/XI10/MM7_d
+ N_XI0/XI41/XI10/NET35_XI0/XI41/XI10/MM7_g N_VSS_XI0/XI41/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM8 N_XI0/XI41/XI10/NET35_XI0/XI41/XI10/MM8_d
+ N_WL<79>_XI0/XI41/XI10/MM8_g N_BLN<5>_XI0/XI41/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI10/MM5 N_XI0/XI41/XI10/NET34_XI0/XI41/XI10/MM5_d
+ N_XI0/XI41/XI10/NET33_XI0/XI41/XI10/MM5_g N_VDD_XI0/XI41/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI10/MM4 N_XI0/XI41/XI10/NET33_XI0/XI41/XI10/MM4_d
+ N_XI0/XI41/XI10/NET34_XI0/XI41/XI10/MM4_g N_VDD_XI0/XI41/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI10/MM10 N_XI0/XI41/XI10/NET35_XI0/XI41/XI10/MM10_d
+ N_XI0/XI41/XI10/NET36_XI0/XI41/XI10/MM10_g N_VDD_XI0/XI41/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI10/MM11 N_XI0/XI41/XI10/NET36_XI0/XI41/XI10/MM11_d
+ N_XI0/XI41/XI10/NET35_XI0/XI41/XI10/MM11_g N_VDD_XI0/XI41/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI11/MM2 N_XI0/XI41/XI11/NET34_XI0/XI41/XI11/MM2_d
+ N_XI0/XI41/XI11/NET33_XI0/XI41/XI11/MM2_g N_VSS_XI0/XI41/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM3 N_XI0/XI41/XI11/NET33_XI0/XI41/XI11/MM3_d
+ N_WL<78>_XI0/XI41/XI11/MM3_g N_BLN<4>_XI0/XI41/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM0 N_XI0/XI41/XI11/NET34_XI0/XI41/XI11/MM0_d
+ N_WL<78>_XI0/XI41/XI11/MM0_g N_BL<4>_XI0/XI41/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM1 N_XI0/XI41/XI11/NET33_XI0/XI41/XI11/MM1_d
+ N_XI0/XI41/XI11/NET34_XI0/XI41/XI11/MM1_g N_VSS_XI0/XI41/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM9 N_XI0/XI41/XI11/NET36_XI0/XI41/XI11/MM9_d
+ N_WL<79>_XI0/XI41/XI11/MM9_g N_BL<4>_XI0/XI41/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM6 N_XI0/XI41/XI11/NET35_XI0/XI41/XI11/MM6_d
+ N_XI0/XI41/XI11/NET36_XI0/XI41/XI11/MM6_g N_VSS_XI0/XI41/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM7 N_XI0/XI41/XI11/NET36_XI0/XI41/XI11/MM7_d
+ N_XI0/XI41/XI11/NET35_XI0/XI41/XI11/MM7_g N_VSS_XI0/XI41/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM8 N_XI0/XI41/XI11/NET35_XI0/XI41/XI11/MM8_d
+ N_WL<79>_XI0/XI41/XI11/MM8_g N_BLN<4>_XI0/XI41/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI11/MM5 N_XI0/XI41/XI11/NET34_XI0/XI41/XI11/MM5_d
+ N_XI0/XI41/XI11/NET33_XI0/XI41/XI11/MM5_g N_VDD_XI0/XI41/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI11/MM4 N_XI0/XI41/XI11/NET33_XI0/XI41/XI11/MM4_d
+ N_XI0/XI41/XI11/NET34_XI0/XI41/XI11/MM4_g N_VDD_XI0/XI41/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI11/MM10 N_XI0/XI41/XI11/NET35_XI0/XI41/XI11/MM10_d
+ N_XI0/XI41/XI11/NET36_XI0/XI41/XI11/MM10_g N_VDD_XI0/XI41/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI11/MM11 N_XI0/XI41/XI11/NET36_XI0/XI41/XI11/MM11_d
+ N_XI0/XI41/XI11/NET35_XI0/XI41/XI11/MM11_g N_VDD_XI0/XI41/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI12/MM2 N_XI0/XI41/XI12/NET34_XI0/XI41/XI12/MM2_d
+ N_XI0/XI41/XI12/NET33_XI0/XI41/XI12/MM2_g N_VSS_XI0/XI41/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM3 N_XI0/XI41/XI12/NET33_XI0/XI41/XI12/MM3_d
+ N_WL<78>_XI0/XI41/XI12/MM3_g N_BLN<3>_XI0/XI41/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM0 N_XI0/XI41/XI12/NET34_XI0/XI41/XI12/MM0_d
+ N_WL<78>_XI0/XI41/XI12/MM0_g N_BL<3>_XI0/XI41/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM1 N_XI0/XI41/XI12/NET33_XI0/XI41/XI12/MM1_d
+ N_XI0/XI41/XI12/NET34_XI0/XI41/XI12/MM1_g N_VSS_XI0/XI41/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM9 N_XI0/XI41/XI12/NET36_XI0/XI41/XI12/MM9_d
+ N_WL<79>_XI0/XI41/XI12/MM9_g N_BL<3>_XI0/XI41/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM6 N_XI0/XI41/XI12/NET35_XI0/XI41/XI12/MM6_d
+ N_XI0/XI41/XI12/NET36_XI0/XI41/XI12/MM6_g N_VSS_XI0/XI41/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM7 N_XI0/XI41/XI12/NET36_XI0/XI41/XI12/MM7_d
+ N_XI0/XI41/XI12/NET35_XI0/XI41/XI12/MM7_g N_VSS_XI0/XI41/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM8 N_XI0/XI41/XI12/NET35_XI0/XI41/XI12/MM8_d
+ N_WL<79>_XI0/XI41/XI12/MM8_g N_BLN<3>_XI0/XI41/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI12/MM5 N_XI0/XI41/XI12/NET34_XI0/XI41/XI12/MM5_d
+ N_XI0/XI41/XI12/NET33_XI0/XI41/XI12/MM5_g N_VDD_XI0/XI41/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI12/MM4 N_XI0/XI41/XI12/NET33_XI0/XI41/XI12/MM4_d
+ N_XI0/XI41/XI12/NET34_XI0/XI41/XI12/MM4_g N_VDD_XI0/XI41/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI12/MM10 N_XI0/XI41/XI12/NET35_XI0/XI41/XI12/MM10_d
+ N_XI0/XI41/XI12/NET36_XI0/XI41/XI12/MM10_g N_VDD_XI0/XI41/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI12/MM11 N_XI0/XI41/XI12/NET36_XI0/XI41/XI12/MM11_d
+ N_XI0/XI41/XI12/NET35_XI0/XI41/XI12/MM11_g N_VDD_XI0/XI41/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI13/MM2 N_XI0/XI41/XI13/NET34_XI0/XI41/XI13/MM2_d
+ N_XI0/XI41/XI13/NET33_XI0/XI41/XI13/MM2_g N_VSS_XI0/XI41/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM3 N_XI0/XI41/XI13/NET33_XI0/XI41/XI13/MM3_d
+ N_WL<78>_XI0/XI41/XI13/MM3_g N_BLN<2>_XI0/XI41/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM0 N_XI0/XI41/XI13/NET34_XI0/XI41/XI13/MM0_d
+ N_WL<78>_XI0/XI41/XI13/MM0_g N_BL<2>_XI0/XI41/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM1 N_XI0/XI41/XI13/NET33_XI0/XI41/XI13/MM1_d
+ N_XI0/XI41/XI13/NET34_XI0/XI41/XI13/MM1_g N_VSS_XI0/XI41/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM9 N_XI0/XI41/XI13/NET36_XI0/XI41/XI13/MM9_d
+ N_WL<79>_XI0/XI41/XI13/MM9_g N_BL<2>_XI0/XI41/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM6 N_XI0/XI41/XI13/NET35_XI0/XI41/XI13/MM6_d
+ N_XI0/XI41/XI13/NET36_XI0/XI41/XI13/MM6_g N_VSS_XI0/XI41/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM7 N_XI0/XI41/XI13/NET36_XI0/XI41/XI13/MM7_d
+ N_XI0/XI41/XI13/NET35_XI0/XI41/XI13/MM7_g N_VSS_XI0/XI41/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM8 N_XI0/XI41/XI13/NET35_XI0/XI41/XI13/MM8_d
+ N_WL<79>_XI0/XI41/XI13/MM8_g N_BLN<2>_XI0/XI41/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI13/MM5 N_XI0/XI41/XI13/NET34_XI0/XI41/XI13/MM5_d
+ N_XI0/XI41/XI13/NET33_XI0/XI41/XI13/MM5_g N_VDD_XI0/XI41/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI13/MM4 N_XI0/XI41/XI13/NET33_XI0/XI41/XI13/MM4_d
+ N_XI0/XI41/XI13/NET34_XI0/XI41/XI13/MM4_g N_VDD_XI0/XI41/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI13/MM10 N_XI0/XI41/XI13/NET35_XI0/XI41/XI13/MM10_d
+ N_XI0/XI41/XI13/NET36_XI0/XI41/XI13/MM10_g N_VDD_XI0/XI41/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI13/MM11 N_XI0/XI41/XI13/NET36_XI0/XI41/XI13/MM11_d
+ N_XI0/XI41/XI13/NET35_XI0/XI41/XI13/MM11_g N_VDD_XI0/XI41/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI14/MM2 N_XI0/XI41/XI14/NET34_XI0/XI41/XI14/MM2_d
+ N_XI0/XI41/XI14/NET33_XI0/XI41/XI14/MM2_g N_VSS_XI0/XI41/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM3 N_XI0/XI41/XI14/NET33_XI0/XI41/XI14/MM3_d
+ N_WL<78>_XI0/XI41/XI14/MM3_g N_BLN<1>_XI0/XI41/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM0 N_XI0/XI41/XI14/NET34_XI0/XI41/XI14/MM0_d
+ N_WL<78>_XI0/XI41/XI14/MM0_g N_BL<1>_XI0/XI41/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM1 N_XI0/XI41/XI14/NET33_XI0/XI41/XI14/MM1_d
+ N_XI0/XI41/XI14/NET34_XI0/XI41/XI14/MM1_g N_VSS_XI0/XI41/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM9 N_XI0/XI41/XI14/NET36_XI0/XI41/XI14/MM9_d
+ N_WL<79>_XI0/XI41/XI14/MM9_g N_BL<1>_XI0/XI41/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM6 N_XI0/XI41/XI14/NET35_XI0/XI41/XI14/MM6_d
+ N_XI0/XI41/XI14/NET36_XI0/XI41/XI14/MM6_g N_VSS_XI0/XI41/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM7 N_XI0/XI41/XI14/NET36_XI0/XI41/XI14/MM7_d
+ N_XI0/XI41/XI14/NET35_XI0/XI41/XI14/MM7_g N_VSS_XI0/XI41/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM8 N_XI0/XI41/XI14/NET35_XI0/XI41/XI14/MM8_d
+ N_WL<79>_XI0/XI41/XI14/MM8_g N_BLN<1>_XI0/XI41/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI14/MM5 N_XI0/XI41/XI14/NET34_XI0/XI41/XI14/MM5_d
+ N_XI0/XI41/XI14/NET33_XI0/XI41/XI14/MM5_g N_VDD_XI0/XI41/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI14/MM4 N_XI0/XI41/XI14/NET33_XI0/XI41/XI14/MM4_d
+ N_XI0/XI41/XI14/NET34_XI0/XI41/XI14/MM4_g N_VDD_XI0/XI41/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI14/MM10 N_XI0/XI41/XI14/NET35_XI0/XI41/XI14/MM10_d
+ N_XI0/XI41/XI14/NET36_XI0/XI41/XI14/MM10_g N_VDD_XI0/XI41/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI14/MM11 N_XI0/XI41/XI14/NET36_XI0/XI41/XI14/MM11_d
+ N_XI0/XI41/XI14/NET35_XI0/XI41/XI14/MM11_g N_VDD_XI0/XI41/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI15/MM2 N_XI0/XI41/XI15/NET34_XI0/XI41/XI15/MM2_d
+ N_XI0/XI41/XI15/NET33_XI0/XI41/XI15/MM2_g N_VSS_XI0/XI41/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM3 N_XI0/XI41/XI15/NET33_XI0/XI41/XI15/MM3_d
+ N_WL<78>_XI0/XI41/XI15/MM3_g N_BLN<0>_XI0/XI41/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM0 N_XI0/XI41/XI15/NET34_XI0/XI41/XI15/MM0_d
+ N_WL<78>_XI0/XI41/XI15/MM0_g N_BL<0>_XI0/XI41/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM1 N_XI0/XI41/XI15/NET33_XI0/XI41/XI15/MM1_d
+ N_XI0/XI41/XI15/NET34_XI0/XI41/XI15/MM1_g N_VSS_XI0/XI41/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM9 N_XI0/XI41/XI15/NET36_XI0/XI41/XI15/MM9_d
+ N_WL<79>_XI0/XI41/XI15/MM9_g N_BL<0>_XI0/XI41/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM6 N_XI0/XI41/XI15/NET35_XI0/XI41/XI15/MM6_d
+ N_XI0/XI41/XI15/NET36_XI0/XI41/XI15/MM6_g N_VSS_XI0/XI41/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM7 N_XI0/XI41/XI15/NET36_XI0/XI41/XI15/MM7_d
+ N_XI0/XI41/XI15/NET35_XI0/XI41/XI15/MM7_g N_VSS_XI0/XI41/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM8 N_XI0/XI41/XI15/NET35_XI0/XI41/XI15/MM8_d
+ N_WL<79>_XI0/XI41/XI15/MM8_g N_BLN<0>_XI0/XI41/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI41/XI15/MM5 N_XI0/XI41/XI15/NET34_XI0/XI41/XI15/MM5_d
+ N_XI0/XI41/XI15/NET33_XI0/XI41/XI15/MM5_g N_VDD_XI0/XI41/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI15/MM4 N_XI0/XI41/XI15/NET33_XI0/XI41/XI15/MM4_d
+ N_XI0/XI41/XI15/NET34_XI0/XI41/XI15/MM4_g N_VDD_XI0/XI41/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI15/MM10 N_XI0/XI41/XI15/NET35_XI0/XI41/XI15/MM10_d
+ N_XI0/XI41/XI15/NET36_XI0/XI41/XI15/MM10_g N_VDD_XI0/XI41/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI41/XI15/MM11 N_XI0/XI41/XI15/NET36_XI0/XI41/XI15/MM11_d
+ N_XI0/XI41/XI15/NET35_XI0/XI41/XI15/MM11_g N_VDD_XI0/XI41/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI0/MM2 N_XI0/XI42/XI0/NET34_XI0/XI42/XI0/MM2_d
+ N_XI0/XI42/XI0/NET33_XI0/XI42/XI0/MM2_g N_VSS_XI0/XI42/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM3 N_XI0/XI42/XI0/NET33_XI0/XI42/XI0/MM3_d
+ N_WL<80>_XI0/XI42/XI0/MM3_g N_BLN<15>_XI0/XI42/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM0 N_XI0/XI42/XI0/NET34_XI0/XI42/XI0/MM0_d
+ N_WL<80>_XI0/XI42/XI0/MM0_g N_BL<15>_XI0/XI42/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM1 N_XI0/XI42/XI0/NET33_XI0/XI42/XI0/MM1_d
+ N_XI0/XI42/XI0/NET34_XI0/XI42/XI0/MM1_g N_VSS_XI0/XI42/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM9 N_XI0/XI42/XI0/NET36_XI0/XI42/XI0/MM9_d
+ N_WL<81>_XI0/XI42/XI0/MM9_g N_BL<15>_XI0/XI42/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM6 N_XI0/XI42/XI0/NET35_XI0/XI42/XI0/MM6_d
+ N_XI0/XI42/XI0/NET36_XI0/XI42/XI0/MM6_g N_VSS_XI0/XI42/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM7 N_XI0/XI42/XI0/NET36_XI0/XI42/XI0/MM7_d
+ N_XI0/XI42/XI0/NET35_XI0/XI42/XI0/MM7_g N_VSS_XI0/XI42/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM8 N_XI0/XI42/XI0/NET35_XI0/XI42/XI0/MM8_d
+ N_WL<81>_XI0/XI42/XI0/MM8_g N_BLN<15>_XI0/XI42/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI0/MM5 N_XI0/XI42/XI0/NET34_XI0/XI42/XI0/MM5_d
+ N_XI0/XI42/XI0/NET33_XI0/XI42/XI0/MM5_g N_VDD_XI0/XI42/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI0/MM4 N_XI0/XI42/XI0/NET33_XI0/XI42/XI0/MM4_d
+ N_XI0/XI42/XI0/NET34_XI0/XI42/XI0/MM4_g N_VDD_XI0/XI42/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI0/MM10 N_XI0/XI42/XI0/NET35_XI0/XI42/XI0/MM10_d
+ N_XI0/XI42/XI0/NET36_XI0/XI42/XI0/MM10_g N_VDD_XI0/XI42/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI0/MM11 N_XI0/XI42/XI0/NET36_XI0/XI42/XI0/MM11_d
+ N_XI0/XI42/XI0/NET35_XI0/XI42/XI0/MM11_g N_VDD_XI0/XI42/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI1/MM2 N_XI0/XI42/XI1/NET34_XI0/XI42/XI1/MM2_d
+ N_XI0/XI42/XI1/NET33_XI0/XI42/XI1/MM2_g N_VSS_XI0/XI42/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM3 N_XI0/XI42/XI1/NET33_XI0/XI42/XI1/MM3_d
+ N_WL<80>_XI0/XI42/XI1/MM3_g N_BLN<14>_XI0/XI42/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM0 N_XI0/XI42/XI1/NET34_XI0/XI42/XI1/MM0_d
+ N_WL<80>_XI0/XI42/XI1/MM0_g N_BL<14>_XI0/XI42/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM1 N_XI0/XI42/XI1/NET33_XI0/XI42/XI1/MM1_d
+ N_XI0/XI42/XI1/NET34_XI0/XI42/XI1/MM1_g N_VSS_XI0/XI42/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM9 N_XI0/XI42/XI1/NET36_XI0/XI42/XI1/MM9_d
+ N_WL<81>_XI0/XI42/XI1/MM9_g N_BL<14>_XI0/XI42/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM6 N_XI0/XI42/XI1/NET35_XI0/XI42/XI1/MM6_d
+ N_XI0/XI42/XI1/NET36_XI0/XI42/XI1/MM6_g N_VSS_XI0/XI42/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM7 N_XI0/XI42/XI1/NET36_XI0/XI42/XI1/MM7_d
+ N_XI0/XI42/XI1/NET35_XI0/XI42/XI1/MM7_g N_VSS_XI0/XI42/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM8 N_XI0/XI42/XI1/NET35_XI0/XI42/XI1/MM8_d
+ N_WL<81>_XI0/XI42/XI1/MM8_g N_BLN<14>_XI0/XI42/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI1/MM5 N_XI0/XI42/XI1/NET34_XI0/XI42/XI1/MM5_d
+ N_XI0/XI42/XI1/NET33_XI0/XI42/XI1/MM5_g N_VDD_XI0/XI42/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI1/MM4 N_XI0/XI42/XI1/NET33_XI0/XI42/XI1/MM4_d
+ N_XI0/XI42/XI1/NET34_XI0/XI42/XI1/MM4_g N_VDD_XI0/XI42/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI1/MM10 N_XI0/XI42/XI1/NET35_XI0/XI42/XI1/MM10_d
+ N_XI0/XI42/XI1/NET36_XI0/XI42/XI1/MM10_g N_VDD_XI0/XI42/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI1/MM11 N_XI0/XI42/XI1/NET36_XI0/XI42/XI1/MM11_d
+ N_XI0/XI42/XI1/NET35_XI0/XI42/XI1/MM11_g N_VDD_XI0/XI42/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI2/MM2 N_XI0/XI42/XI2/NET34_XI0/XI42/XI2/MM2_d
+ N_XI0/XI42/XI2/NET33_XI0/XI42/XI2/MM2_g N_VSS_XI0/XI42/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM3 N_XI0/XI42/XI2/NET33_XI0/XI42/XI2/MM3_d
+ N_WL<80>_XI0/XI42/XI2/MM3_g N_BLN<13>_XI0/XI42/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM0 N_XI0/XI42/XI2/NET34_XI0/XI42/XI2/MM0_d
+ N_WL<80>_XI0/XI42/XI2/MM0_g N_BL<13>_XI0/XI42/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM1 N_XI0/XI42/XI2/NET33_XI0/XI42/XI2/MM1_d
+ N_XI0/XI42/XI2/NET34_XI0/XI42/XI2/MM1_g N_VSS_XI0/XI42/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM9 N_XI0/XI42/XI2/NET36_XI0/XI42/XI2/MM9_d
+ N_WL<81>_XI0/XI42/XI2/MM9_g N_BL<13>_XI0/XI42/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM6 N_XI0/XI42/XI2/NET35_XI0/XI42/XI2/MM6_d
+ N_XI0/XI42/XI2/NET36_XI0/XI42/XI2/MM6_g N_VSS_XI0/XI42/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM7 N_XI0/XI42/XI2/NET36_XI0/XI42/XI2/MM7_d
+ N_XI0/XI42/XI2/NET35_XI0/XI42/XI2/MM7_g N_VSS_XI0/XI42/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM8 N_XI0/XI42/XI2/NET35_XI0/XI42/XI2/MM8_d
+ N_WL<81>_XI0/XI42/XI2/MM8_g N_BLN<13>_XI0/XI42/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI2/MM5 N_XI0/XI42/XI2/NET34_XI0/XI42/XI2/MM5_d
+ N_XI0/XI42/XI2/NET33_XI0/XI42/XI2/MM5_g N_VDD_XI0/XI42/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI2/MM4 N_XI0/XI42/XI2/NET33_XI0/XI42/XI2/MM4_d
+ N_XI0/XI42/XI2/NET34_XI0/XI42/XI2/MM4_g N_VDD_XI0/XI42/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI2/MM10 N_XI0/XI42/XI2/NET35_XI0/XI42/XI2/MM10_d
+ N_XI0/XI42/XI2/NET36_XI0/XI42/XI2/MM10_g N_VDD_XI0/XI42/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI2/MM11 N_XI0/XI42/XI2/NET36_XI0/XI42/XI2/MM11_d
+ N_XI0/XI42/XI2/NET35_XI0/XI42/XI2/MM11_g N_VDD_XI0/XI42/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI3/MM2 N_XI0/XI42/XI3/NET34_XI0/XI42/XI3/MM2_d
+ N_XI0/XI42/XI3/NET33_XI0/XI42/XI3/MM2_g N_VSS_XI0/XI42/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM3 N_XI0/XI42/XI3/NET33_XI0/XI42/XI3/MM3_d
+ N_WL<80>_XI0/XI42/XI3/MM3_g N_BLN<12>_XI0/XI42/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM0 N_XI0/XI42/XI3/NET34_XI0/XI42/XI3/MM0_d
+ N_WL<80>_XI0/XI42/XI3/MM0_g N_BL<12>_XI0/XI42/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM1 N_XI0/XI42/XI3/NET33_XI0/XI42/XI3/MM1_d
+ N_XI0/XI42/XI3/NET34_XI0/XI42/XI3/MM1_g N_VSS_XI0/XI42/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM9 N_XI0/XI42/XI3/NET36_XI0/XI42/XI3/MM9_d
+ N_WL<81>_XI0/XI42/XI3/MM9_g N_BL<12>_XI0/XI42/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM6 N_XI0/XI42/XI3/NET35_XI0/XI42/XI3/MM6_d
+ N_XI0/XI42/XI3/NET36_XI0/XI42/XI3/MM6_g N_VSS_XI0/XI42/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM7 N_XI0/XI42/XI3/NET36_XI0/XI42/XI3/MM7_d
+ N_XI0/XI42/XI3/NET35_XI0/XI42/XI3/MM7_g N_VSS_XI0/XI42/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM8 N_XI0/XI42/XI3/NET35_XI0/XI42/XI3/MM8_d
+ N_WL<81>_XI0/XI42/XI3/MM8_g N_BLN<12>_XI0/XI42/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI3/MM5 N_XI0/XI42/XI3/NET34_XI0/XI42/XI3/MM5_d
+ N_XI0/XI42/XI3/NET33_XI0/XI42/XI3/MM5_g N_VDD_XI0/XI42/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI3/MM4 N_XI0/XI42/XI3/NET33_XI0/XI42/XI3/MM4_d
+ N_XI0/XI42/XI3/NET34_XI0/XI42/XI3/MM4_g N_VDD_XI0/XI42/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI3/MM10 N_XI0/XI42/XI3/NET35_XI0/XI42/XI3/MM10_d
+ N_XI0/XI42/XI3/NET36_XI0/XI42/XI3/MM10_g N_VDD_XI0/XI42/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI3/MM11 N_XI0/XI42/XI3/NET36_XI0/XI42/XI3/MM11_d
+ N_XI0/XI42/XI3/NET35_XI0/XI42/XI3/MM11_g N_VDD_XI0/XI42/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI4/MM2 N_XI0/XI42/XI4/NET34_XI0/XI42/XI4/MM2_d
+ N_XI0/XI42/XI4/NET33_XI0/XI42/XI4/MM2_g N_VSS_XI0/XI42/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM3 N_XI0/XI42/XI4/NET33_XI0/XI42/XI4/MM3_d
+ N_WL<80>_XI0/XI42/XI4/MM3_g N_BLN<11>_XI0/XI42/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM0 N_XI0/XI42/XI4/NET34_XI0/XI42/XI4/MM0_d
+ N_WL<80>_XI0/XI42/XI4/MM0_g N_BL<11>_XI0/XI42/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM1 N_XI0/XI42/XI4/NET33_XI0/XI42/XI4/MM1_d
+ N_XI0/XI42/XI4/NET34_XI0/XI42/XI4/MM1_g N_VSS_XI0/XI42/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM9 N_XI0/XI42/XI4/NET36_XI0/XI42/XI4/MM9_d
+ N_WL<81>_XI0/XI42/XI4/MM9_g N_BL<11>_XI0/XI42/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM6 N_XI0/XI42/XI4/NET35_XI0/XI42/XI4/MM6_d
+ N_XI0/XI42/XI4/NET36_XI0/XI42/XI4/MM6_g N_VSS_XI0/XI42/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM7 N_XI0/XI42/XI4/NET36_XI0/XI42/XI4/MM7_d
+ N_XI0/XI42/XI4/NET35_XI0/XI42/XI4/MM7_g N_VSS_XI0/XI42/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM8 N_XI0/XI42/XI4/NET35_XI0/XI42/XI4/MM8_d
+ N_WL<81>_XI0/XI42/XI4/MM8_g N_BLN<11>_XI0/XI42/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI4/MM5 N_XI0/XI42/XI4/NET34_XI0/XI42/XI4/MM5_d
+ N_XI0/XI42/XI4/NET33_XI0/XI42/XI4/MM5_g N_VDD_XI0/XI42/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI4/MM4 N_XI0/XI42/XI4/NET33_XI0/XI42/XI4/MM4_d
+ N_XI0/XI42/XI4/NET34_XI0/XI42/XI4/MM4_g N_VDD_XI0/XI42/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI4/MM10 N_XI0/XI42/XI4/NET35_XI0/XI42/XI4/MM10_d
+ N_XI0/XI42/XI4/NET36_XI0/XI42/XI4/MM10_g N_VDD_XI0/XI42/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI4/MM11 N_XI0/XI42/XI4/NET36_XI0/XI42/XI4/MM11_d
+ N_XI0/XI42/XI4/NET35_XI0/XI42/XI4/MM11_g N_VDD_XI0/XI42/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI5/MM2 N_XI0/XI42/XI5/NET34_XI0/XI42/XI5/MM2_d
+ N_XI0/XI42/XI5/NET33_XI0/XI42/XI5/MM2_g N_VSS_XI0/XI42/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM3 N_XI0/XI42/XI5/NET33_XI0/XI42/XI5/MM3_d
+ N_WL<80>_XI0/XI42/XI5/MM3_g N_BLN<10>_XI0/XI42/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM0 N_XI0/XI42/XI5/NET34_XI0/XI42/XI5/MM0_d
+ N_WL<80>_XI0/XI42/XI5/MM0_g N_BL<10>_XI0/XI42/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM1 N_XI0/XI42/XI5/NET33_XI0/XI42/XI5/MM1_d
+ N_XI0/XI42/XI5/NET34_XI0/XI42/XI5/MM1_g N_VSS_XI0/XI42/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM9 N_XI0/XI42/XI5/NET36_XI0/XI42/XI5/MM9_d
+ N_WL<81>_XI0/XI42/XI5/MM9_g N_BL<10>_XI0/XI42/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM6 N_XI0/XI42/XI5/NET35_XI0/XI42/XI5/MM6_d
+ N_XI0/XI42/XI5/NET36_XI0/XI42/XI5/MM6_g N_VSS_XI0/XI42/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM7 N_XI0/XI42/XI5/NET36_XI0/XI42/XI5/MM7_d
+ N_XI0/XI42/XI5/NET35_XI0/XI42/XI5/MM7_g N_VSS_XI0/XI42/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM8 N_XI0/XI42/XI5/NET35_XI0/XI42/XI5/MM8_d
+ N_WL<81>_XI0/XI42/XI5/MM8_g N_BLN<10>_XI0/XI42/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI5/MM5 N_XI0/XI42/XI5/NET34_XI0/XI42/XI5/MM5_d
+ N_XI0/XI42/XI5/NET33_XI0/XI42/XI5/MM5_g N_VDD_XI0/XI42/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI5/MM4 N_XI0/XI42/XI5/NET33_XI0/XI42/XI5/MM4_d
+ N_XI0/XI42/XI5/NET34_XI0/XI42/XI5/MM4_g N_VDD_XI0/XI42/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI5/MM10 N_XI0/XI42/XI5/NET35_XI0/XI42/XI5/MM10_d
+ N_XI0/XI42/XI5/NET36_XI0/XI42/XI5/MM10_g N_VDD_XI0/XI42/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI5/MM11 N_XI0/XI42/XI5/NET36_XI0/XI42/XI5/MM11_d
+ N_XI0/XI42/XI5/NET35_XI0/XI42/XI5/MM11_g N_VDD_XI0/XI42/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI6/MM2 N_XI0/XI42/XI6/NET34_XI0/XI42/XI6/MM2_d
+ N_XI0/XI42/XI6/NET33_XI0/XI42/XI6/MM2_g N_VSS_XI0/XI42/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM3 N_XI0/XI42/XI6/NET33_XI0/XI42/XI6/MM3_d
+ N_WL<80>_XI0/XI42/XI6/MM3_g N_BLN<9>_XI0/XI42/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM0 N_XI0/XI42/XI6/NET34_XI0/XI42/XI6/MM0_d
+ N_WL<80>_XI0/XI42/XI6/MM0_g N_BL<9>_XI0/XI42/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM1 N_XI0/XI42/XI6/NET33_XI0/XI42/XI6/MM1_d
+ N_XI0/XI42/XI6/NET34_XI0/XI42/XI6/MM1_g N_VSS_XI0/XI42/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM9 N_XI0/XI42/XI6/NET36_XI0/XI42/XI6/MM9_d
+ N_WL<81>_XI0/XI42/XI6/MM9_g N_BL<9>_XI0/XI42/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM6 N_XI0/XI42/XI6/NET35_XI0/XI42/XI6/MM6_d
+ N_XI0/XI42/XI6/NET36_XI0/XI42/XI6/MM6_g N_VSS_XI0/XI42/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM7 N_XI0/XI42/XI6/NET36_XI0/XI42/XI6/MM7_d
+ N_XI0/XI42/XI6/NET35_XI0/XI42/XI6/MM7_g N_VSS_XI0/XI42/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM8 N_XI0/XI42/XI6/NET35_XI0/XI42/XI6/MM8_d
+ N_WL<81>_XI0/XI42/XI6/MM8_g N_BLN<9>_XI0/XI42/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI6/MM5 N_XI0/XI42/XI6/NET34_XI0/XI42/XI6/MM5_d
+ N_XI0/XI42/XI6/NET33_XI0/XI42/XI6/MM5_g N_VDD_XI0/XI42/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI6/MM4 N_XI0/XI42/XI6/NET33_XI0/XI42/XI6/MM4_d
+ N_XI0/XI42/XI6/NET34_XI0/XI42/XI6/MM4_g N_VDD_XI0/XI42/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI6/MM10 N_XI0/XI42/XI6/NET35_XI0/XI42/XI6/MM10_d
+ N_XI0/XI42/XI6/NET36_XI0/XI42/XI6/MM10_g N_VDD_XI0/XI42/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI6/MM11 N_XI0/XI42/XI6/NET36_XI0/XI42/XI6/MM11_d
+ N_XI0/XI42/XI6/NET35_XI0/XI42/XI6/MM11_g N_VDD_XI0/XI42/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI7/MM2 N_XI0/XI42/XI7/NET34_XI0/XI42/XI7/MM2_d
+ N_XI0/XI42/XI7/NET33_XI0/XI42/XI7/MM2_g N_VSS_XI0/XI42/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM3 N_XI0/XI42/XI7/NET33_XI0/XI42/XI7/MM3_d
+ N_WL<80>_XI0/XI42/XI7/MM3_g N_BLN<8>_XI0/XI42/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM0 N_XI0/XI42/XI7/NET34_XI0/XI42/XI7/MM0_d
+ N_WL<80>_XI0/XI42/XI7/MM0_g N_BL<8>_XI0/XI42/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM1 N_XI0/XI42/XI7/NET33_XI0/XI42/XI7/MM1_d
+ N_XI0/XI42/XI7/NET34_XI0/XI42/XI7/MM1_g N_VSS_XI0/XI42/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM9 N_XI0/XI42/XI7/NET36_XI0/XI42/XI7/MM9_d
+ N_WL<81>_XI0/XI42/XI7/MM9_g N_BL<8>_XI0/XI42/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM6 N_XI0/XI42/XI7/NET35_XI0/XI42/XI7/MM6_d
+ N_XI0/XI42/XI7/NET36_XI0/XI42/XI7/MM6_g N_VSS_XI0/XI42/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM7 N_XI0/XI42/XI7/NET36_XI0/XI42/XI7/MM7_d
+ N_XI0/XI42/XI7/NET35_XI0/XI42/XI7/MM7_g N_VSS_XI0/XI42/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM8 N_XI0/XI42/XI7/NET35_XI0/XI42/XI7/MM8_d
+ N_WL<81>_XI0/XI42/XI7/MM8_g N_BLN<8>_XI0/XI42/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI7/MM5 N_XI0/XI42/XI7/NET34_XI0/XI42/XI7/MM5_d
+ N_XI0/XI42/XI7/NET33_XI0/XI42/XI7/MM5_g N_VDD_XI0/XI42/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI7/MM4 N_XI0/XI42/XI7/NET33_XI0/XI42/XI7/MM4_d
+ N_XI0/XI42/XI7/NET34_XI0/XI42/XI7/MM4_g N_VDD_XI0/XI42/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI7/MM10 N_XI0/XI42/XI7/NET35_XI0/XI42/XI7/MM10_d
+ N_XI0/XI42/XI7/NET36_XI0/XI42/XI7/MM10_g N_VDD_XI0/XI42/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI7/MM11 N_XI0/XI42/XI7/NET36_XI0/XI42/XI7/MM11_d
+ N_XI0/XI42/XI7/NET35_XI0/XI42/XI7/MM11_g N_VDD_XI0/XI42/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI8/MM2 N_XI0/XI42/XI8/NET34_XI0/XI42/XI8/MM2_d
+ N_XI0/XI42/XI8/NET33_XI0/XI42/XI8/MM2_g N_VSS_XI0/XI42/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM3 N_XI0/XI42/XI8/NET33_XI0/XI42/XI8/MM3_d
+ N_WL<80>_XI0/XI42/XI8/MM3_g N_BLN<7>_XI0/XI42/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM0 N_XI0/XI42/XI8/NET34_XI0/XI42/XI8/MM0_d
+ N_WL<80>_XI0/XI42/XI8/MM0_g N_BL<7>_XI0/XI42/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM1 N_XI0/XI42/XI8/NET33_XI0/XI42/XI8/MM1_d
+ N_XI0/XI42/XI8/NET34_XI0/XI42/XI8/MM1_g N_VSS_XI0/XI42/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM9 N_XI0/XI42/XI8/NET36_XI0/XI42/XI8/MM9_d
+ N_WL<81>_XI0/XI42/XI8/MM9_g N_BL<7>_XI0/XI42/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM6 N_XI0/XI42/XI8/NET35_XI0/XI42/XI8/MM6_d
+ N_XI0/XI42/XI8/NET36_XI0/XI42/XI8/MM6_g N_VSS_XI0/XI42/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM7 N_XI0/XI42/XI8/NET36_XI0/XI42/XI8/MM7_d
+ N_XI0/XI42/XI8/NET35_XI0/XI42/XI8/MM7_g N_VSS_XI0/XI42/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM8 N_XI0/XI42/XI8/NET35_XI0/XI42/XI8/MM8_d
+ N_WL<81>_XI0/XI42/XI8/MM8_g N_BLN<7>_XI0/XI42/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI8/MM5 N_XI0/XI42/XI8/NET34_XI0/XI42/XI8/MM5_d
+ N_XI0/XI42/XI8/NET33_XI0/XI42/XI8/MM5_g N_VDD_XI0/XI42/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI8/MM4 N_XI0/XI42/XI8/NET33_XI0/XI42/XI8/MM4_d
+ N_XI0/XI42/XI8/NET34_XI0/XI42/XI8/MM4_g N_VDD_XI0/XI42/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI8/MM10 N_XI0/XI42/XI8/NET35_XI0/XI42/XI8/MM10_d
+ N_XI0/XI42/XI8/NET36_XI0/XI42/XI8/MM10_g N_VDD_XI0/XI42/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI8/MM11 N_XI0/XI42/XI8/NET36_XI0/XI42/XI8/MM11_d
+ N_XI0/XI42/XI8/NET35_XI0/XI42/XI8/MM11_g N_VDD_XI0/XI42/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI9/MM2 N_XI0/XI42/XI9/NET34_XI0/XI42/XI9/MM2_d
+ N_XI0/XI42/XI9/NET33_XI0/XI42/XI9/MM2_g N_VSS_XI0/XI42/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM3 N_XI0/XI42/XI9/NET33_XI0/XI42/XI9/MM3_d
+ N_WL<80>_XI0/XI42/XI9/MM3_g N_BLN<6>_XI0/XI42/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM0 N_XI0/XI42/XI9/NET34_XI0/XI42/XI9/MM0_d
+ N_WL<80>_XI0/XI42/XI9/MM0_g N_BL<6>_XI0/XI42/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM1 N_XI0/XI42/XI9/NET33_XI0/XI42/XI9/MM1_d
+ N_XI0/XI42/XI9/NET34_XI0/XI42/XI9/MM1_g N_VSS_XI0/XI42/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM9 N_XI0/XI42/XI9/NET36_XI0/XI42/XI9/MM9_d
+ N_WL<81>_XI0/XI42/XI9/MM9_g N_BL<6>_XI0/XI42/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM6 N_XI0/XI42/XI9/NET35_XI0/XI42/XI9/MM6_d
+ N_XI0/XI42/XI9/NET36_XI0/XI42/XI9/MM6_g N_VSS_XI0/XI42/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM7 N_XI0/XI42/XI9/NET36_XI0/XI42/XI9/MM7_d
+ N_XI0/XI42/XI9/NET35_XI0/XI42/XI9/MM7_g N_VSS_XI0/XI42/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM8 N_XI0/XI42/XI9/NET35_XI0/XI42/XI9/MM8_d
+ N_WL<81>_XI0/XI42/XI9/MM8_g N_BLN<6>_XI0/XI42/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI9/MM5 N_XI0/XI42/XI9/NET34_XI0/XI42/XI9/MM5_d
+ N_XI0/XI42/XI9/NET33_XI0/XI42/XI9/MM5_g N_VDD_XI0/XI42/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI9/MM4 N_XI0/XI42/XI9/NET33_XI0/XI42/XI9/MM4_d
+ N_XI0/XI42/XI9/NET34_XI0/XI42/XI9/MM4_g N_VDD_XI0/XI42/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI9/MM10 N_XI0/XI42/XI9/NET35_XI0/XI42/XI9/MM10_d
+ N_XI0/XI42/XI9/NET36_XI0/XI42/XI9/MM10_g N_VDD_XI0/XI42/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI9/MM11 N_XI0/XI42/XI9/NET36_XI0/XI42/XI9/MM11_d
+ N_XI0/XI42/XI9/NET35_XI0/XI42/XI9/MM11_g N_VDD_XI0/XI42/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI10/MM2 N_XI0/XI42/XI10/NET34_XI0/XI42/XI10/MM2_d
+ N_XI0/XI42/XI10/NET33_XI0/XI42/XI10/MM2_g N_VSS_XI0/XI42/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM3 N_XI0/XI42/XI10/NET33_XI0/XI42/XI10/MM3_d
+ N_WL<80>_XI0/XI42/XI10/MM3_g N_BLN<5>_XI0/XI42/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM0 N_XI0/XI42/XI10/NET34_XI0/XI42/XI10/MM0_d
+ N_WL<80>_XI0/XI42/XI10/MM0_g N_BL<5>_XI0/XI42/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM1 N_XI0/XI42/XI10/NET33_XI0/XI42/XI10/MM1_d
+ N_XI0/XI42/XI10/NET34_XI0/XI42/XI10/MM1_g N_VSS_XI0/XI42/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM9 N_XI0/XI42/XI10/NET36_XI0/XI42/XI10/MM9_d
+ N_WL<81>_XI0/XI42/XI10/MM9_g N_BL<5>_XI0/XI42/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM6 N_XI0/XI42/XI10/NET35_XI0/XI42/XI10/MM6_d
+ N_XI0/XI42/XI10/NET36_XI0/XI42/XI10/MM6_g N_VSS_XI0/XI42/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM7 N_XI0/XI42/XI10/NET36_XI0/XI42/XI10/MM7_d
+ N_XI0/XI42/XI10/NET35_XI0/XI42/XI10/MM7_g N_VSS_XI0/XI42/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM8 N_XI0/XI42/XI10/NET35_XI0/XI42/XI10/MM8_d
+ N_WL<81>_XI0/XI42/XI10/MM8_g N_BLN<5>_XI0/XI42/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI10/MM5 N_XI0/XI42/XI10/NET34_XI0/XI42/XI10/MM5_d
+ N_XI0/XI42/XI10/NET33_XI0/XI42/XI10/MM5_g N_VDD_XI0/XI42/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI10/MM4 N_XI0/XI42/XI10/NET33_XI0/XI42/XI10/MM4_d
+ N_XI0/XI42/XI10/NET34_XI0/XI42/XI10/MM4_g N_VDD_XI0/XI42/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI10/MM10 N_XI0/XI42/XI10/NET35_XI0/XI42/XI10/MM10_d
+ N_XI0/XI42/XI10/NET36_XI0/XI42/XI10/MM10_g N_VDD_XI0/XI42/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI10/MM11 N_XI0/XI42/XI10/NET36_XI0/XI42/XI10/MM11_d
+ N_XI0/XI42/XI10/NET35_XI0/XI42/XI10/MM11_g N_VDD_XI0/XI42/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI11/MM2 N_XI0/XI42/XI11/NET34_XI0/XI42/XI11/MM2_d
+ N_XI0/XI42/XI11/NET33_XI0/XI42/XI11/MM2_g N_VSS_XI0/XI42/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM3 N_XI0/XI42/XI11/NET33_XI0/XI42/XI11/MM3_d
+ N_WL<80>_XI0/XI42/XI11/MM3_g N_BLN<4>_XI0/XI42/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM0 N_XI0/XI42/XI11/NET34_XI0/XI42/XI11/MM0_d
+ N_WL<80>_XI0/XI42/XI11/MM0_g N_BL<4>_XI0/XI42/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM1 N_XI0/XI42/XI11/NET33_XI0/XI42/XI11/MM1_d
+ N_XI0/XI42/XI11/NET34_XI0/XI42/XI11/MM1_g N_VSS_XI0/XI42/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM9 N_XI0/XI42/XI11/NET36_XI0/XI42/XI11/MM9_d
+ N_WL<81>_XI0/XI42/XI11/MM9_g N_BL<4>_XI0/XI42/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM6 N_XI0/XI42/XI11/NET35_XI0/XI42/XI11/MM6_d
+ N_XI0/XI42/XI11/NET36_XI0/XI42/XI11/MM6_g N_VSS_XI0/XI42/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM7 N_XI0/XI42/XI11/NET36_XI0/XI42/XI11/MM7_d
+ N_XI0/XI42/XI11/NET35_XI0/XI42/XI11/MM7_g N_VSS_XI0/XI42/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM8 N_XI0/XI42/XI11/NET35_XI0/XI42/XI11/MM8_d
+ N_WL<81>_XI0/XI42/XI11/MM8_g N_BLN<4>_XI0/XI42/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI11/MM5 N_XI0/XI42/XI11/NET34_XI0/XI42/XI11/MM5_d
+ N_XI0/XI42/XI11/NET33_XI0/XI42/XI11/MM5_g N_VDD_XI0/XI42/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI11/MM4 N_XI0/XI42/XI11/NET33_XI0/XI42/XI11/MM4_d
+ N_XI0/XI42/XI11/NET34_XI0/XI42/XI11/MM4_g N_VDD_XI0/XI42/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI11/MM10 N_XI0/XI42/XI11/NET35_XI0/XI42/XI11/MM10_d
+ N_XI0/XI42/XI11/NET36_XI0/XI42/XI11/MM10_g N_VDD_XI0/XI42/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI11/MM11 N_XI0/XI42/XI11/NET36_XI0/XI42/XI11/MM11_d
+ N_XI0/XI42/XI11/NET35_XI0/XI42/XI11/MM11_g N_VDD_XI0/XI42/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI12/MM2 N_XI0/XI42/XI12/NET34_XI0/XI42/XI12/MM2_d
+ N_XI0/XI42/XI12/NET33_XI0/XI42/XI12/MM2_g N_VSS_XI0/XI42/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM3 N_XI0/XI42/XI12/NET33_XI0/XI42/XI12/MM3_d
+ N_WL<80>_XI0/XI42/XI12/MM3_g N_BLN<3>_XI0/XI42/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM0 N_XI0/XI42/XI12/NET34_XI0/XI42/XI12/MM0_d
+ N_WL<80>_XI0/XI42/XI12/MM0_g N_BL<3>_XI0/XI42/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM1 N_XI0/XI42/XI12/NET33_XI0/XI42/XI12/MM1_d
+ N_XI0/XI42/XI12/NET34_XI0/XI42/XI12/MM1_g N_VSS_XI0/XI42/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM9 N_XI0/XI42/XI12/NET36_XI0/XI42/XI12/MM9_d
+ N_WL<81>_XI0/XI42/XI12/MM9_g N_BL<3>_XI0/XI42/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM6 N_XI0/XI42/XI12/NET35_XI0/XI42/XI12/MM6_d
+ N_XI0/XI42/XI12/NET36_XI0/XI42/XI12/MM6_g N_VSS_XI0/XI42/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM7 N_XI0/XI42/XI12/NET36_XI0/XI42/XI12/MM7_d
+ N_XI0/XI42/XI12/NET35_XI0/XI42/XI12/MM7_g N_VSS_XI0/XI42/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM8 N_XI0/XI42/XI12/NET35_XI0/XI42/XI12/MM8_d
+ N_WL<81>_XI0/XI42/XI12/MM8_g N_BLN<3>_XI0/XI42/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI12/MM5 N_XI0/XI42/XI12/NET34_XI0/XI42/XI12/MM5_d
+ N_XI0/XI42/XI12/NET33_XI0/XI42/XI12/MM5_g N_VDD_XI0/XI42/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI12/MM4 N_XI0/XI42/XI12/NET33_XI0/XI42/XI12/MM4_d
+ N_XI0/XI42/XI12/NET34_XI0/XI42/XI12/MM4_g N_VDD_XI0/XI42/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI12/MM10 N_XI0/XI42/XI12/NET35_XI0/XI42/XI12/MM10_d
+ N_XI0/XI42/XI12/NET36_XI0/XI42/XI12/MM10_g N_VDD_XI0/XI42/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI12/MM11 N_XI0/XI42/XI12/NET36_XI0/XI42/XI12/MM11_d
+ N_XI0/XI42/XI12/NET35_XI0/XI42/XI12/MM11_g N_VDD_XI0/XI42/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI13/MM2 N_XI0/XI42/XI13/NET34_XI0/XI42/XI13/MM2_d
+ N_XI0/XI42/XI13/NET33_XI0/XI42/XI13/MM2_g N_VSS_XI0/XI42/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM3 N_XI0/XI42/XI13/NET33_XI0/XI42/XI13/MM3_d
+ N_WL<80>_XI0/XI42/XI13/MM3_g N_BLN<2>_XI0/XI42/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM0 N_XI0/XI42/XI13/NET34_XI0/XI42/XI13/MM0_d
+ N_WL<80>_XI0/XI42/XI13/MM0_g N_BL<2>_XI0/XI42/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM1 N_XI0/XI42/XI13/NET33_XI0/XI42/XI13/MM1_d
+ N_XI0/XI42/XI13/NET34_XI0/XI42/XI13/MM1_g N_VSS_XI0/XI42/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM9 N_XI0/XI42/XI13/NET36_XI0/XI42/XI13/MM9_d
+ N_WL<81>_XI0/XI42/XI13/MM9_g N_BL<2>_XI0/XI42/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM6 N_XI0/XI42/XI13/NET35_XI0/XI42/XI13/MM6_d
+ N_XI0/XI42/XI13/NET36_XI0/XI42/XI13/MM6_g N_VSS_XI0/XI42/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM7 N_XI0/XI42/XI13/NET36_XI0/XI42/XI13/MM7_d
+ N_XI0/XI42/XI13/NET35_XI0/XI42/XI13/MM7_g N_VSS_XI0/XI42/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM8 N_XI0/XI42/XI13/NET35_XI0/XI42/XI13/MM8_d
+ N_WL<81>_XI0/XI42/XI13/MM8_g N_BLN<2>_XI0/XI42/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI13/MM5 N_XI0/XI42/XI13/NET34_XI0/XI42/XI13/MM5_d
+ N_XI0/XI42/XI13/NET33_XI0/XI42/XI13/MM5_g N_VDD_XI0/XI42/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI13/MM4 N_XI0/XI42/XI13/NET33_XI0/XI42/XI13/MM4_d
+ N_XI0/XI42/XI13/NET34_XI0/XI42/XI13/MM4_g N_VDD_XI0/XI42/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI13/MM10 N_XI0/XI42/XI13/NET35_XI0/XI42/XI13/MM10_d
+ N_XI0/XI42/XI13/NET36_XI0/XI42/XI13/MM10_g N_VDD_XI0/XI42/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI13/MM11 N_XI0/XI42/XI13/NET36_XI0/XI42/XI13/MM11_d
+ N_XI0/XI42/XI13/NET35_XI0/XI42/XI13/MM11_g N_VDD_XI0/XI42/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI14/MM2 N_XI0/XI42/XI14/NET34_XI0/XI42/XI14/MM2_d
+ N_XI0/XI42/XI14/NET33_XI0/XI42/XI14/MM2_g N_VSS_XI0/XI42/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM3 N_XI0/XI42/XI14/NET33_XI0/XI42/XI14/MM3_d
+ N_WL<80>_XI0/XI42/XI14/MM3_g N_BLN<1>_XI0/XI42/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM0 N_XI0/XI42/XI14/NET34_XI0/XI42/XI14/MM0_d
+ N_WL<80>_XI0/XI42/XI14/MM0_g N_BL<1>_XI0/XI42/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM1 N_XI0/XI42/XI14/NET33_XI0/XI42/XI14/MM1_d
+ N_XI0/XI42/XI14/NET34_XI0/XI42/XI14/MM1_g N_VSS_XI0/XI42/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM9 N_XI0/XI42/XI14/NET36_XI0/XI42/XI14/MM9_d
+ N_WL<81>_XI0/XI42/XI14/MM9_g N_BL<1>_XI0/XI42/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM6 N_XI0/XI42/XI14/NET35_XI0/XI42/XI14/MM6_d
+ N_XI0/XI42/XI14/NET36_XI0/XI42/XI14/MM6_g N_VSS_XI0/XI42/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM7 N_XI0/XI42/XI14/NET36_XI0/XI42/XI14/MM7_d
+ N_XI0/XI42/XI14/NET35_XI0/XI42/XI14/MM7_g N_VSS_XI0/XI42/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM8 N_XI0/XI42/XI14/NET35_XI0/XI42/XI14/MM8_d
+ N_WL<81>_XI0/XI42/XI14/MM8_g N_BLN<1>_XI0/XI42/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI14/MM5 N_XI0/XI42/XI14/NET34_XI0/XI42/XI14/MM5_d
+ N_XI0/XI42/XI14/NET33_XI0/XI42/XI14/MM5_g N_VDD_XI0/XI42/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI14/MM4 N_XI0/XI42/XI14/NET33_XI0/XI42/XI14/MM4_d
+ N_XI0/XI42/XI14/NET34_XI0/XI42/XI14/MM4_g N_VDD_XI0/XI42/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI14/MM10 N_XI0/XI42/XI14/NET35_XI0/XI42/XI14/MM10_d
+ N_XI0/XI42/XI14/NET36_XI0/XI42/XI14/MM10_g N_VDD_XI0/XI42/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI14/MM11 N_XI0/XI42/XI14/NET36_XI0/XI42/XI14/MM11_d
+ N_XI0/XI42/XI14/NET35_XI0/XI42/XI14/MM11_g N_VDD_XI0/XI42/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI15/MM2 N_XI0/XI42/XI15/NET34_XI0/XI42/XI15/MM2_d
+ N_XI0/XI42/XI15/NET33_XI0/XI42/XI15/MM2_g N_VSS_XI0/XI42/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM3 N_XI0/XI42/XI15/NET33_XI0/XI42/XI15/MM3_d
+ N_WL<80>_XI0/XI42/XI15/MM3_g N_BLN<0>_XI0/XI42/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM0 N_XI0/XI42/XI15/NET34_XI0/XI42/XI15/MM0_d
+ N_WL<80>_XI0/XI42/XI15/MM0_g N_BL<0>_XI0/XI42/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM1 N_XI0/XI42/XI15/NET33_XI0/XI42/XI15/MM1_d
+ N_XI0/XI42/XI15/NET34_XI0/XI42/XI15/MM1_g N_VSS_XI0/XI42/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM9 N_XI0/XI42/XI15/NET36_XI0/XI42/XI15/MM9_d
+ N_WL<81>_XI0/XI42/XI15/MM9_g N_BL<0>_XI0/XI42/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM6 N_XI0/XI42/XI15/NET35_XI0/XI42/XI15/MM6_d
+ N_XI0/XI42/XI15/NET36_XI0/XI42/XI15/MM6_g N_VSS_XI0/XI42/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM7 N_XI0/XI42/XI15/NET36_XI0/XI42/XI15/MM7_d
+ N_XI0/XI42/XI15/NET35_XI0/XI42/XI15/MM7_g N_VSS_XI0/XI42/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM8 N_XI0/XI42/XI15/NET35_XI0/XI42/XI15/MM8_d
+ N_WL<81>_XI0/XI42/XI15/MM8_g N_BLN<0>_XI0/XI42/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI42/XI15/MM5 N_XI0/XI42/XI15/NET34_XI0/XI42/XI15/MM5_d
+ N_XI0/XI42/XI15/NET33_XI0/XI42/XI15/MM5_g N_VDD_XI0/XI42/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI15/MM4 N_XI0/XI42/XI15/NET33_XI0/XI42/XI15/MM4_d
+ N_XI0/XI42/XI15/NET34_XI0/XI42/XI15/MM4_g N_VDD_XI0/XI42/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI15/MM10 N_XI0/XI42/XI15/NET35_XI0/XI42/XI15/MM10_d
+ N_XI0/XI42/XI15/NET36_XI0/XI42/XI15/MM10_g N_VDD_XI0/XI42/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI42/XI15/MM11 N_XI0/XI42/XI15/NET36_XI0/XI42/XI15/MM11_d
+ N_XI0/XI42/XI15/NET35_XI0/XI42/XI15/MM11_g N_VDD_XI0/XI42/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI0/MM2 N_XI0/XI43/XI0/NET34_XI0/XI43/XI0/MM2_d
+ N_XI0/XI43/XI0/NET33_XI0/XI43/XI0/MM2_g N_VSS_XI0/XI43/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM3 N_XI0/XI43/XI0/NET33_XI0/XI43/XI0/MM3_d
+ N_WL<82>_XI0/XI43/XI0/MM3_g N_BLN<15>_XI0/XI43/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM0 N_XI0/XI43/XI0/NET34_XI0/XI43/XI0/MM0_d
+ N_WL<82>_XI0/XI43/XI0/MM0_g N_BL<15>_XI0/XI43/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM1 N_XI0/XI43/XI0/NET33_XI0/XI43/XI0/MM1_d
+ N_XI0/XI43/XI0/NET34_XI0/XI43/XI0/MM1_g N_VSS_XI0/XI43/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM9 N_XI0/XI43/XI0/NET36_XI0/XI43/XI0/MM9_d
+ N_WL<83>_XI0/XI43/XI0/MM9_g N_BL<15>_XI0/XI43/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM6 N_XI0/XI43/XI0/NET35_XI0/XI43/XI0/MM6_d
+ N_XI0/XI43/XI0/NET36_XI0/XI43/XI0/MM6_g N_VSS_XI0/XI43/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM7 N_XI0/XI43/XI0/NET36_XI0/XI43/XI0/MM7_d
+ N_XI0/XI43/XI0/NET35_XI0/XI43/XI0/MM7_g N_VSS_XI0/XI43/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM8 N_XI0/XI43/XI0/NET35_XI0/XI43/XI0/MM8_d
+ N_WL<83>_XI0/XI43/XI0/MM8_g N_BLN<15>_XI0/XI43/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI0/MM5 N_XI0/XI43/XI0/NET34_XI0/XI43/XI0/MM5_d
+ N_XI0/XI43/XI0/NET33_XI0/XI43/XI0/MM5_g N_VDD_XI0/XI43/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI0/MM4 N_XI0/XI43/XI0/NET33_XI0/XI43/XI0/MM4_d
+ N_XI0/XI43/XI0/NET34_XI0/XI43/XI0/MM4_g N_VDD_XI0/XI43/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI0/MM10 N_XI0/XI43/XI0/NET35_XI0/XI43/XI0/MM10_d
+ N_XI0/XI43/XI0/NET36_XI0/XI43/XI0/MM10_g N_VDD_XI0/XI43/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI0/MM11 N_XI0/XI43/XI0/NET36_XI0/XI43/XI0/MM11_d
+ N_XI0/XI43/XI0/NET35_XI0/XI43/XI0/MM11_g N_VDD_XI0/XI43/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI1/MM2 N_XI0/XI43/XI1/NET34_XI0/XI43/XI1/MM2_d
+ N_XI0/XI43/XI1/NET33_XI0/XI43/XI1/MM2_g N_VSS_XI0/XI43/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM3 N_XI0/XI43/XI1/NET33_XI0/XI43/XI1/MM3_d
+ N_WL<82>_XI0/XI43/XI1/MM3_g N_BLN<14>_XI0/XI43/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM0 N_XI0/XI43/XI1/NET34_XI0/XI43/XI1/MM0_d
+ N_WL<82>_XI0/XI43/XI1/MM0_g N_BL<14>_XI0/XI43/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM1 N_XI0/XI43/XI1/NET33_XI0/XI43/XI1/MM1_d
+ N_XI0/XI43/XI1/NET34_XI0/XI43/XI1/MM1_g N_VSS_XI0/XI43/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM9 N_XI0/XI43/XI1/NET36_XI0/XI43/XI1/MM9_d
+ N_WL<83>_XI0/XI43/XI1/MM9_g N_BL<14>_XI0/XI43/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM6 N_XI0/XI43/XI1/NET35_XI0/XI43/XI1/MM6_d
+ N_XI0/XI43/XI1/NET36_XI0/XI43/XI1/MM6_g N_VSS_XI0/XI43/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM7 N_XI0/XI43/XI1/NET36_XI0/XI43/XI1/MM7_d
+ N_XI0/XI43/XI1/NET35_XI0/XI43/XI1/MM7_g N_VSS_XI0/XI43/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM8 N_XI0/XI43/XI1/NET35_XI0/XI43/XI1/MM8_d
+ N_WL<83>_XI0/XI43/XI1/MM8_g N_BLN<14>_XI0/XI43/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI1/MM5 N_XI0/XI43/XI1/NET34_XI0/XI43/XI1/MM5_d
+ N_XI0/XI43/XI1/NET33_XI0/XI43/XI1/MM5_g N_VDD_XI0/XI43/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI1/MM4 N_XI0/XI43/XI1/NET33_XI0/XI43/XI1/MM4_d
+ N_XI0/XI43/XI1/NET34_XI0/XI43/XI1/MM4_g N_VDD_XI0/XI43/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI1/MM10 N_XI0/XI43/XI1/NET35_XI0/XI43/XI1/MM10_d
+ N_XI0/XI43/XI1/NET36_XI0/XI43/XI1/MM10_g N_VDD_XI0/XI43/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI1/MM11 N_XI0/XI43/XI1/NET36_XI0/XI43/XI1/MM11_d
+ N_XI0/XI43/XI1/NET35_XI0/XI43/XI1/MM11_g N_VDD_XI0/XI43/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI2/MM2 N_XI0/XI43/XI2/NET34_XI0/XI43/XI2/MM2_d
+ N_XI0/XI43/XI2/NET33_XI0/XI43/XI2/MM2_g N_VSS_XI0/XI43/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM3 N_XI0/XI43/XI2/NET33_XI0/XI43/XI2/MM3_d
+ N_WL<82>_XI0/XI43/XI2/MM3_g N_BLN<13>_XI0/XI43/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM0 N_XI0/XI43/XI2/NET34_XI0/XI43/XI2/MM0_d
+ N_WL<82>_XI0/XI43/XI2/MM0_g N_BL<13>_XI0/XI43/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM1 N_XI0/XI43/XI2/NET33_XI0/XI43/XI2/MM1_d
+ N_XI0/XI43/XI2/NET34_XI0/XI43/XI2/MM1_g N_VSS_XI0/XI43/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM9 N_XI0/XI43/XI2/NET36_XI0/XI43/XI2/MM9_d
+ N_WL<83>_XI0/XI43/XI2/MM9_g N_BL<13>_XI0/XI43/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM6 N_XI0/XI43/XI2/NET35_XI0/XI43/XI2/MM6_d
+ N_XI0/XI43/XI2/NET36_XI0/XI43/XI2/MM6_g N_VSS_XI0/XI43/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM7 N_XI0/XI43/XI2/NET36_XI0/XI43/XI2/MM7_d
+ N_XI0/XI43/XI2/NET35_XI0/XI43/XI2/MM7_g N_VSS_XI0/XI43/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM8 N_XI0/XI43/XI2/NET35_XI0/XI43/XI2/MM8_d
+ N_WL<83>_XI0/XI43/XI2/MM8_g N_BLN<13>_XI0/XI43/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI2/MM5 N_XI0/XI43/XI2/NET34_XI0/XI43/XI2/MM5_d
+ N_XI0/XI43/XI2/NET33_XI0/XI43/XI2/MM5_g N_VDD_XI0/XI43/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI2/MM4 N_XI0/XI43/XI2/NET33_XI0/XI43/XI2/MM4_d
+ N_XI0/XI43/XI2/NET34_XI0/XI43/XI2/MM4_g N_VDD_XI0/XI43/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI2/MM10 N_XI0/XI43/XI2/NET35_XI0/XI43/XI2/MM10_d
+ N_XI0/XI43/XI2/NET36_XI0/XI43/XI2/MM10_g N_VDD_XI0/XI43/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI2/MM11 N_XI0/XI43/XI2/NET36_XI0/XI43/XI2/MM11_d
+ N_XI0/XI43/XI2/NET35_XI0/XI43/XI2/MM11_g N_VDD_XI0/XI43/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI3/MM2 N_XI0/XI43/XI3/NET34_XI0/XI43/XI3/MM2_d
+ N_XI0/XI43/XI3/NET33_XI0/XI43/XI3/MM2_g N_VSS_XI0/XI43/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM3 N_XI0/XI43/XI3/NET33_XI0/XI43/XI3/MM3_d
+ N_WL<82>_XI0/XI43/XI3/MM3_g N_BLN<12>_XI0/XI43/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM0 N_XI0/XI43/XI3/NET34_XI0/XI43/XI3/MM0_d
+ N_WL<82>_XI0/XI43/XI3/MM0_g N_BL<12>_XI0/XI43/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM1 N_XI0/XI43/XI3/NET33_XI0/XI43/XI3/MM1_d
+ N_XI0/XI43/XI3/NET34_XI0/XI43/XI3/MM1_g N_VSS_XI0/XI43/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM9 N_XI0/XI43/XI3/NET36_XI0/XI43/XI3/MM9_d
+ N_WL<83>_XI0/XI43/XI3/MM9_g N_BL<12>_XI0/XI43/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM6 N_XI0/XI43/XI3/NET35_XI0/XI43/XI3/MM6_d
+ N_XI0/XI43/XI3/NET36_XI0/XI43/XI3/MM6_g N_VSS_XI0/XI43/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM7 N_XI0/XI43/XI3/NET36_XI0/XI43/XI3/MM7_d
+ N_XI0/XI43/XI3/NET35_XI0/XI43/XI3/MM7_g N_VSS_XI0/XI43/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM8 N_XI0/XI43/XI3/NET35_XI0/XI43/XI3/MM8_d
+ N_WL<83>_XI0/XI43/XI3/MM8_g N_BLN<12>_XI0/XI43/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI3/MM5 N_XI0/XI43/XI3/NET34_XI0/XI43/XI3/MM5_d
+ N_XI0/XI43/XI3/NET33_XI0/XI43/XI3/MM5_g N_VDD_XI0/XI43/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI3/MM4 N_XI0/XI43/XI3/NET33_XI0/XI43/XI3/MM4_d
+ N_XI0/XI43/XI3/NET34_XI0/XI43/XI3/MM4_g N_VDD_XI0/XI43/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI3/MM10 N_XI0/XI43/XI3/NET35_XI0/XI43/XI3/MM10_d
+ N_XI0/XI43/XI3/NET36_XI0/XI43/XI3/MM10_g N_VDD_XI0/XI43/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI3/MM11 N_XI0/XI43/XI3/NET36_XI0/XI43/XI3/MM11_d
+ N_XI0/XI43/XI3/NET35_XI0/XI43/XI3/MM11_g N_VDD_XI0/XI43/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI4/MM2 N_XI0/XI43/XI4/NET34_XI0/XI43/XI4/MM2_d
+ N_XI0/XI43/XI4/NET33_XI0/XI43/XI4/MM2_g N_VSS_XI0/XI43/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM3 N_XI0/XI43/XI4/NET33_XI0/XI43/XI4/MM3_d
+ N_WL<82>_XI0/XI43/XI4/MM3_g N_BLN<11>_XI0/XI43/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM0 N_XI0/XI43/XI4/NET34_XI0/XI43/XI4/MM0_d
+ N_WL<82>_XI0/XI43/XI4/MM0_g N_BL<11>_XI0/XI43/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM1 N_XI0/XI43/XI4/NET33_XI0/XI43/XI4/MM1_d
+ N_XI0/XI43/XI4/NET34_XI0/XI43/XI4/MM1_g N_VSS_XI0/XI43/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM9 N_XI0/XI43/XI4/NET36_XI0/XI43/XI4/MM9_d
+ N_WL<83>_XI0/XI43/XI4/MM9_g N_BL<11>_XI0/XI43/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM6 N_XI0/XI43/XI4/NET35_XI0/XI43/XI4/MM6_d
+ N_XI0/XI43/XI4/NET36_XI0/XI43/XI4/MM6_g N_VSS_XI0/XI43/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM7 N_XI0/XI43/XI4/NET36_XI0/XI43/XI4/MM7_d
+ N_XI0/XI43/XI4/NET35_XI0/XI43/XI4/MM7_g N_VSS_XI0/XI43/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM8 N_XI0/XI43/XI4/NET35_XI0/XI43/XI4/MM8_d
+ N_WL<83>_XI0/XI43/XI4/MM8_g N_BLN<11>_XI0/XI43/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI4/MM5 N_XI0/XI43/XI4/NET34_XI0/XI43/XI4/MM5_d
+ N_XI0/XI43/XI4/NET33_XI0/XI43/XI4/MM5_g N_VDD_XI0/XI43/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI4/MM4 N_XI0/XI43/XI4/NET33_XI0/XI43/XI4/MM4_d
+ N_XI0/XI43/XI4/NET34_XI0/XI43/XI4/MM4_g N_VDD_XI0/XI43/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI4/MM10 N_XI0/XI43/XI4/NET35_XI0/XI43/XI4/MM10_d
+ N_XI0/XI43/XI4/NET36_XI0/XI43/XI4/MM10_g N_VDD_XI0/XI43/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI4/MM11 N_XI0/XI43/XI4/NET36_XI0/XI43/XI4/MM11_d
+ N_XI0/XI43/XI4/NET35_XI0/XI43/XI4/MM11_g N_VDD_XI0/XI43/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI5/MM2 N_XI0/XI43/XI5/NET34_XI0/XI43/XI5/MM2_d
+ N_XI0/XI43/XI5/NET33_XI0/XI43/XI5/MM2_g N_VSS_XI0/XI43/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM3 N_XI0/XI43/XI5/NET33_XI0/XI43/XI5/MM3_d
+ N_WL<82>_XI0/XI43/XI5/MM3_g N_BLN<10>_XI0/XI43/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM0 N_XI0/XI43/XI5/NET34_XI0/XI43/XI5/MM0_d
+ N_WL<82>_XI0/XI43/XI5/MM0_g N_BL<10>_XI0/XI43/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM1 N_XI0/XI43/XI5/NET33_XI0/XI43/XI5/MM1_d
+ N_XI0/XI43/XI5/NET34_XI0/XI43/XI5/MM1_g N_VSS_XI0/XI43/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM9 N_XI0/XI43/XI5/NET36_XI0/XI43/XI5/MM9_d
+ N_WL<83>_XI0/XI43/XI5/MM9_g N_BL<10>_XI0/XI43/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM6 N_XI0/XI43/XI5/NET35_XI0/XI43/XI5/MM6_d
+ N_XI0/XI43/XI5/NET36_XI0/XI43/XI5/MM6_g N_VSS_XI0/XI43/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM7 N_XI0/XI43/XI5/NET36_XI0/XI43/XI5/MM7_d
+ N_XI0/XI43/XI5/NET35_XI0/XI43/XI5/MM7_g N_VSS_XI0/XI43/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM8 N_XI0/XI43/XI5/NET35_XI0/XI43/XI5/MM8_d
+ N_WL<83>_XI0/XI43/XI5/MM8_g N_BLN<10>_XI0/XI43/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI5/MM5 N_XI0/XI43/XI5/NET34_XI0/XI43/XI5/MM5_d
+ N_XI0/XI43/XI5/NET33_XI0/XI43/XI5/MM5_g N_VDD_XI0/XI43/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI5/MM4 N_XI0/XI43/XI5/NET33_XI0/XI43/XI5/MM4_d
+ N_XI0/XI43/XI5/NET34_XI0/XI43/XI5/MM4_g N_VDD_XI0/XI43/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI5/MM10 N_XI0/XI43/XI5/NET35_XI0/XI43/XI5/MM10_d
+ N_XI0/XI43/XI5/NET36_XI0/XI43/XI5/MM10_g N_VDD_XI0/XI43/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI5/MM11 N_XI0/XI43/XI5/NET36_XI0/XI43/XI5/MM11_d
+ N_XI0/XI43/XI5/NET35_XI0/XI43/XI5/MM11_g N_VDD_XI0/XI43/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI6/MM2 N_XI0/XI43/XI6/NET34_XI0/XI43/XI6/MM2_d
+ N_XI0/XI43/XI6/NET33_XI0/XI43/XI6/MM2_g N_VSS_XI0/XI43/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM3 N_XI0/XI43/XI6/NET33_XI0/XI43/XI6/MM3_d
+ N_WL<82>_XI0/XI43/XI6/MM3_g N_BLN<9>_XI0/XI43/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM0 N_XI0/XI43/XI6/NET34_XI0/XI43/XI6/MM0_d
+ N_WL<82>_XI0/XI43/XI6/MM0_g N_BL<9>_XI0/XI43/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM1 N_XI0/XI43/XI6/NET33_XI0/XI43/XI6/MM1_d
+ N_XI0/XI43/XI6/NET34_XI0/XI43/XI6/MM1_g N_VSS_XI0/XI43/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM9 N_XI0/XI43/XI6/NET36_XI0/XI43/XI6/MM9_d
+ N_WL<83>_XI0/XI43/XI6/MM9_g N_BL<9>_XI0/XI43/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM6 N_XI0/XI43/XI6/NET35_XI0/XI43/XI6/MM6_d
+ N_XI0/XI43/XI6/NET36_XI0/XI43/XI6/MM6_g N_VSS_XI0/XI43/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM7 N_XI0/XI43/XI6/NET36_XI0/XI43/XI6/MM7_d
+ N_XI0/XI43/XI6/NET35_XI0/XI43/XI6/MM7_g N_VSS_XI0/XI43/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM8 N_XI0/XI43/XI6/NET35_XI0/XI43/XI6/MM8_d
+ N_WL<83>_XI0/XI43/XI6/MM8_g N_BLN<9>_XI0/XI43/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI6/MM5 N_XI0/XI43/XI6/NET34_XI0/XI43/XI6/MM5_d
+ N_XI0/XI43/XI6/NET33_XI0/XI43/XI6/MM5_g N_VDD_XI0/XI43/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI6/MM4 N_XI0/XI43/XI6/NET33_XI0/XI43/XI6/MM4_d
+ N_XI0/XI43/XI6/NET34_XI0/XI43/XI6/MM4_g N_VDD_XI0/XI43/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI6/MM10 N_XI0/XI43/XI6/NET35_XI0/XI43/XI6/MM10_d
+ N_XI0/XI43/XI6/NET36_XI0/XI43/XI6/MM10_g N_VDD_XI0/XI43/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI6/MM11 N_XI0/XI43/XI6/NET36_XI0/XI43/XI6/MM11_d
+ N_XI0/XI43/XI6/NET35_XI0/XI43/XI6/MM11_g N_VDD_XI0/XI43/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI7/MM2 N_XI0/XI43/XI7/NET34_XI0/XI43/XI7/MM2_d
+ N_XI0/XI43/XI7/NET33_XI0/XI43/XI7/MM2_g N_VSS_XI0/XI43/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM3 N_XI0/XI43/XI7/NET33_XI0/XI43/XI7/MM3_d
+ N_WL<82>_XI0/XI43/XI7/MM3_g N_BLN<8>_XI0/XI43/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM0 N_XI0/XI43/XI7/NET34_XI0/XI43/XI7/MM0_d
+ N_WL<82>_XI0/XI43/XI7/MM0_g N_BL<8>_XI0/XI43/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM1 N_XI0/XI43/XI7/NET33_XI0/XI43/XI7/MM1_d
+ N_XI0/XI43/XI7/NET34_XI0/XI43/XI7/MM1_g N_VSS_XI0/XI43/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM9 N_XI0/XI43/XI7/NET36_XI0/XI43/XI7/MM9_d
+ N_WL<83>_XI0/XI43/XI7/MM9_g N_BL<8>_XI0/XI43/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM6 N_XI0/XI43/XI7/NET35_XI0/XI43/XI7/MM6_d
+ N_XI0/XI43/XI7/NET36_XI0/XI43/XI7/MM6_g N_VSS_XI0/XI43/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM7 N_XI0/XI43/XI7/NET36_XI0/XI43/XI7/MM7_d
+ N_XI0/XI43/XI7/NET35_XI0/XI43/XI7/MM7_g N_VSS_XI0/XI43/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM8 N_XI0/XI43/XI7/NET35_XI0/XI43/XI7/MM8_d
+ N_WL<83>_XI0/XI43/XI7/MM8_g N_BLN<8>_XI0/XI43/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI7/MM5 N_XI0/XI43/XI7/NET34_XI0/XI43/XI7/MM5_d
+ N_XI0/XI43/XI7/NET33_XI0/XI43/XI7/MM5_g N_VDD_XI0/XI43/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI7/MM4 N_XI0/XI43/XI7/NET33_XI0/XI43/XI7/MM4_d
+ N_XI0/XI43/XI7/NET34_XI0/XI43/XI7/MM4_g N_VDD_XI0/XI43/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI7/MM10 N_XI0/XI43/XI7/NET35_XI0/XI43/XI7/MM10_d
+ N_XI0/XI43/XI7/NET36_XI0/XI43/XI7/MM10_g N_VDD_XI0/XI43/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI7/MM11 N_XI0/XI43/XI7/NET36_XI0/XI43/XI7/MM11_d
+ N_XI0/XI43/XI7/NET35_XI0/XI43/XI7/MM11_g N_VDD_XI0/XI43/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI8/MM2 N_XI0/XI43/XI8/NET34_XI0/XI43/XI8/MM2_d
+ N_XI0/XI43/XI8/NET33_XI0/XI43/XI8/MM2_g N_VSS_XI0/XI43/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM3 N_XI0/XI43/XI8/NET33_XI0/XI43/XI8/MM3_d
+ N_WL<82>_XI0/XI43/XI8/MM3_g N_BLN<7>_XI0/XI43/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM0 N_XI0/XI43/XI8/NET34_XI0/XI43/XI8/MM0_d
+ N_WL<82>_XI0/XI43/XI8/MM0_g N_BL<7>_XI0/XI43/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM1 N_XI0/XI43/XI8/NET33_XI0/XI43/XI8/MM1_d
+ N_XI0/XI43/XI8/NET34_XI0/XI43/XI8/MM1_g N_VSS_XI0/XI43/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM9 N_XI0/XI43/XI8/NET36_XI0/XI43/XI8/MM9_d
+ N_WL<83>_XI0/XI43/XI8/MM9_g N_BL<7>_XI0/XI43/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM6 N_XI0/XI43/XI8/NET35_XI0/XI43/XI8/MM6_d
+ N_XI0/XI43/XI8/NET36_XI0/XI43/XI8/MM6_g N_VSS_XI0/XI43/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM7 N_XI0/XI43/XI8/NET36_XI0/XI43/XI8/MM7_d
+ N_XI0/XI43/XI8/NET35_XI0/XI43/XI8/MM7_g N_VSS_XI0/XI43/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM8 N_XI0/XI43/XI8/NET35_XI0/XI43/XI8/MM8_d
+ N_WL<83>_XI0/XI43/XI8/MM8_g N_BLN<7>_XI0/XI43/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI8/MM5 N_XI0/XI43/XI8/NET34_XI0/XI43/XI8/MM5_d
+ N_XI0/XI43/XI8/NET33_XI0/XI43/XI8/MM5_g N_VDD_XI0/XI43/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI8/MM4 N_XI0/XI43/XI8/NET33_XI0/XI43/XI8/MM4_d
+ N_XI0/XI43/XI8/NET34_XI0/XI43/XI8/MM4_g N_VDD_XI0/XI43/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI8/MM10 N_XI0/XI43/XI8/NET35_XI0/XI43/XI8/MM10_d
+ N_XI0/XI43/XI8/NET36_XI0/XI43/XI8/MM10_g N_VDD_XI0/XI43/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI8/MM11 N_XI0/XI43/XI8/NET36_XI0/XI43/XI8/MM11_d
+ N_XI0/XI43/XI8/NET35_XI0/XI43/XI8/MM11_g N_VDD_XI0/XI43/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI9/MM2 N_XI0/XI43/XI9/NET34_XI0/XI43/XI9/MM2_d
+ N_XI0/XI43/XI9/NET33_XI0/XI43/XI9/MM2_g N_VSS_XI0/XI43/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM3 N_XI0/XI43/XI9/NET33_XI0/XI43/XI9/MM3_d
+ N_WL<82>_XI0/XI43/XI9/MM3_g N_BLN<6>_XI0/XI43/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM0 N_XI0/XI43/XI9/NET34_XI0/XI43/XI9/MM0_d
+ N_WL<82>_XI0/XI43/XI9/MM0_g N_BL<6>_XI0/XI43/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM1 N_XI0/XI43/XI9/NET33_XI0/XI43/XI9/MM1_d
+ N_XI0/XI43/XI9/NET34_XI0/XI43/XI9/MM1_g N_VSS_XI0/XI43/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM9 N_XI0/XI43/XI9/NET36_XI0/XI43/XI9/MM9_d
+ N_WL<83>_XI0/XI43/XI9/MM9_g N_BL<6>_XI0/XI43/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM6 N_XI0/XI43/XI9/NET35_XI0/XI43/XI9/MM6_d
+ N_XI0/XI43/XI9/NET36_XI0/XI43/XI9/MM6_g N_VSS_XI0/XI43/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM7 N_XI0/XI43/XI9/NET36_XI0/XI43/XI9/MM7_d
+ N_XI0/XI43/XI9/NET35_XI0/XI43/XI9/MM7_g N_VSS_XI0/XI43/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM8 N_XI0/XI43/XI9/NET35_XI0/XI43/XI9/MM8_d
+ N_WL<83>_XI0/XI43/XI9/MM8_g N_BLN<6>_XI0/XI43/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI9/MM5 N_XI0/XI43/XI9/NET34_XI0/XI43/XI9/MM5_d
+ N_XI0/XI43/XI9/NET33_XI0/XI43/XI9/MM5_g N_VDD_XI0/XI43/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI9/MM4 N_XI0/XI43/XI9/NET33_XI0/XI43/XI9/MM4_d
+ N_XI0/XI43/XI9/NET34_XI0/XI43/XI9/MM4_g N_VDD_XI0/XI43/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI9/MM10 N_XI0/XI43/XI9/NET35_XI0/XI43/XI9/MM10_d
+ N_XI0/XI43/XI9/NET36_XI0/XI43/XI9/MM10_g N_VDD_XI0/XI43/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI9/MM11 N_XI0/XI43/XI9/NET36_XI0/XI43/XI9/MM11_d
+ N_XI0/XI43/XI9/NET35_XI0/XI43/XI9/MM11_g N_VDD_XI0/XI43/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI10/MM2 N_XI0/XI43/XI10/NET34_XI0/XI43/XI10/MM2_d
+ N_XI0/XI43/XI10/NET33_XI0/XI43/XI10/MM2_g N_VSS_XI0/XI43/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM3 N_XI0/XI43/XI10/NET33_XI0/XI43/XI10/MM3_d
+ N_WL<82>_XI0/XI43/XI10/MM3_g N_BLN<5>_XI0/XI43/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM0 N_XI0/XI43/XI10/NET34_XI0/XI43/XI10/MM0_d
+ N_WL<82>_XI0/XI43/XI10/MM0_g N_BL<5>_XI0/XI43/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM1 N_XI0/XI43/XI10/NET33_XI0/XI43/XI10/MM1_d
+ N_XI0/XI43/XI10/NET34_XI0/XI43/XI10/MM1_g N_VSS_XI0/XI43/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM9 N_XI0/XI43/XI10/NET36_XI0/XI43/XI10/MM9_d
+ N_WL<83>_XI0/XI43/XI10/MM9_g N_BL<5>_XI0/XI43/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM6 N_XI0/XI43/XI10/NET35_XI0/XI43/XI10/MM6_d
+ N_XI0/XI43/XI10/NET36_XI0/XI43/XI10/MM6_g N_VSS_XI0/XI43/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM7 N_XI0/XI43/XI10/NET36_XI0/XI43/XI10/MM7_d
+ N_XI0/XI43/XI10/NET35_XI0/XI43/XI10/MM7_g N_VSS_XI0/XI43/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM8 N_XI0/XI43/XI10/NET35_XI0/XI43/XI10/MM8_d
+ N_WL<83>_XI0/XI43/XI10/MM8_g N_BLN<5>_XI0/XI43/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI10/MM5 N_XI0/XI43/XI10/NET34_XI0/XI43/XI10/MM5_d
+ N_XI0/XI43/XI10/NET33_XI0/XI43/XI10/MM5_g N_VDD_XI0/XI43/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI10/MM4 N_XI0/XI43/XI10/NET33_XI0/XI43/XI10/MM4_d
+ N_XI0/XI43/XI10/NET34_XI0/XI43/XI10/MM4_g N_VDD_XI0/XI43/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI10/MM10 N_XI0/XI43/XI10/NET35_XI0/XI43/XI10/MM10_d
+ N_XI0/XI43/XI10/NET36_XI0/XI43/XI10/MM10_g N_VDD_XI0/XI43/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI10/MM11 N_XI0/XI43/XI10/NET36_XI0/XI43/XI10/MM11_d
+ N_XI0/XI43/XI10/NET35_XI0/XI43/XI10/MM11_g N_VDD_XI0/XI43/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI11/MM2 N_XI0/XI43/XI11/NET34_XI0/XI43/XI11/MM2_d
+ N_XI0/XI43/XI11/NET33_XI0/XI43/XI11/MM2_g N_VSS_XI0/XI43/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM3 N_XI0/XI43/XI11/NET33_XI0/XI43/XI11/MM3_d
+ N_WL<82>_XI0/XI43/XI11/MM3_g N_BLN<4>_XI0/XI43/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM0 N_XI0/XI43/XI11/NET34_XI0/XI43/XI11/MM0_d
+ N_WL<82>_XI0/XI43/XI11/MM0_g N_BL<4>_XI0/XI43/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM1 N_XI0/XI43/XI11/NET33_XI0/XI43/XI11/MM1_d
+ N_XI0/XI43/XI11/NET34_XI0/XI43/XI11/MM1_g N_VSS_XI0/XI43/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM9 N_XI0/XI43/XI11/NET36_XI0/XI43/XI11/MM9_d
+ N_WL<83>_XI0/XI43/XI11/MM9_g N_BL<4>_XI0/XI43/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM6 N_XI0/XI43/XI11/NET35_XI0/XI43/XI11/MM6_d
+ N_XI0/XI43/XI11/NET36_XI0/XI43/XI11/MM6_g N_VSS_XI0/XI43/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM7 N_XI0/XI43/XI11/NET36_XI0/XI43/XI11/MM7_d
+ N_XI0/XI43/XI11/NET35_XI0/XI43/XI11/MM7_g N_VSS_XI0/XI43/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM8 N_XI0/XI43/XI11/NET35_XI0/XI43/XI11/MM8_d
+ N_WL<83>_XI0/XI43/XI11/MM8_g N_BLN<4>_XI0/XI43/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI11/MM5 N_XI0/XI43/XI11/NET34_XI0/XI43/XI11/MM5_d
+ N_XI0/XI43/XI11/NET33_XI0/XI43/XI11/MM5_g N_VDD_XI0/XI43/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI11/MM4 N_XI0/XI43/XI11/NET33_XI0/XI43/XI11/MM4_d
+ N_XI0/XI43/XI11/NET34_XI0/XI43/XI11/MM4_g N_VDD_XI0/XI43/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI11/MM10 N_XI0/XI43/XI11/NET35_XI0/XI43/XI11/MM10_d
+ N_XI0/XI43/XI11/NET36_XI0/XI43/XI11/MM10_g N_VDD_XI0/XI43/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI11/MM11 N_XI0/XI43/XI11/NET36_XI0/XI43/XI11/MM11_d
+ N_XI0/XI43/XI11/NET35_XI0/XI43/XI11/MM11_g N_VDD_XI0/XI43/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI12/MM2 N_XI0/XI43/XI12/NET34_XI0/XI43/XI12/MM2_d
+ N_XI0/XI43/XI12/NET33_XI0/XI43/XI12/MM2_g N_VSS_XI0/XI43/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM3 N_XI0/XI43/XI12/NET33_XI0/XI43/XI12/MM3_d
+ N_WL<82>_XI0/XI43/XI12/MM3_g N_BLN<3>_XI0/XI43/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM0 N_XI0/XI43/XI12/NET34_XI0/XI43/XI12/MM0_d
+ N_WL<82>_XI0/XI43/XI12/MM0_g N_BL<3>_XI0/XI43/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM1 N_XI0/XI43/XI12/NET33_XI0/XI43/XI12/MM1_d
+ N_XI0/XI43/XI12/NET34_XI0/XI43/XI12/MM1_g N_VSS_XI0/XI43/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM9 N_XI0/XI43/XI12/NET36_XI0/XI43/XI12/MM9_d
+ N_WL<83>_XI0/XI43/XI12/MM9_g N_BL<3>_XI0/XI43/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM6 N_XI0/XI43/XI12/NET35_XI0/XI43/XI12/MM6_d
+ N_XI0/XI43/XI12/NET36_XI0/XI43/XI12/MM6_g N_VSS_XI0/XI43/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM7 N_XI0/XI43/XI12/NET36_XI0/XI43/XI12/MM7_d
+ N_XI0/XI43/XI12/NET35_XI0/XI43/XI12/MM7_g N_VSS_XI0/XI43/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM8 N_XI0/XI43/XI12/NET35_XI0/XI43/XI12/MM8_d
+ N_WL<83>_XI0/XI43/XI12/MM8_g N_BLN<3>_XI0/XI43/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI12/MM5 N_XI0/XI43/XI12/NET34_XI0/XI43/XI12/MM5_d
+ N_XI0/XI43/XI12/NET33_XI0/XI43/XI12/MM5_g N_VDD_XI0/XI43/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI12/MM4 N_XI0/XI43/XI12/NET33_XI0/XI43/XI12/MM4_d
+ N_XI0/XI43/XI12/NET34_XI0/XI43/XI12/MM4_g N_VDD_XI0/XI43/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI12/MM10 N_XI0/XI43/XI12/NET35_XI0/XI43/XI12/MM10_d
+ N_XI0/XI43/XI12/NET36_XI0/XI43/XI12/MM10_g N_VDD_XI0/XI43/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI12/MM11 N_XI0/XI43/XI12/NET36_XI0/XI43/XI12/MM11_d
+ N_XI0/XI43/XI12/NET35_XI0/XI43/XI12/MM11_g N_VDD_XI0/XI43/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI13/MM2 N_XI0/XI43/XI13/NET34_XI0/XI43/XI13/MM2_d
+ N_XI0/XI43/XI13/NET33_XI0/XI43/XI13/MM2_g N_VSS_XI0/XI43/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM3 N_XI0/XI43/XI13/NET33_XI0/XI43/XI13/MM3_d
+ N_WL<82>_XI0/XI43/XI13/MM3_g N_BLN<2>_XI0/XI43/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM0 N_XI0/XI43/XI13/NET34_XI0/XI43/XI13/MM0_d
+ N_WL<82>_XI0/XI43/XI13/MM0_g N_BL<2>_XI0/XI43/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM1 N_XI0/XI43/XI13/NET33_XI0/XI43/XI13/MM1_d
+ N_XI0/XI43/XI13/NET34_XI0/XI43/XI13/MM1_g N_VSS_XI0/XI43/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM9 N_XI0/XI43/XI13/NET36_XI0/XI43/XI13/MM9_d
+ N_WL<83>_XI0/XI43/XI13/MM9_g N_BL<2>_XI0/XI43/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM6 N_XI0/XI43/XI13/NET35_XI0/XI43/XI13/MM6_d
+ N_XI0/XI43/XI13/NET36_XI0/XI43/XI13/MM6_g N_VSS_XI0/XI43/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM7 N_XI0/XI43/XI13/NET36_XI0/XI43/XI13/MM7_d
+ N_XI0/XI43/XI13/NET35_XI0/XI43/XI13/MM7_g N_VSS_XI0/XI43/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM8 N_XI0/XI43/XI13/NET35_XI0/XI43/XI13/MM8_d
+ N_WL<83>_XI0/XI43/XI13/MM8_g N_BLN<2>_XI0/XI43/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI13/MM5 N_XI0/XI43/XI13/NET34_XI0/XI43/XI13/MM5_d
+ N_XI0/XI43/XI13/NET33_XI0/XI43/XI13/MM5_g N_VDD_XI0/XI43/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI13/MM4 N_XI0/XI43/XI13/NET33_XI0/XI43/XI13/MM4_d
+ N_XI0/XI43/XI13/NET34_XI0/XI43/XI13/MM4_g N_VDD_XI0/XI43/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI13/MM10 N_XI0/XI43/XI13/NET35_XI0/XI43/XI13/MM10_d
+ N_XI0/XI43/XI13/NET36_XI0/XI43/XI13/MM10_g N_VDD_XI0/XI43/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI13/MM11 N_XI0/XI43/XI13/NET36_XI0/XI43/XI13/MM11_d
+ N_XI0/XI43/XI13/NET35_XI0/XI43/XI13/MM11_g N_VDD_XI0/XI43/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI14/MM2 N_XI0/XI43/XI14/NET34_XI0/XI43/XI14/MM2_d
+ N_XI0/XI43/XI14/NET33_XI0/XI43/XI14/MM2_g N_VSS_XI0/XI43/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM3 N_XI0/XI43/XI14/NET33_XI0/XI43/XI14/MM3_d
+ N_WL<82>_XI0/XI43/XI14/MM3_g N_BLN<1>_XI0/XI43/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM0 N_XI0/XI43/XI14/NET34_XI0/XI43/XI14/MM0_d
+ N_WL<82>_XI0/XI43/XI14/MM0_g N_BL<1>_XI0/XI43/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM1 N_XI0/XI43/XI14/NET33_XI0/XI43/XI14/MM1_d
+ N_XI0/XI43/XI14/NET34_XI0/XI43/XI14/MM1_g N_VSS_XI0/XI43/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM9 N_XI0/XI43/XI14/NET36_XI0/XI43/XI14/MM9_d
+ N_WL<83>_XI0/XI43/XI14/MM9_g N_BL<1>_XI0/XI43/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM6 N_XI0/XI43/XI14/NET35_XI0/XI43/XI14/MM6_d
+ N_XI0/XI43/XI14/NET36_XI0/XI43/XI14/MM6_g N_VSS_XI0/XI43/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM7 N_XI0/XI43/XI14/NET36_XI0/XI43/XI14/MM7_d
+ N_XI0/XI43/XI14/NET35_XI0/XI43/XI14/MM7_g N_VSS_XI0/XI43/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM8 N_XI0/XI43/XI14/NET35_XI0/XI43/XI14/MM8_d
+ N_WL<83>_XI0/XI43/XI14/MM8_g N_BLN<1>_XI0/XI43/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI14/MM5 N_XI0/XI43/XI14/NET34_XI0/XI43/XI14/MM5_d
+ N_XI0/XI43/XI14/NET33_XI0/XI43/XI14/MM5_g N_VDD_XI0/XI43/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI14/MM4 N_XI0/XI43/XI14/NET33_XI0/XI43/XI14/MM4_d
+ N_XI0/XI43/XI14/NET34_XI0/XI43/XI14/MM4_g N_VDD_XI0/XI43/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI14/MM10 N_XI0/XI43/XI14/NET35_XI0/XI43/XI14/MM10_d
+ N_XI0/XI43/XI14/NET36_XI0/XI43/XI14/MM10_g N_VDD_XI0/XI43/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI14/MM11 N_XI0/XI43/XI14/NET36_XI0/XI43/XI14/MM11_d
+ N_XI0/XI43/XI14/NET35_XI0/XI43/XI14/MM11_g N_VDD_XI0/XI43/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI15/MM2 N_XI0/XI43/XI15/NET34_XI0/XI43/XI15/MM2_d
+ N_XI0/XI43/XI15/NET33_XI0/XI43/XI15/MM2_g N_VSS_XI0/XI43/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM3 N_XI0/XI43/XI15/NET33_XI0/XI43/XI15/MM3_d
+ N_WL<82>_XI0/XI43/XI15/MM3_g N_BLN<0>_XI0/XI43/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM0 N_XI0/XI43/XI15/NET34_XI0/XI43/XI15/MM0_d
+ N_WL<82>_XI0/XI43/XI15/MM0_g N_BL<0>_XI0/XI43/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM1 N_XI0/XI43/XI15/NET33_XI0/XI43/XI15/MM1_d
+ N_XI0/XI43/XI15/NET34_XI0/XI43/XI15/MM1_g N_VSS_XI0/XI43/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM9 N_XI0/XI43/XI15/NET36_XI0/XI43/XI15/MM9_d
+ N_WL<83>_XI0/XI43/XI15/MM9_g N_BL<0>_XI0/XI43/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM6 N_XI0/XI43/XI15/NET35_XI0/XI43/XI15/MM6_d
+ N_XI0/XI43/XI15/NET36_XI0/XI43/XI15/MM6_g N_VSS_XI0/XI43/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM7 N_XI0/XI43/XI15/NET36_XI0/XI43/XI15/MM7_d
+ N_XI0/XI43/XI15/NET35_XI0/XI43/XI15/MM7_g N_VSS_XI0/XI43/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM8 N_XI0/XI43/XI15/NET35_XI0/XI43/XI15/MM8_d
+ N_WL<83>_XI0/XI43/XI15/MM8_g N_BLN<0>_XI0/XI43/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI43/XI15/MM5 N_XI0/XI43/XI15/NET34_XI0/XI43/XI15/MM5_d
+ N_XI0/XI43/XI15/NET33_XI0/XI43/XI15/MM5_g N_VDD_XI0/XI43/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI15/MM4 N_XI0/XI43/XI15/NET33_XI0/XI43/XI15/MM4_d
+ N_XI0/XI43/XI15/NET34_XI0/XI43/XI15/MM4_g N_VDD_XI0/XI43/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI15/MM10 N_XI0/XI43/XI15/NET35_XI0/XI43/XI15/MM10_d
+ N_XI0/XI43/XI15/NET36_XI0/XI43/XI15/MM10_g N_VDD_XI0/XI43/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI43/XI15/MM11 N_XI0/XI43/XI15/NET36_XI0/XI43/XI15/MM11_d
+ N_XI0/XI43/XI15/NET35_XI0/XI43/XI15/MM11_g N_VDD_XI0/XI43/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI0/MM2 N_XI0/XI44/XI0/NET34_XI0/XI44/XI0/MM2_d
+ N_XI0/XI44/XI0/NET33_XI0/XI44/XI0/MM2_g N_VSS_XI0/XI44/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM3 N_XI0/XI44/XI0/NET33_XI0/XI44/XI0/MM3_d
+ N_WL<84>_XI0/XI44/XI0/MM3_g N_BLN<15>_XI0/XI44/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM0 N_XI0/XI44/XI0/NET34_XI0/XI44/XI0/MM0_d
+ N_WL<84>_XI0/XI44/XI0/MM0_g N_BL<15>_XI0/XI44/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM1 N_XI0/XI44/XI0/NET33_XI0/XI44/XI0/MM1_d
+ N_XI0/XI44/XI0/NET34_XI0/XI44/XI0/MM1_g N_VSS_XI0/XI44/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM9 N_XI0/XI44/XI0/NET36_XI0/XI44/XI0/MM9_d
+ N_WL<85>_XI0/XI44/XI0/MM9_g N_BL<15>_XI0/XI44/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM6 N_XI0/XI44/XI0/NET35_XI0/XI44/XI0/MM6_d
+ N_XI0/XI44/XI0/NET36_XI0/XI44/XI0/MM6_g N_VSS_XI0/XI44/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM7 N_XI0/XI44/XI0/NET36_XI0/XI44/XI0/MM7_d
+ N_XI0/XI44/XI0/NET35_XI0/XI44/XI0/MM7_g N_VSS_XI0/XI44/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM8 N_XI0/XI44/XI0/NET35_XI0/XI44/XI0/MM8_d
+ N_WL<85>_XI0/XI44/XI0/MM8_g N_BLN<15>_XI0/XI44/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI0/MM5 N_XI0/XI44/XI0/NET34_XI0/XI44/XI0/MM5_d
+ N_XI0/XI44/XI0/NET33_XI0/XI44/XI0/MM5_g N_VDD_XI0/XI44/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI0/MM4 N_XI0/XI44/XI0/NET33_XI0/XI44/XI0/MM4_d
+ N_XI0/XI44/XI0/NET34_XI0/XI44/XI0/MM4_g N_VDD_XI0/XI44/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI0/MM10 N_XI0/XI44/XI0/NET35_XI0/XI44/XI0/MM10_d
+ N_XI0/XI44/XI0/NET36_XI0/XI44/XI0/MM10_g N_VDD_XI0/XI44/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI0/MM11 N_XI0/XI44/XI0/NET36_XI0/XI44/XI0/MM11_d
+ N_XI0/XI44/XI0/NET35_XI0/XI44/XI0/MM11_g N_VDD_XI0/XI44/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI1/MM2 N_XI0/XI44/XI1/NET34_XI0/XI44/XI1/MM2_d
+ N_XI0/XI44/XI1/NET33_XI0/XI44/XI1/MM2_g N_VSS_XI0/XI44/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM3 N_XI0/XI44/XI1/NET33_XI0/XI44/XI1/MM3_d
+ N_WL<84>_XI0/XI44/XI1/MM3_g N_BLN<14>_XI0/XI44/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM0 N_XI0/XI44/XI1/NET34_XI0/XI44/XI1/MM0_d
+ N_WL<84>_XI0/XI44/XI1/MM0_g N_BL<14>_XI0/XI44/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM1 N_XI0/XI44/XI1/NET33_XI0/XI44/XI1/MM1_d
+ N_XI0/XI44/XI1/NET34_XI0/XI44/XI1/MM1_g N_VSS_XI0/XI44/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM9 N_XI0/XI44/XI1/NET36_XI0/XI44/XI1/MM9_d
+ N_WL<85>_XI0/XI44/XI1/MM9_g N_BL<14>_XI0/XI44/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM6 N_XI0/XI44/XI1/NET35_XI0/XI44/XI1/MM6_d
+ N_XI0/XI44/XI1/NET36_XI0/XI44/XI1/MM6_g N_VSS_XI0/XI44/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM7 N_XI0/XI44/XI1/NET36_XI0/XI44/XI1/MM7_d
+ N_XI0/XI44/XI1/NET35_XI0/XI44/XI1/MM7_g N_VSS_XI0/XI44/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM8 N_XI0/XI44/XI1/NET35_XI0/XI44/XI1/MM8_d
+ N_WL<85>_XI0/XI44/XI1/MM8_g N_BLN<14>_XI0/XI44/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI1/MM5 N_XI0/XI44/XI1/NET34_XI0/XI44/XI1/MM5_d
+ N_XI0/XI44/XI1/NET33_XI0/XI44/XI1/MM5_g N_VDD_XI0/XI44/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI1/MM4 N_XI0/XI44/XI1/NET33_XI0/XI44/XI1/MM4_d
+ N_XI0/XI44/XI1/NET34_XI0/XI44/XI1/MM4_g N_VDD_XI0/XI44/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI1/MM10 N_XI0/XI44/XI1/NET35_XI0/XI44/XI1/MM10_d
+ N_XI0/XI44/XI1/NET36_XI0/XI44/XI1/MM10_g N_VDD_XI0/XI44/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI1/MM11 N_XI0/XI44/XI1/NET36_XI0/XI44/XI1/MM11_d
+ N_XI0/XI44/XI1/NET35_XI0/XI44/XI1/MM11_g N_VDD_XI0/XI44/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI2/MM2 N_XI0/XI44/XI2/NET34_XI0/XI44/XI2/MM2_d
+ N_XI0/XI44/XI2/NET33_XI0/XI44/XI2/MM2_g N_VSS_XI0/XI44/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM3 N_XI0/XI44/XI2/NET33_XI0/XI44/XI2/MM3_d
+ N_WL<84>_XI0/XI44/XI2/MM3_g N_BLN<13>_XI0/XI44/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM0 N_XI0/XI44/XI2/NET34_XI0/XI44/XI2/MM0_d
+ N_WL<84>_XI0/XI44/XI2/MM0_g N_BL<13>_XI0/XI44/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM1 N_XI0/XI44/XI2/NET33_XI0/XI44/XI2/MM1_d
+ N_XI0/XI44/XI2/NET34_XI0/XI44/XI2/MM1_g N_VSS_XI0/XI44/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM9 N_XI0/XI44/XI2/NET36_XI0/XI44/XI2/MM9_d
+ N_WL<85>_XI0/XI44/XI2/MM9_g N_BL<13>_XI0/XI44/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM6 N_XI0/XI44/XI2/NET35_XI0/XI44/XI2/MM6_d
+ N_XI0/XI44/XI2/NET36_XI0/XI44/XI2/MM6_g N_VSS_XI0/XI44/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM7 N_XI0/XI44/XI2/NET36_XI0/XI44/XI2/MM7_d
+ N_XI0/XI44/XI2/NET35_XI0/XI44/XI2/MM7_g N_VSS_XI0/XI44/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM8 N_XI0/XI44/XI2/NET35_XI0/XI44/XI2/MM8_d
+ N_WL<85>_XI0/XI44/XI2/MM8_g N_BLN<13>_XI0/XI44/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI2/MM5 N_XI0/XI44/XI2/NET34_XI0/XI44/XI2/MM5_d
+ N_XI0/XI44/XI2/NET33_XI0/XI44/XI2/MM5_g N_VDD_XI0/XI44/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI2/MM4 N_XI0/XI44/XI2/NET33_XI0/XI44/XI2/MM4_d
+ N_XI0/XI44/XI2/NET34_XI0/XI44/XI2/MM4_g N_VDD_XI0/XI44/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI2/MM10 N_XI0/XI44/XI2/NET35_XI0/XI44/XI2/MM10_d
+ N_XI0/XI44/XI2/NET36_XI0/XI44/XI2/MM10_g N_VDD_XI0/XI44/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI2/MM11 N_XI0/XI44/XI2/NET36_XI0/XI44/XI2/MM11_d
+ N_XI0/XI44/XI2/NET35_XI0/XI44/XI2/MM11_g N_VDD_XI0/XI44/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI3/MM2 N_XI0/XI44/XI3/NET34_XI0/XI44/XI3/MM2_d
+ N_XI0/XI44/XI3/NET33_XI0/XI44/XI3/MM2_g N_VSS_XI0/XI44/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM3 N_XI0/XI44/XI3/NET33_XI0/XI44/XI3/MM3_d
+ N_WL<84>_XI0/XI44/XI3/MM3_g N_BLN<12>_XI0/XI44/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM0 N_XI0/XI44/XI3/NET34_XI0/XI44/XI3/MM0_d
+ N_WL<84>_XI0/XI44/XI3/MM0_g N_BL<12>_XI0/XI44/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM1 N_XI0/XI44/XI3/NET33_XI0/XI44/XI3/MM1_d
+ N_XI0/XI44/XI3/NET34_XI0/XI44/XI3/MM1_g N_VSS_XI0/XI44/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM9 N_XI0/XI44/XI3/NET36_XI0/XI44/XI3/MM9_d
+ N_WL<85>_XI0/XI44/XI3/MM9_g N_BL<12>_XI0/XI44/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM6 N_XI0/XI44/XI3/NET35_XI0/XI44/XI3/MM6_d
+ N_XI0/XI44/XI3/NET36_XI0/XI44/XI3/MM6_g N_VSS_XI0/XI44/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM7 N_XI0/XI44/XI3/NET36_XI0/XI44/XI3/MM7_d
+ N_XI0/XI44/XI3/NET35_XI0/XI44/XI3/MM7_g N_VSS_XI0/XI44/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM8 N_XI0/XI44/XI3/NET35_XI0/XI44/XI3/MM8_d
+ N_WL<85>_XI0/XI44/XI3/MM8_g N_BLN<12>_XI0/XI44/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI3/MM5 N_XI0/XI44/XI3/NET34_XI0/XI44/XI3/MM5_d
+ N_XI0/XI44/XI3/NET33_XI0/XI44/XI3/MM5_g N_VDD_XI0/XI44/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI3/MM4 N_XI0/XI44/XI3/NET33_XI0/XI44/XI3/MM4_d
+ N_XI0/XI44/XI3/NET34_XI0/XI44/XI3/MM4_g N_VDD_XI0/XI44/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI3/MM10 N_XI0/XI44/XI3/NET35_XI0/XI44/XI3/MM10_d
+ N_XI0/XI44/XI3/NET36_XI0/XI44/XI3/MM10_g N_VDD_XI0/XI44/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI3/MM11 N_XI0/XI44/XI3/NET36_XI0/XI44/XI3/MM11_d
+ N_XI0/XI44/XI3/NET35_XI0/XI44/XI3/MM11_g N_VDD_XI0/XI44/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI4/MM2 N_XI0/XI44/XI4/NET34_XI0/XI44/XI4/MM2_d
+ N_XI0/XI44/XI4/NET33_XI0/XI44/XI4/MM2_g N_VSS_XI0/XI44/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM3 N_XI0/XI44/XI4/NET33_XI0/XI44/XI4/MM3_d
+ N_WL<84>_XI0/XI44/XI4/MM3_g N_BLN<11>_XI0/XI44/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM0 N_XI0/XI44/XI4/NET34_XI0/XI44/XI4/MM0_d
+ N_WL<84>_XI0/XI44/XI4/MM0_g N_BL<11>_XI0/XI44/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM1 N_XI0/XI44/XI4/NET33_XI0/XI44/XI4/MM1_d
+ N_XI0/XI44/XI4/NET34_XI0/XI44/XI4/MM1_g N_VSS_XI0/XI44/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM9 N_XI0/XI44/XI4/NET36_XI0/XI44/XI4/MM9_d
+ N_WL<85>_XI0/XI44/XI4/MM9_g N_BL<11>_XI0/XI44/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM6 N_XI0/XI44/XI4/NET35_XI0/XI44/XI4/MM6_d
+ N_XI0/XI44/XI4/NET36_XI0/XI44/XI4/MM6_g N_VSS_XI0/XI44/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM7 N_XI0/XI44/XI4/NET36_XI0/XI44/XI4/MM7_d
+ N_XI0/XI44/XI4/NET35_XI0/XI44/XI4/MM7_g N_VSS_XI0/XI44/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM8 N_XI0/XI44/XI4/NET35_XI0/XI44/XI4/MM8_d
+ N_WL<85>_XI0/XI44/XI4/MM8_g N_BLN<11>_XI0/XI44/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI4/MM5 N_XI0/XI44/XI4/NET34_XI0/XI44/XI4/MM5_d
+ N_XI0/XI44/XI4/NET33_XI0/XI44/XI4/MM5_g N_VDD_XI0/XI44/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI4/MM4 N_XI0/XI44/XI4/NET33_XI0/XI44/XI4/MM4_d
+ N_XI0/XI44/XI4/NET34_XI0/XI44/XI4/MM4_g N_VDD_XI0/XI44/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI4/MM10 N_XI0/XI44/XI4/NET35_XI0/XI44/XI4/MM10_d
+ N_XI0/XI44/XI4/NET36_XI0/XI44/XI4/MM10_g N_VDD_XI0/XI44/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI4/MM11 N_XI0/XI44/XI4/NET36_XI0/XI44/XI4/MM11_d
+ N_XI0/XI44/XI4/NET35_XI0/XI44/XI4/MM11_g N_VDD_XI0/XI44/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI5/MM2 N_XI0/XI44/XI5/NET34_XI0/XI44/XI5/MM2_d
+ N_XI0/XI44/XI5/NET33_XI0/XI44/XI5/MM2_g N_VSS_XI0/XI44/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM3 N_XI0/XI44/XI5/NET33_XI0/XI44/XI5/MM3_d
+ N_WL<84>_XI0/XI44/XI5/MM3_g N_BLN<10>_XI0/XI44/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM0 N_XI0/XI44/XI5/NET34_XI0/XI44/XI5/MM0_d
+ N_WL<84>_XI0/XI44/XI5/MM0_g N_BL<10>_XI0/XI44/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM1 N_XI0/XI44/XI5/NET33_XI0/XI44/XI5/MM1_d
+ N_XI0/XI44/XI5/NET34_XI0/XI44/XI5/MM1_g N_VSS_XI0/XI44/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM9 N_XI0/XI44/XI5/NET36_XI0/XI44/XI5/MM9_d
+ N_WL<85>_XI0/XI44/XI5/MM9_g N_BL<10>_XI0/XI44/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM6 N_XI0/XI44/XI5/NET35_XI0/XI44/XI5/MM6_d
+ N_XI0/XI44/XI5/NET36_XI0/XI44/XI5/MM6_g N_VSS_XI0/XI44/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM7 N_XI0/XI44/XI5/NET36_XI0/XI44/XI5/MM7_d
+ N_XI0/XI44/XI5/NET35_XI0/XI44/XI5/MM7_g N_VSS_XI0/XI44/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM8 N_XI0/XI44/XI5/NET35_XI0/XI44/XI5/MM8_d
+ N_WL<85>_XI0/XI44/XI5/MM8_g N_BLN<10>_XI0/XI44/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI5/MM5 N_XI0/XI44/XI5/NET34_XI0/XI44/XI5/MM5_d
+ N_XI0/XI44/XI5/NET33_XI0/XI44/XI5/MM5_g N_VDD_XI0/XI44/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI5/MM4 N_XI0/XI44/XI5/NET33_XI0/XI44/XI5/MM4_d
+ N_XI0/XI44/XI5/NET34_XI0/XI44/XI5/MM4_g N_VDD_XI0/XI44/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI5/MM10 N_XI0/XI44/XI5/NET35_XI0/XI44/XI5/MM10_d
+ N_XI0/XI44/XI5/NET36_XI0/XI44/XI5/MM10_g N_VDD_XI0/XI44/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI5/MM11 N_XI0/XI44/XI5/NET36_XI0/XI44/XI5/MM11_d
+ N_XI0/XI44/XI5/NET35_XI0/XI44/XI5/MM11_g N_VDD_XI0/XI44/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI6/MM2 N_XI0/XI44/XI6/NET34_XI0/XI44/XI6/MM2_d
+ N_XI0/XI44/XI6/NET33_XI0/XI44/XI6/MM2_g N_VSS_XI0/XI44/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM3 N_XI0/XI44/XI6/NET33_XI0/XI44/XI6/MM3_d
+ N_WL<84>_XI0/XI44/XI6/MM3_g N_BLN<9>_XI0/XI44/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM0 N_XI0/XI44/XI6/NET34_XI0/XI44/XI6/MM0_d
+ N_WL<84>_XI0/XI44/XI6/MM0_g N_BL<9>_XI0/XI44/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM1 N_XI0/XI44/XI6/NET33_XI0/XI44/XI6/MM1_d
+ N_XI0/XI44/XI6/NET34_XI0/XI44/XI6/MM1_g N_VSS_XI0/XI44/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM9 N_XI0/XI44/XI6/NET36_XI0/XI44/XI6/MM9_d
+ N_WL<85>_XI0/XI44/XI6/MM9_g N_BL<9>_XI0/XI44/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM6 N_XI0/XI44/XI6/NET35_XI0/XI44/XI6/MM6_d
+ N_XI0/XI44/XI6/NET36_XI0/XI44/XI6/MM6_g N_VSS_XI0/XI44/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM7 N_XI0/XI44/XI6/NET36_XI0/XI44/XI6/MM7_d
+ N_XI0/XI44/XI6/NET35_XI0/XI44/XI6/MM7_g N_VSS_XI0/XI44/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM8 N_XI0/XI44/XI6/NET35_XI0/XI44/XI6/MM8_d
+ N_WL<85>_XI0/XI44/XI6/MM8_g N_BLN<9>_XI0/XI44/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI6/MM5 N_XI0/XI44/XI6/NET34_XI0/XI44/XI6/MM5_d
+ N_XI0/XI44/XI6/NET33_XI0/XI44/XI6/MM5_g N_VDD_XI0/XI44/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI6/MM4 N_XI0/XI44/XI6/NET33_XI0/XI44/XI6/MM4_d
+ N_XI0/XI44/XI6/NET34_XI0/XI44/XI6/MM4_g N_VDD_XI0/XI44/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI6/MM10 N_XI0/XI44/XI6/NET35_XI0/XI44/XI6/MM10_d
+ N_XI0/XI44/XI6/NET36_XI0/XI44/XI6/MM10_g N_VDD_XI0/XI44/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI6/MM11 N_XI0/XI44/XI6/NET36_XI0/XI44/XI6/MM11_d
+ N_XI0/XI44/XI6/NET35_XI0/XI44/XI6/MM11_g N_VDD_XI0/XI44/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI7/MM2 N_XI0/XI44/XI7/NET34_XI0/XI44/XI7/MM2_d
+ N_XI0/XI44/XI7/NET33_XI0/XI44/XI7/MM2_g N_VSS_XI0/XI44/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM3 N_XI0/XI44/XI7/NET33_XI0/XI44/XI7/MM3_d
+ N_WL<84>_XI0/XI44/XI7/MM3_g N_BLN<8>_XI0/XI44/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM0 N_XI0/XI44/XI7/NET34_XI0/XI44/XI7/MM0_d
+ N_WL<84>_XI0/XI44/XI7/MM0_g N_BL<8>_XI0/XI44/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM1 N_XI0/XI44/XI7/NET33_XI0/XI44/XI7/MM1_d
+ N_XI0/XI44/XI7/NET34_XI0/XI44/XI7/MM1_g N_VSS_XI0/XI44/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM9 N_XI0/XI44/XI7/NET36_XI0/XI44/XI7/MM9_d
+ N_WL<85>_XI0/XI44/XI7/MM9_g N_BL<8>_XI0/XI44/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM6 N_XI0/XI44/XI7/NET35_XI0/XI44/XI7/MM6_d
+ N_XI0/XI44/XI7/NET36_XI0/XI44/XI7/MM6_g N_VSS_XI0/XI44/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM7 N_XI0/XI44/XI7/NET36_XI0/XI44/XI7/MM7_d
+ N_XI0/XI44/XI7/NET35_XI0/XI44/XI7/MM7_g N_VSS_XI0/XI44/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM8 N_XI0/XI44/XI7/NET35_XI0/XI44/XI7/MM8_d
+ N_WL<85>_XI0/XI44/XI7/MM8_g N_BLN<8>_XI0/XI44/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI7/MM5 N_XI0/XI44/XI7/NET34_XI0/XI44/XI7/MM5_d
+ N_XI0/XI44/XI7/NET33_XI0/XI44/XI7/MM5_g N_VDD_XI0/XI44/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI7/MM4 N_XI0/XI44/XI7/NET33_XI0/XI44/XI7/MM4_d
+ N_XI0/XI44/XI7/NET34_XI0/XI44/XI7/MM4_g N_VDD_XI0/XI44/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI7/MM10 N_XI0/XI44/XI7/NET35_XI0/XI44/XI7/MM10_d
+ N_XI0/XI44/XI7/NET36_XI0/XI44/XI7/MM10_g N_VDD_XI0/XI44/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI7/MM11 N_XI0/XI44/XI7/NET36_XI0/XI44/XI7/MM11_d
+ N_XI0/XI44/XI7/NET35_XI0/XI44/XI7/MM11_g N_VDD_XI0/XI44/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI8/MM2 N_XI0/XI44/XI8/NET34_XI0/XI44/XI8/MM2_d
+ N_XI0/XI44/XI8/NET33_XI0/XI44/XI8/MM2_g N_VSS_XI0/XI44/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM3 N_XI0/XI44/XI8/NET33_XI0/XI44/XI8/MM3_d
+ N_WL<84>_XI0/XI44/XI8/MM3_g N_BLN<7>_XI0/XI44/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM0 N_XI0/XI44/XI8/NET34_XI0/XI44/XI8/MM0_d
+ N_WL<84>_XI0/XI44/XI8/MM0_g N_BL<7>_XI0/XI44/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM1 N_XI0/XI44/XI8/NET33_XI0/XI44/XI8/MM1_d
+ N_XI0/XI44/XI8/NET34_XI0/XI44/XI8/MM1_g N_VSS_XI0/XI44/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM9 N_XI0/XI44/XI8/NET36_XI0/XI44/XI8/MM9_d
+ N_WL<85>_XI0/XI44/XI8/MM9_g N_BL<7>_XI0/XI44/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM6 N_XI0/XI44/XI8/NET35_XI0/XI44/XI8/MM6_d
+ N_XI0/XI44/XI8/NET36_XI0/XI44/XI8/MM6_g N_VSS_XI0/XI44/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM7 N_XI0/XI44/XI8/NET36_XI0/XI44/XI8/MM7_d
+ N_XI0/XI44/XI8/NET35_XI0/XI44/XI8/MM7_g N_VSS_XI0/XI44/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM8 N_XI0/XI44/XI8/NET35_XI0/XI44/XI8/MM8_d
+ N_WL<85>_XI0/XI44/XI8/MM8_g N_BLN<7>_XI0/XI44/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI8/MM5 N_XI0/XI44/XI8/NET34_XI0/XI44/XI8/MM5_d
+ N_XI0/XI44/XI8/NET33_XI0/XI44/XI8/MM5_g N_VDD_XI0/XI44/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI8/MM4 N_XI0/XI44/XI8/NET33_XI0/XI44/XI8/MM4_d
+ N_XI0/XI44/XI8/NET34_XI0/XI44/XI8/MM4_g N_VDD_XI0/XI44/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI8/MM10 N_XI0/XI44/XI8/NET35_XI0/XI44/XI8/MM10_d
+ N_XI0/XI44/XI8/NET36_XI0/XI44/XI8/MM10_g N_VDD_XI0/XI44/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI8/MM11 N_XI0/XI44/XI8/NET36_XI0/XI44/XI8/MM11_d
+ N_XI0/XI44/XI8/NET35_XI0/XI44/XI8/MM11_g N_VDD_XI0/XI44/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI9/MM2 N_XI0/XI44/XI9/NET34_XI0/XI44/XI9/MM2_d
+ N_XI0/XI44/XI9/NET33_XI0/XI44/XI9/MM2_g N_VSS_XI0/XI44/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM3 N_XI0/XI44/XI9/NET33_XI0/XI44/XI9/MM3_d
+ N_WL<84>_XI0/XI44/XI9/MM3_g N_BLN<6>_XI0/XI44/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM0 N_XI0/XI44/XI9/NET34_XI0/XI44/XI9/MM0_d
+ N_WL<84>_XI0/XI44/XI9/MM0_g N_BL<6>_XI0/XI44/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM1 N_XI0/XI44/XI9/NET33_XI0/XI44/XI9/MM1_d
+ N_XI0/XI44/XI9/NET34_XI0/XI44/XI9/MM1_g N_VSS_XI0/XI44/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM9 N_XI0/XI44/XI9/NET36_XI0/XI44/XI9/MM9_d
+ N_WL<85>_XI0/XI44/XI9/MM9_g N_BL<6>_XI0/XI44/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM6 N_XI0/XI44/XI9/NET35_XI0/XI44/XI9/MM6_d
+ N_XI0/XI44/XI9/NET36_XI0/XI44/XI9/MM6_g N_VSS_XI0/XI44/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM7 N_XI0/XI44/XI9/NET36_XI0/XI44/XI9/MM7_d
+ N_XI0/XI44/XI9/NET35_XI0/XI44/XI9/MM7_g N_VSS_XI0/XI44/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM8 N_XI0/XI44/XI9/NET35_XI0/XI44/XI9/MM8_d
+ N_WL<85>_XI0/XI44/XI9/MM8_g N_BLN<6>_XI0/XI44/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI9/MM5 N_XI0/XI44/XI9/NET34_XI0/XI44/XI9/MM5_d
+ N_XI0/XI44/XI9/NET33_XI0/XI44/XI9/MM5_g N_VDD_XI0/XI44/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI9/MM4 N_XI0/XI44/XI9/NET33_XI0/XI44/XI9/MM4_d
+ N_XI0/XI44/XI9/NET34_XI0/XI44/XI9/MM4_g N_VDD_XI0/XI44/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI9/MM10 N_XI0/XI44/XI9/NET35_XI0/XI44/XI9/MM10_d
+ N_XI0/XI44/XI9/NET36_XI0/XI44/XI9/MM10_g N_VDD_XI0/XI44/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI9/MM11 N_XI0/XI44/XI9/NET36_XI0/XI44/XI9/MM11_d
+ N_XI0/XI44/XI9/NET35_XI0/XI44/XI9/MM11_g N_VDD_XI0/XI44/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI10/MM2 N_XI0/XI44/XI10/NET34_XI0/XI44/XI10/MM2_d
+ N_XI0/XI44/XI10/NET33_XI0/XI44/XI10/MM2_g N_VSS_XI0/XI44/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM3 N_XI0/XI44/XI10/NET33_XI0/XI44/XI10/MM3_d
+ N_WL<84>_XI0/XI44/XI10/MM3_g N_BLN<5>_XI0/XI44/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM0 N_XI0/XI44/XI10/NET34_XI0/XI44/XI10/MM0_d
+ N_WL<84>_XI0/XI44/XI10/MM0_g N_BL<5>_XI0/XI44/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM1 N_XI0/XI44/XI10/NET33_XI0/XI44/XI10/MM1_d
+ N_XI0/XI44/XI10/NET34_XI0/XI44/XI10/MM1_g N_VSS_XI0/XI44/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM9 N_XI0/XI44/XI10/NET36_XI0/XI44/XI10/MM9_d
+ N_WL<85>_XI0/XI44/XI10/MM9_g N_BL<5>_XI0/XI44/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM6 N_XI0/XI44/XI10/NET35_XI0/XI44/XI10/MM6_d
+ N_XI0/XI44/XI10/NET36_XI0/XI44/XI10/MM6_g N_VSS_XI0/XI44/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM7 N_XI0/XI44/XI10/NET36_XI0/XI44/XI10/MM7_d
+ N_XI0/XI44/XI10/NET35_XI0/XI44/XI10/MM7_g N_VSS_XI0/XI44/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM8 N_XI0/XI44/XI10/NET35_XI0/XI44/XI10/MM8_d
+ N_WL<85>_XI0/XI44/XI10/MM8_g N_BLN<5>_XI0/XI44/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI10/MM5 N_XI0/XI44/XI10/NET34_XI0/XI44/XI10/MM5_d
+ N_XI0/XI44/XI10/NET33_XI0/XI44/XI10/MM5_g N_VDD_XI0/XI44/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI10/MM4 N_XI0/XI44/XI10/NET33_XI0/XI44/XI10/MM4_d
+ N_XI0/XI44/XI10/NET34_XI0/XI44/XI10/MM4_g N_VDD_XI0/XI44/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI10/MM10 N_XI0/XI44/XI10/NET35_XI0/XI44/XI10/MM10_d
+ N_XI0/XI44/XI10/NET36_XI0/XI44/XI10/MM10_g N_VDD_XI0/XI44/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI10/MM11 N_XI0/XI44/XI10/NET36_XI0/XI44/XI10/MM11_d
+ N_XI0/XI44/XI10/NET35_XI0/XI44/XI10/MM11_g N_VDD_XI0/XI44/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI11/MM2 N_XI0/XI44/XI11/NET34_XI0/XI44/XI11/MM2_d
+ N_XI0/XI44/XI11/NET33_XI0/XI44/XI11/MM2_g N_VSS_XI0/XI44/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM3 N_XI0/XI44/XI11/NET33_XI0/XI44/XI11/MM3_d
+ N_WL<84>_XI0/XI44/XI11/MM3_g N_BLN<4>_XI0/XI44/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM0 N_XI0/XI44/XI11/NET34_XI0/XI44/XI11/MM0_d
+ N_WL<84>_XI0/XI44/XI11/MM0_g N_BL<4>_XI0/XI44/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM1 N_XI0/XI44/XI11/NET33_XI0/XI44/XI11/MM1_d
+ N_XI0/XI44/XI11/NET34_XI0/XI44/XI11/MM1_g N_VSS_XI0/XI44/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM9 N_XI0/XI44/XI11/NET36_XI0/XI44/XI11/MM9_d
+ N_WL<85>_XI0/XI44/XI11/MM9_g N_BL<4>_XI0/XI44/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM6 N_XI0/XI44/XI11/NET35_XI0/XI44/XI11/MM6_d
+ N_XI0/XI44/XI11/NET36_XI0/XI44/XI11/MM6_g N_VSS_XI0/XI44/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM7 N_XI0/XI44/XI11/NET36_XI0/XI44/XI11/MM7_d
+ N_XI0/XI44/XI11/NET35_XI0/XI44/XI11/MM7_g N_VSS_XI0/XI44/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM8 N_XI0/XI44/XI11/NET35_XI0/XI44/XI11/MM8_d
+ N_WL<85>_XI0/XI44/XI11/MM8_g N_BLN<4>_XI0/XI44/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI11/MM5 N_XI0/XI44/XI11/NET34_XI0/XI44/XI11/MM5_d
+ N_XI0/XI44/XI11/NET33_XI0/XI44/XI11/MM5_g N_VDD_XI0/XI44/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI11/MM4 N_XI0/XI44/XI11/NET33_XI0/XI44/XI11/MM4_d
+ N_XI0/XI44/XI11/NET34_XI0/XI44/XI11/MM4_g N_VDD_XI0/XI44/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI11/MM10 N_XI0/XI44/XI11/NET35_XI0/XI44/XI11/MM10_d
+ N_XI0/XI44/XI11/NET36_XI0/XI44/XI11/MM10_g N_VDD_XI0/XI44/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI11/MM11 N_XI0/XI44/XI11/NET36_XI0/XI44/XI11/MM11_d
+ N_XI0/XI44/XI11/NET35_XI0/XI44/XI11/MM11_g N_VDD_XI0/XI44/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI12/MM2 N_XI0/XI44/XI12/NET34_XI0/XI44/XI12/MM2_d
+ N_XI0/XI44/XI12/NET33_XI0/XI44/XI12/MM2_g N_VSS_XI0/XI44/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM3 N_XI0/XI44/XI12/NET33_XI0/XI44/XI12/MM3_d
+ N_WL<84>_XI0/XI44/XI12/MM3_g N_BLN<3>_XI0/XI44/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM0 N_XI0/XI44/XI12/NET34_XI0/XI44/XI12/MM0_d
+ N_WL<84>_XI0/XI44/XI12/MM0_g N_BL<3>_XI0/XI44/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM1 N_XI0/XI44/XI12/NET33_XI0/XI44/XI12/MM1_d
+ N_XI0/XI44/XI12/NET34_XI0/XI44/XI12/MM1_g N_VSS_XI0/XI44/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM9 N_XI0/XI44/XI12/NET36_XI0/XI44/XI12/MM9_d
+ N_WL<85>_XI0/XI44/XI12/MM9_g N_BL<3>_XI0/XI44/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM6 N_XI0/XI44/XI12/NET35_XI0/XI44/XI12/MM6_d
+ N_XI0/XI44/XI12/NET36_XI0/XI44/XI12/MM6_g N_VSS_XI0/XI44/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM7 N_XI0/XI44/XI12/NET36_XI0/XI44/XI12/MM7_d
+ N_XI0/XI44/XI12/NET35_XI0/XI44/XI12/MM7_g N_VSS_XI0/XI44/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM8 N_XI0/XI44/XI12/NET35_XI0/XI44/XI12/MM8_d
+ N_WL<85>_XI0/XI44/XI12/MM8_g N_BLN<3>_XI0/XI44/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI12/MM5 N_XI0/XI44/XI12/NET34_XI0/XI44/XI12/MM5_d
+ N_XI0/XI44/XI12/NET33_XI0/XI44/XI12/MM5_g N_VDD_XI0/XI44/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI12/MM4 N_XI0/XI44/XI12/NET33_XI0/XI44/XI12/MM4_d
+ N_XI0/XI44/XI12/NET34_XI0/XI44/XI12/MM4_g N_VDD_XI0/XI44/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI12/MM10 N_XI0/XI44/XI12/NET35_XI0/XI44/XI12/MM10_d
+ N_XI0/XI44/XI12/NET36_XI0/XI44/XI12/MM10_g N_VDD_XI0/XI44/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI12/MM11 N_XI0/XI44/XI12/NET36_XI0/XI44/XI12/MM11_d
+ N_XI0/XI44/XI12/NET35_XI0/XI44/XI12/MM11_g N_VDD_XI0/XI44/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI13/MM2 N_XI0/XI44/XI13/NET34_XI0/XI44/XI13/MM2_d
+ N_XI0/XI44/XI13/NET33_XI0/XI44/XI13/MM2_g N_VSS_XI0/XI44/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM3 N_XI0/XI44/XI13/NET33_XI0/XI44/XI13/MM3_d
+ N_WL<84>_XI0/XI44/XI13/MM3_g N_BLN<2>_XI0/XI44/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM0 N_XI0/XI44/XI13/NET34_XI0/XI44/XI13/MM0_d
+ N_WL<84>_XI0/XI44/XI13/MM0_g N_BL<2>_XI0/XI44/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM1 N_XI0/XI44/XI13/NET33_XI0/XI44/XI13/MM1_d
+ N_XI0/XI44/XI13/NET34_XI0/XI44/XI13/MM1_g N_VSS_XI0/XI44/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM9 N_XI0/XI44/XI13/NET36_XI0/XI44/XI13/MM9_d
+ N_WL<85>_XI0/XI44/XI13/MM9_g N_BL<2>_XI0/XI44/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM6 N_XI0/XI44/XI13/NET35_XI0/XI44/XI13/MM6_d
+ N_XI0/XI44/XI13/NET36_XI0/XI44/XI13/MM6_g N_VSS_XI0/XI44/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM7 N_XI0/XI44/XI13/NET36_XI0/XI44/XI13/MM7_d
+ N_XI0/XI44/XI13/NET35_XI0/XI44/XI13/MM7_g N_VSS_XI0/XI44/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM8 N_XI0/XI44/XI13/NET35_XI0/XI44/XI13/MM8_d
+ N_WL<85>_XI0/XI44/XI13/MM8_g N_BLN<2>_XI0/XI44/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI13/MM5 N_XI0/XI44/XI13/NET34_XI0/XI44/XI13/MM5_d
+ N_XI0/XI44/XI13/NET33_XI0/XI44/XI13/MM5_g N_VDD_XI0/XI44/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI13/MM4 N_XI0/XI44/XI13/NET33_XI0/XI44/XI13/MM4_d
+ N_XI0/XI44/XI13/NET34_XI0/XI44/XI13/MM4_g N_VDD_XI0/XI44/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI13/MM10 N_XI0/XI44/XI13/NET35_XI0/XI44/XI13/MM10_d
+ N_XI0/XI44/XI13/NET36_XI0/XI44/XI13/MM10_g N_VDD_XI0/XI44/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI13/MM11 N_XI0/XI44/XI13/NET36_XI0/XI44/XI13/MM11_d
+ N_XI0/XI44/XI13/NET35_XI0/XI44/XI13/MM11_g N_VDD_XI0/XI44/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI14/MM2 N_XI0/XI44/XI14/NET34_XI0/XI44/XI14/MM2_d
+ N_XI0/XI44/XI14/NET33_XI0/XI44/XI14/MM2_g N_VSS_XI0/XI44/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM3 N_XI0/XI44/XI14/NET33_XI0/XI44/XI14/MM3_d
+ N_WL<84>_XI0/XI44/XI14/MM3_g N_BLN<1>_XI0/XI44/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM0 N_XI0/XI44/XI14/NET34_XI0/XI44/XI14/MM0_d
+ N_WL<84>_XI0/XI44/XI14/MM0_g N_BL<1>_XI0/XI44/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM1 N_XI0/XI44/XI14/NET33_XI0/XI44/XI14/MM1_d
+ N_XI0/XI44/XI14/NET34_XI0/XI44/XI14/MM1_g N_VSS_XI0/XI44/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM9 N_XI0/XI44/XI14/NET36_XI0/XI44/XI14/MM9_d
+ N_WL<85>_XI0/XI44/XI14/MM9_g N_BL<1>_XI0/XI44/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM6 N_XI0/XI44/XI14/NET35_XI0/XI44/XI14/MM6_d
+ N_XI0/XI44/XI14/NET36_XI0/XI44/XI14/MM6_g N_VSS_XI0/XI44/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM7 N_XI0/XI44/XI14/NET36_XI0/XI44/XI14/MM7_d
+ N_XI0/XI44/XI14/NET35_XI0/XI44/XI14/MM7_g N_VSS_XI0/XI44/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM8 N_XI0/XI44/XI14/NET35_XI0/XI44/XI14/MM8_d
+ N_WL<85>_XI0/XI44/XI14/MM8_g N_BLN<1>_XI0/XI44/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI14/MM5 N_XI0/XI44/XI14/NET34_XI0/XI44/XI14/MM5_d
+ N_XI0/XI44/XI14/NET33_XI0/XI44/XI14/MM5_g N_VDD_XI0/XI44/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI14/MM4 N_XI0/XI44/XI14/NET33_XI0/XI44/XI14/MM4_d
+ N_XI0/XI44/XI14/NET34_XI0/XI44/XI14/MM4_g N_VDD_XI0/XI44/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI14/MM10 N_XI0/XI44/XI14/NET35_XI0/XI44/XI14/MM10_d
+ N_XI0/XI44/XI14/NET36_XI0/XI44/XI14/MM10_g N_VDD_XI0/XI44/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI14/MM11 N_XI0/XI44/XI14/NET36_XI0/XI44/XI14/MM11_d
+ N_XI0/XI44/XI14/NET35_XI0/XI44/XI14/MM11_g N_VDD_XI0/XI44/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI15/MM2 N_XI0/XI44/XI15/NET34_XI0/XI44/XI15/MM2_d
+ N_XI0/XI44/XI15/NET33_XI0/XI44/XI15/MM2_g N_VSS_XI0/XI44/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM3 N_XI0/XI44/XI15/NET33_XI0/XI44/XI15/MM3_d
+ N_WL<84>_XI0/XI44/XI15/MM3_g N_BLN<0>_XI0/XI44/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM0 N_XI0/XI44/XI15/NET34_XI0/XI44/XI15/MM0_d
+ N_WL<84>_XI0/XI44/XI15/MM0_g N_BL<0>_XI0/XI44/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM1 N_XI0/XI44/XI15/NET33_XI0/XI44/XI15/MM1_d
+ N_XI0/XI44/XI15/NET34_XI0/XI44/XI15/MM1_g N_VSS_XI0/XI44/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM9 N_XI0/XI44/XI15/NET36_XI0/XI44/XI15/MM9_d
+ N_WL<85>_XI0/XI44/XI15/MM9_g N_BL<0>_XI0/XI44/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM6 N_XI0/XI44/XI15/NET35_XI0/XI44/XI15/MM6_d
+ N_XI0/XI44/XI15/NET36_XI0/XI44/XI15/MM6_g N_VSS_XI0/XI44/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM7 N_XI0/XI44/XI15/NET36_XI0/XI44/XI15/MM7_d
+ N_XI0/XI44/XI15/NET35_XI0/XI44/XI15/MM7_g N_VSS_XI0/XI44/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM8 N_XI0/XI44/XI15/NET35_XI0/XI44/XI15/MM8_d
+ N_WL<85>_XI0/XI44/XI15/MM8_g N_BLN<0>_XI0/XI44/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI44/XI15/MM5 N_XI0/XI44/XI15/NET34_XI0/XI44/XI15/MM5_d
+ N_XI0/XI44/XI15/NET33_XI0/XI44/XI15/MM5_g N_VDD_XI0/XI44/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI15/MM4 N_XI0/XI44/XI15/NET33_XI0/XI44/XI15/MM4_d
+ N_XI0/XI44/XI15/NET34_XI0/XI44/XI15/MM4_g N_VDD_XI0/XI44/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI15/MM10 N_XI0/XI44/XI15/NET35_XI0/XI44/XI15/MM10_d
+ N_XI0/XI44/XI15/NET36_XI0/XI44/XI15/MM10_g N_VDD_XI0/XI44/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI44/XI15/MM11 N_XI0/XI44/XI15/NET36_XI0/XI44/XI15/MM11_d
+ N_XI0/XI44/XI15/NET35_XI0/XI44/XI15/MM11_g N_VDD_XI0/XI44/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI0/MM2 N_XI0/XI45/XI0/NET34_XI0/XI45/XI0/MM2_d
+ N_XI0/XI45/XI0/NET33_XI0/XI45/XI0/MM2_g N_VSS_XI0/XI45/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM3 N_XI0/XI45/XI0/NET33_XI0/XI45/XI0/MM3_d
+ N_WL<86>_XI0/XI45/XI0/MM3_g N_BLN<15>_XI0/XI45/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM0 N_XI0/XI45/XI0/NET34_XI0/XI45/XI0/MM0_d
+ N_WL<86>_XI0/XI45/XI0/MM0_g N_BL<15>_XI0/XI45/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM1 N_XI0/XI45/XI0/NET33_XI0/XI45/XI0/MM1_d
+ N_XI0/XI45/XI0/NET34_XI0/XI45/XI0/MM1_g N_VSS_XI0/XI45/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM9 N_XI0/XI45/XI0/NET36_XI0/XI45/XI0/MM9_d
+ N_WL<87>_XI0/XI45/XI0/MM9_g N_BL<15>_XI0/XI45/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM6 N_XI0/XI45/XI0/NET35_XI0/XI45/XI0/MM6_d
+ N_XI0/XI45/XI0/NET36_XI0/XI45/XI0/MM6_g N_VSS_XI0/XI45/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM7 N_XI0/XI45/XI0/NET36_XI0/XI45/XI0/MM7_d
+ N_XI0/XI45/XI0/NET35_XI0/XI45/XI0/MM7_g N_VSS_XI0/XI45/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM8 N_XI0/XI45/XI0/NET35_XI0/XI45/XI0/MM8_d
+ N_WL<87>_XI0/XI45/XI0/MM8_g N_BLN<15>_XI0/XI45/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI0/MM5 N_XI0/XI45/XI0/NET34_XI0/XI45/XI0/MM5_d
+ N_XI0/XI45/XI0/NET33_XI0/XI45/XI0/MM5_g N_VDD_XI0/XI45/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI0/MM4 N_XI0/XI45/XI0/NET33_XI0/XI45/XI0/MM4_d
+ N_XI0/XI45/XI0/NET34_XI0/XI45/XI0/MM4_g N_VDD_XI0/XI45/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI0/MM10 N_XI0/XI45/XI0/NET35_XI0/XI45/XI0/MM10_d
+ N_XI0/XI45/XI0/NET36_XI0/XI45/XI0/MM10_g N_VDD_XI0/XI45/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI0/MM11 N_XI0/XI45/XI0/NET36_XI0/XI45/XI0/MM11_d
+ N_XI0/XI45/XI0/NET35_XI0/XI45/XI0/MM11_g N_VDD_XI0/XI45/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI1/MM2 N_XI0/XI45/XI1/NET34_XI0/XI45/XI1/MM2_d
+ N_XI0/XI45/XI1/NET33_XI0/XI45/XI1/MM2_g N_VSS_XI0/XI45/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM3 N_XI0/XI45/XI1/NET33_XI0/XI45/XI1/MM3_d
+ N_WL<86>_XI0/XI45/XI1/MM3_g N_BLN<14>_XI0/XI45/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM0 N_XI0/XI45/XI1/NET34_XI0/XI45/XI1/MM0_d
+ N_WL<86>_XI0/XI45/XI1/MM0_g N_BL<14>_XI0/XI45/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM1 N_XI0/XI45/XI1/NET33_XI0/XI45/XI1/MM1_d
+ N_XI0/XI45/XI1/NET34_XI0/XI45/XI1/MM1_g N_VSS_XI0/XI45/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM9 N_XI0/XI45/XI1/NET36_XI0/XI45/XI1/MM9_d
+ N_WL<87>_XI0/XI45/XI1/MM9_g N_BL<14>_XI0/XI45/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM6 N_XI0/XI45/XI1/NET35_XI0/XI45/XI1/MM6_d
+ N_XI0/XI45/XI1/NET36_XI0/XI45/XI1/MM6_g N_VSS_XI0/XI45/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM7 N_XI0/XI45/XI1/NET36_XI0/XI45/XI1/MM7_d
+ N_XI0/XI45/XI1/NET35_XI0/XI45/XI1/MM7_g N_VSS_XI0/XI45/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM8 N_XI0/XI45/XI1/NET35_XI0/XI45/XI1/MM8_d
+ N_WL<87>_XI0/XI45/XI1/MM8_g N_BLN<14>_XI0/XI45/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI1/MM5 N_XI0/XI45/XI1/NET34_XI0/XI45/XI1/MM5_d
+ N_XI0/XI45/XI1/NET33_XI0/XI45/XI1/MM5_g N_VDD_XI0/XI45/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI1/MM4 N_XI0/XI45/XI1/NET33_XI0/XI45/XI1/MM4_d
+ N_XI0/XI45/XI1/NET34_XI0/XI45/XI1/MM4_g N_VDD_XI0/XI45/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI1/MM10 N_XI0/XI45/XI1/NET35_XI0/XI45/XI1/MM10_d
+ N_XI0/XI45/XI1/NET36_XI0/XI45/XI1/MM10_g N_VDD_XI0/XI45/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI1/MM11 N_XI0/XI45/XI1/NET36_XI0/XI45/XI1/MM11_d
+ N_XI0/XI45/XI1/NET35_XI0/XI45/XI1/MM11_g N_VDD_XI0/XI45/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI2/MM2 N_XI0/XI45/XI2/NET34_XI0/XI45/XI2/MM2_d
+ N_XI0/XI45/XI2/NET33_XI0/XI45/XI2/MM2_g N_VSS_XI0/XI45/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM3 N_XI0/XI45/XI2/NET33_XI0/XI45/XI2/MM3_d
+ N_WL<86>_XI0/XI45/XI2/MM3_g N_BLN<13>_XI0/XI45/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM0 N_XI0/XI45/XI2/NET34_XI0/XI45/XI2/MM0_d
+ N_WL<86>_XI0/XI45/XI2/MM0_g N_BL<13>_XI0/XI45/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM1 N_XI0/XI45/XI2/NET33_XI0/XI45/XI2/MM1_d
+ N_XI0/XI45/XI2/NET34_XI0/XI45/XI2/MM1_g N_VSS_XI0/XI45/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM9 N_XI0/XI45/XI2/NET36_XI0/XI45/XI2/MM9_d
+ N_WL<87>_XI0/XI45/XI2/MM9_g N_BL<13>_XI0/XI45/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM6 N_XI0/XI45/XI2/NET35_XI0/XI45/XI2/MM6_d
+ N_XI0/XI45/XI2/NET36_XI0/XI45/XI2/MM6_g N_VSS_XI0/XI45/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM7 N_XI0/XI45/XI2/NET36_XI0/XI45/XI2/MM7_d
+ N_XI0/XI45/XI2/NET35_XI0/XI45/XI2/MM7_g N_VSS_XI0/XI45/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM8 N_XI0/XI45/XI2/NET35_XI0/XI45/XI2/MM8_d
+ N_WL<87>_XI0/XI45/XI2/MM8_g N_BLN<13>_XI0/XI45/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI2/MM5 N_XI0/XI45/XI2/NET34_XI0/XI45/XI2/MM5_d
+ N_XI0/XI45/XI2/NET33_XI0/XI45/XI2/MM5_g N_VDD_XI0/XI45/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI2/MM4 N_XI0/XI45/XI2/NET33_XI0/XI45/XI2/MM4_d
+ N_XI0/XI45/XI2/NET34_XI0/XI45/XI2/MM4_g N_VDD_XI0/XI45/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI2/MM10 N_XI0/XI45/XI2/NET35_XI0/XI45/XI2/MM10_d
+ N_XI0/XI45/XI2/NET36_XI0/XI45/XI2/MM10_g N_VDD_XI0/XI45/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI2/MM11 N_XI0/XI45/XI2/NET36_XI0/XI45/XI2/MM11_d
+ N_XI0/XI45/XI2/NET35_XI0/XI45/XI2/MM11_g N_VDD_XI0/XI45/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI3/MM2 N_XI0/XI45/XI3/NET34_XI0/XI45/XI3/MM2_d
+ N_XI0/XI45/XI3/NET33_XI0/XI45/XI3/MM2_g N_VSS_XI0/XI45/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM3 N_XI0/XI45/XI3/NET33_XI0/XI45/XI3/MM3_d
+ N_WL<86>_XI0/XI45/XI3/MM3_g N_BLN<12>_XI0/XI45/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM0 N_XI0/XI45/XI3/NET34_XI0/XI45/XI3/MM0_d
+ N_WL<86>_XI0/XI45/XI3/MM0_g N_BL<12>_XI0/XI45/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM1 N_XI0/XI45/XI3/NET33_XI0/XI45/XI3/MM1_d
+ N_XI0/XI45/XI3/NET34_XI0/XI45/XI3/MM1_g N_VSS_XI0/XI45/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM9 N_XI0/XI45/XI3/NET36_XI0/XI45/XI3/MM9_d
+ N_WL<87>_XI0/XI45/XI3/MM9_g N_BL<12>_XI0/XI45/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM6 N_XI0/XI45/XI3/NET35_XI0/XI45/XI3/MM6_d
+ N_XI0/XI45/XI3/NET36_XI0/XI45/XI3/MM6_g N_VSS_XI0/XI45/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM7 N_XI0/XI45/XI3/NET36_XI0/XI45/XI3/MM7_d
+ N_XI0/XI45/XI3/NET35_XI0/XI45/XI3/MM7_g N_VSS_XI0/XI45/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM8 N_XI0/XI45/XI3/NET35_XI0/XI45/XI3/MM8_d
+ N_WL<87>_XI0/XI45/XI3/MM8_g N_BLN<12>_XI0/XI45/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI3/MM5 N_XI0/XI45/XI3/NET34_XI0/XI45/XI3/MM5_d
+ N_XI0/XI45/XI3/NET33_XI0/XI45/XI3/MM5_g N_VDD_XI0/XI45/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI3/MM4 N_XI0/XI45/XI3/NET33_XI0/XI45/XI3/MM4_d
+ N_XI0/XI45/XI3/NET34_XI0/XI45/XI3/MM4_g N_VDD_XI0/XI45/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI3/MM10 N_XI0/XI45/XI3/NET35_XI0/XI45/XI3/MM10_d
+ N_XI0/XI45/XI3/NET36_XI0/XI45/XI3/MM10_g N_VDD_XI0/XI45/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI3/MM11 N_XI0/XI45/XI3/NET36_XI0/XI45/XI3/MM11_d
+ N_XI0/XI45/XI3/NET35_XI0/XI45/XI3/MM11_g N_VDD_XI0/XI45/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI4/MM2 N_XI0/XI45/XI4/NET34_XI0/XI45/XI4/MM2_d
+ N_XI0/XI45/XI4/NET33_XI0/XI45/XI4/MM2_g N_VSS_XI0/XI45/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM3 N_XI0/XI45/XI4/NET33_XI0/XI45/XI4/MM3_d
+ N_WL<86>_XI0/XI45/XI4/MM3_g N_BLN<11>_XI0/XI45/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM0 N_XI0/XI45/XI4/NET34_XI0/XI45/XI4/MM0_d
+ N_WL<86>_XI0/XI45/XI4/MM0_g N_BL<11>_XI0/XI45/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM1 N_XI0/XI45/XI4/NET33_XI0/XI45/XI4/MM1_d
+ N_XI0/XI45/XI4/NET34_XI0/XI45/XI4/MM1_g N_VSS_XI0/XI45/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM9 N_XI0/XI45/XI4/NET36_XI0/XI45/XI4/MM9_d
+ N_WL<87>_XI0/XI45/XI4/MM9_g N_BL<11>_XI0/XI45/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM6 N_XI0/XI45/XI4/NET35_XI0/XI45/XI4/MM6_d
+ N_XI0/XI45/XI4/NET36_XI0/XI45/XI4/MM6_g N_VSS_XI0/XI45/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM7 N_XI0/XI45/XI4/NET36_XI0/XI45/XI4/MM7_d
+ N_XI0/XI45/XI4/NET35_XI0/XI45/XI4/MM7_g N_VSS_XI0/XI45/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM8 N_XI0/XI45/XI4/NET35_XI0/XI45/XI4/MM8_d
+ N_WL<87>_XI0/XI45/XI4/MM8_g N_BLN<11>_XI0/XI45/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI4/MM5 N_XI0/XI45/XI4/NET34_XI0/XI45/XI4/MM5_d
+ N_XI0/XI45/XI4/NET33_XI0/XI45/XI4/MM5_g N_VDD_XI0/XI45/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI4/MM4 N_XI0/XI45/XI4/NET33_XI0/XI45/XI4/MM4_d
+ N_XI0/XI45/XI4/NET34_XI0/XI45/XI4/MM4_g N_VDD_XI0/XI45/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI4/MM10 N_XI0/XI45/XI4/NET35_XI0/XI45/XI4/MM10_d
+ N_XI0/XI45/XI4/NET36_XI0/XI45/XI4/MM10_g N_VDD_XI0/XI45/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI4/MM11 N_XI0/XI45/XI4/NET36_XI0/XI45/XI4/MM11_d
+ N_XI0/XI45/XI4/NET35_XI0/XI45/XI4/MM11_g N_VDD_XI0/XI45/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI5/MM2 N_XI0/XI45/XI5/NET34_XI0/XI45/XI5/MM2_d
+ N_XI0/XI45/XI5/NET33_XI0/XI45/XI5/MM2_g N_VSS_XI0/XI45/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM3 N_XI0/XI45/XI5/NET33_XI0/XI45/XI5/MM3_d
+ N_WL<86>_XI0/XI45/XI5/MM3_g N_BLN<10>_XI0/XI45/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM0 N_XI0/XI45/XI5/NET34_XI0/XI45/XI5/MM0_d
+ N_WL<86>_XI0/XI45/XI5/MM0_g N_BL<10>_XI0/XI45/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM1 N_XI0/XI45/XI5/NET33_XI0/XI45/XI5/MM1_d
+ N_XI0/XI45/XI5/NET34_XI0/XI45/XI5/MM1_g N_VSS_XI0/XI45/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM9 N_XI0/XI45/XI5/NET36_XI0/XI45/XI5/MM9_d
+ N_WL<87>_XI0/XI45/XI5/MM9_g N_BL<10>_XI0/XI45/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM6 N_XI0/XI45/XI5/NET35_XI0/XI45/XI5/MM6_d
+ N_XI0/XI45/XI5/NET36_XI0/XI45/XI5/MM6_g N_VSS_XI0/XI45/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM7 N_XI0/XI45/XI5/NET36_XI0/XI45/XI5/MM7_d
+ N_XI0/XI45/XI5/NET35_XI0/XI45/XI5/MM7_g N_VSS_XI0/XI45/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM8 N_XI0/XI45/XI5/NET35_XI0/XI45/XI5/MM8_d
+ N_WL<87>_XI0/XI45/XI5/MM8_g N_BLN<10>_XI0/XI45/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI5/MM5 N_XI0/XI45/XI5/NET34_XI0/XI45/XI5/MM5_d
+ N_XI0/XI45/XI5/NET33_XI0/XI45/XI5/MM5_g N_VDD_XI0/XI45/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI5/MM4 N_XI0/XI45/XI5/NET33_XI0/XI45/XI5/MM4_d
+ N_XI0/XI45/XI5/NET34_XI0/XI45/XI5/MM4_g N_VDD_XI0/XI45/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI5/MM10 N_XI0/XI45/XI5/NET35_XI0/XI45/XI5/MM10_d
+ N_XI0/XI45/XI5/NET36_XI0/XI45/XI5/MM10_g N_VDD_XI0/XI45/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI5/MM11 N_XI0/XI45/XI5/NET36_XI0/XI45/XI5/MM11_d
+ N_XI0/XI45/XI5/NET35_XI0/XI45/XI5/MM11_g N_VDD_XI0/XI45/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI6/MM2 N_XI0/XI45/XI6/NET34_XI0/XI45/XI6/MM2_d
+ N_XI0/XI45/XI6/NET33_XI0/XI45/XI6/MM2_g N_VSS_XI0/XI45/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM3 N_XI0/XI45/XI6/NET33_XI0/XI45/XI6/MM3_d
+ N_WL<86>_XI0/XI45/XI6/MM3_g N_BLN<9>_XI0/XI45/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM0 N_XI0/XI45/XI6/NET34_XI0/XI45/XI6/MM0_d
+ N_WL<86>_XI0/XI45/XI6/MM0_g N_BL<9>_XI0/XI45/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM1 N_XI0/XI45/XI6/NET33_XI0/XI45/XI6/MM1_d
+ N_XI0/XI45/XI6/NET34_XI0/XI45/XI6/MM1_g N_VSS_XI0/XI45/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM9 N_XI0/XI45/XI6/NET36_XI0/XI45/XI6/MM9_d
+ N_WL<87>_XI0/XI45/XI6/MM9_g N_BL<9>_XI0/XI45/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM6 N_XI0/XI45/XI6/NET35_XI0/XI45/XI6/MM6_d
+ N_XI0/XI45/XI6/NET36_XI0/XI45/XI6/MM6_g N_VSS_XI0/XI45/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM7 N_XI0/XI45/XI6/NET36_XI0/XI45/XI6/MM7_d
+ N_XI0/XI45/XI6/NET35_XI0/XI45/XI6/MM7_g N_VSS_XI0/XI45/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM8 N_XI0/XI45/XI6/NET35_XI0/XI45/XI6/MM8_d
+ N_WL<87>_XI0/XI45/XI6/MM8_g N_BLN<9>_XI0/XI45/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI6/MM5 N_XI0/XI45/XI6/NET34_XI0/XI45/XI6/MM5_d
+ N_XI0/XI45/XI6/NET33_XI0/XI45/XI6/MM5_g N_VDD_XI0/XI45/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI6/MM4 N_XI0/XI45/XI6/NET33_XI0/XI45/XI6/MM4_d
+ N_XI0/XI45/XI6/NET34_XI0/XI45/XI6/MM4_g N_VDD_XI0/XI45/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI6/MM10 N_XI0/XI45/XI6/NET35_XI0/XI45/XI6/MM10_d
+ N_XI0/XI45/XI6/NET36_XI0/XI45/XI6/MM10_g N_VDD_XI0/XI45/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI6/MM11 N_XI0/XI45/XI6/NET36_XI0/XI45/XI6/MM11_d
+ N_XI0/XI45/XI6/NET35_XI0/XI45/XI6/MM11_g N_VDD_XI0/XI45/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI7/MM2 N_XI0/XI45/XI7/NET34_XI0/XI45/XI7/MM2_d
+ N_XI0/XI45/XI7/NET33_XI0/XI45/XI7/MM2_g N_VSS_XI0/XI45/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM3 N_XI0/XI45/XI7/NET33_XI0/XI45/XI7/MM3_d
+ N_WL<86>_XI0/XI45/XI7/MM3_g N_BLN<8>_XI0/XI45/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM0 N_XI0/XI45/XI7/NET34_XI0/XI45/XI7/MM0_d
+ N_WL<86>_XI0/XI45/XI7/MM0_g N_BL<8>_XI0/XI45/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM1 N_XI0/XI45/XI7/NET33_XI0/XI45/XI7/MM1_d
+ N_XI0/XI45/XI7/NET34_XI0/XI45/XI7/MM1_g N_VSS_XI0/XI45/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM9 N_XI0/XI45/XI7/NET36_XI0/XI45/XI7/MM9_d
+ N_WL<87>_XI0/XI45/XI7/MM9_g N_BL<8>_XI0/XI45/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM6 N_XI0/XI45/XI7/NET35_XI0/XI45/XI7/MM6_d
+ N_XI0/XI45/XI7/NET36_XI0/XI45/XI7/MM6_g N_VSS_XI0/XI45/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM7 N_XI0/XI45/XI7/NET36_XI0/XI45/XI7/MM7_d
+ N_XI0/XI45/XI7/NET35_XI0/XI45/XI7/MM7_g N_VSS_XI0/XI45/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM8 N_XI0/XI45/XI7/NET35_XI0/XI45/XI7/MM8_d
+ N_WL<87>_XI0/XI45/XI7/MM8_g N_BLN<8>_XI0/XI45/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI7/MM5 N_XI0/XI45/XI7/NET34_XI0/XI45/XI7/MM5_d
+ N_XI0/XI45/XI7/NET33_XI0/XI45/XI7/MM5_g N_VDD_XI0/XI45/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI7/MM4 N_XI0/XI45/XI7/NET33_XI0/XI45/XI7/MM4_d
+ N_XI0/XI45/XI7/NET34_XI0/XI45/XI7/MM4_g N_VDD_XI0/XI45/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI7/MM10 N_XI0/XI45/XI7/NET35_XI0/XI45/XI7/MM10_d
+ N_XI0/XI45/XI7/NET36_XI0/XI45/XI7/MM10_g N_VDD_XI0/XI45/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI7/MM11 N_XI0/XI45/XI7/NET36_XI0/XI45/XI7/MM11_d
+ N_XI0/XI45/XI7/NET35_XI0/XI45/XI7/MM11_g N_VDD_XI0/XI45/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI8/MM2 N_XI0/XI45/XI8/NET34_XI0/XI45/XI8/MM2_d
+ N_XI0/XI45/XI8/NET33_XI0/XI45/XI8/MM2_g N_VSS_XI0/XI45/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM3 N_XI0/XI45/XI8/NET33_XI0/XI45/XI8/MM3_d
+ N_WL<86>_XI0/XI45/XI8/MM3_g N_BLN<7>_XI0/XI45/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM0 N_XI0/XI45/XI8/NET34_XI0/XI45/XI8/MM0_d
+ N_WL<86>_XI0/XI45/XI8/MM0_g N_BL<7>_XI0/XI45/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM1 N_XI0/XI45/XI8/NET33_XI0/XI45/XI8/MM1_d
+ N_XI0/XI45/XI8/NET34_XI0/XI45/XI8/MM1_g N_VSS_XI0/XI45/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM9 N_XI0/XI45/XI8/NET36_XI0/XI45/XI8/MM9_d
+ N_WL<87>_XI0/XI45/XI8/MM9_g N_BL<7>_XI0/XI45/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM6 N_XI0/XI45/XI8/NET35_XI0/XI45/XI8/MM6_d
+ N_XI0/XI45/XI8/NET36_XI0/XI45/XI8/MM6_g N_VSS_XI0/XI45/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM7 N_XI0/XI45/XI8/NET36_XI0/XI45/XI8/MM7_d
+ N_XI0/XI45/XI8/NET35_XI0/XI45/XI8/MM7_g N_VSS_XI0/XI45/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM8 N_XI0/XI45/XI8/NET35_XI0/XI45/XI8/MM8_d
+ N_WL<87>_XI0/XI45/XI8/MM8_g N_BLN<7>_XI0/XI45/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI8/MM5 N_XI0/XI45/XI8/NET34_XI0/XI45/XI8/MM5_d
+ N_XI0/XI45/XI8/NET33_XI0/XI45/XI8/MM5_g N_VDD_XI0/XI45/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI8/MM4 N_XI0/XI45/XI8/NET33_XI0/XI45/XI8/MM4_d
+ N_XI0/XI45/XI8/NET34_XI0/XI45/XI8/MM4_g N_VDD_XI0/XI45/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI8/MM10 N_XI0/XI45/XI8/NET35_XI0/XI45/XI8/MM10_d
+ N_XI0/XI45/XI8/NET36_XI0/XI45/XI8/MM10_g N_VDD_XI0/XI45/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI8/MM11 N_XI0/XI45/XI8/NET36_XI0/XI45/XI8/MM11_d
+ N_XI0/XI45/XI8/NET35_XI0/XI45/XI8/MM11_g N_VDD_XI0/XI45/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI9/MM2 N_XI0/XI45/XI9/NET34_XI0/XI45/XI9/MM2_d
+ N_XI0/XI45/XI9/NET33_XI0/XI45/XI9/MM2_g N_VSS_XI0/XI45/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM3 N_XI0/XI45/XI9/NET33_XI0/XI45/XI9/MM3_d
+ N_WL<86>_XI0/XI45/XI9/MM3_g N_BLN<6>_XI0/XI45/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM0 N_XI0/XI45/XI9/NET34_XI0/XI45/XI9/MM0_d
+ N_WL<86>_XI0/XI45/XI9/MM0_g N_BL<6>_XI0/XI45/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM1 N_XI0/XI45/XI9/NET33_XI0/XI45/XI9/MM1_d
+ N_XI0/XI45/XI9/NET34_XI0/XI45/XI9/MM1_g N_VSS_XI0/XI45/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM9 N_XI0/XI45/XI9/NET36_XI0/XI45/XI9/MM9_d
+ N_WL<87>_XI0/XI45/XI9/MM9_g N_BL<6>_XI0/XI45/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM6 N_XI0/XI45/XI9/NET35_XI0/XI45/XI9/MM6_d
+ N_XI0/XI45/XI9/NET36_XI0/XI45/XI9/MM6_g N_VSS_XI0/XI45/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM7 N_XI0/XI45/XI9/NET36_XI0/XI45/XI9/MM7_d
+ N_XI0/XI45/XI9/NET35_XI0/XI45/XI9/MM7_g N_VSS_XI0/XI45/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM8 N_XI0/XI45/XI9/NET35_XI0/XI45/XI9/MM8_d
+ N_WL<87>_XI0/XI45/XI9/MM8_g N_BLN<6>_XI0/XI45/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI9/MM5 N_XI0/XI45/XI9/NET34_XI0/XI45/XI9/MM5_d
+ N_XI0/XI45/XI9/NET33_XI0/XI45/XI9/MM5_g N_VDD_XI0/XI45/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI9/MM4 N_XI0/XI45/XI9/NET33_XI0/XI45/XI9/MM4_d
+ N_XI0/XI45/XI9/NET34_XI0/XI45/XI9/MM4_g N_VDD_XI0/XI45/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI9/MM10 N_XI0/XI45/XI9/NET35_XI0/XI45/XI9/MM10_d
+ N_XI0/XI45/XI9/NET36_XI0/XI45/XI9/MM10_g N_VDD_XI0/XI45/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI9/MM11 N_XI0/XI45/XI9/NET36_XI0/XI45/XI9/MM11_d
+ N_XI0/XI45/XI9/NET35_XI0/XI45/XI9/MM11_g N_VDD_XI0/XI45/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI10/MM2 N_XI0/XI45/XI10/NET34_XI0/XI45/XI10/MM2_d
+ N_XI0/XI45/XI10/NET33_XI0/XI45/XI10/MM2_g N_VSS_XI0/XI45/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM3 N_XI0/XI45/XI10/NET33_XI0/XI45/XI10/MM3_d
+ N_WL<86>_XI0/XI45/XI10/MM3_g N_BLN<5>_XI0/XI45/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM0 N_XI0/XI45/XI10/NET34_XI0/XI45/XI10/MM0_d
+ N_WL<86>_XI0/XI45/XI10/MM0_g N_BL<5>_XI0/XI45/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM1 N_XI0/XI45/XI10/NET33_XI0/XI45/XI10/MM1_d
+ N_XI0/XI45/XI10/NET34_XI0/XI45/XI10/MM1_g N_VSS_XI0/XI45/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM9 N_XI0/XI45/XI10/NET36_XI0/XI45/XI10/MM9_d
+ N_WL<87>_XI0/XI45/XI10/MM9_g N_BL<5>_XI0/XI45/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM6 N_XI0/XI45/XI10/NET35_XI0/XI45/XI10/MM6_d
+ N_XI0/XI45/XI10/NET36_XI0/XI45/XI10/MM6_g N_VSS_XI0/XI45/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM7 N_XI0/XI45/XI10/NET36_XI0/XI45/XI10/MM7_d
+ N_XI0/XI45/XI10/NET35_XI0/XI45/XI10/MM7_g N_VSS_XI0/XI45/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM8 N_XI0/XI45/XI10/NET35_XI0/XI45/XI10/MM8_d
+ N_WL<87>_XI0/XI45/XI10/MM8_g N_BLN<5>_XI0/XI45/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI10/MM5 N_XI0/XI45/XI10/NET34_XI0/XI45/XI10/MM5_d
+ N_XI0/XI45/XI10/NET33_XI0/XI45/XI10/MM5_g N_VDD_XI0/XI45/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI10/MM4 N_XI0/XI45/XI10/NET33_XI0/XI45/XI10/MM4_d
+ N_XI0/XI45/XI10/NET34_XI0/XI45/XI10/MM4_g N_VDD_XI0/XI45/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI10/MM10 N_XI0/XI45/XI10/NET35_XI0/XI45/XI10/MM10_d
+ N_XI0/XI45/XI10/NET36_XI0/XI45/XI10/MM10_g N_VDD_XI0/XI45/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI10/MM11 N_XI0/XI45/XI10/NET36_XI0/XI45/XI10/MM11_d
+ N_XI0/XI45/XI10/NET35_XI0/XI45/XI10/MM11_g N_VDD_XI0/XI45/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI11/MM2 N_XI0/XI45/XI11/NET34_XI0/XI45/XI11/MM2_d
+ N_XI0/XI45/XI11/NET33_XI0/XI45/XI11/MM2_g N_VSS_XI0/XI45/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM3 N_XI0/XI45/XI11/NET33_XI0/XI45/XI11/MM3_d
+ N_WL<86>_XI0/XI45/XI11/MM3_g N_BLN<4>_XI0/XI45/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM0 N_XI0/XI45/XI11/NET34_XI0/XI45/XI11/MM0_d
+ N_WL<86>_XI0/XI45/XI11/MM0_g N_BL<4>_XI0/XI45/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM1 N_XI0/XI45/XI11/NET33_XI0/XI45/XI11/MM1_d
+ N_XI0/XI45/XI11/NET34_XI0/XI45/XI11/MM1_g N_VSS_XI0/XI45/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM9 N_XI0/XI45/XI11/NET36_XI0/XI45/XI11/MM9_d
+ N_WL<87>_XI0/XI45/XI11/MM9_g N_BL<4>_XI0/XI45/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM6 N_XI0/XI45/XI11/NET35_XI0/XI45/XI11/MM6_d
+ N_XI0/XI45/XI11/NET36_XI0/XI45/XI11/MM6_g N_VSS_XI0/XI45/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM7 N_XI0/XI45/XI11/NET36_XI0/XI45/XI11/MM7_d
+ N_XI0/XI45/XI11/NET35_XI0/XI45/XI11/MM7_g N_VSS_XI0/XI45/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM8 N_XI0/XI45/XI11/NET35_XI0/XI45/XI11/MM8_d
+ N_WL<87>_XI0/XI45/XI11/MM8_g N_BLN<4>_XI0/XI45/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI11/MM5 N_XI0/XI45/XI11/NET34_XI0/XI45/XI11/MM5_d
+ N_XI0/XI45/XI11/NET33_XI0/XI45/XI11/MM5_g N_VDD_XI0/XI45/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI11/MM4 N_XI0/XI45/XI11/NET33_XI0/XI45/XI11/MM4_d
+ N_XI0/XI45/XI11/NET34_XI0/XI45/XI11/MM4_g N_VDD_XI0/XI45/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI11/MM10 N_XI0/XI45/XI11/NET35_XI0/XI45/XI11/MM10_d
+ N_XI0/XI45/XI11/NET36_XI0/XI45/XI11/MM10_g N_VDD_XI0/XI45/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI11/MM11 N_XI0/XI45/XI11/NET36_XI0/XI45/XI11/MM11_d
+ N_XI0/XI45/XI11/NET35_XI0/XI45/XI11/MM11_g N_VDD_XI0/XI45/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI12/MM2 N_XI0/XI45/XI12/NET34_XI0/XI45/XI12/MM2_d
+ N_XI0/XI45/XI12/NET33_XI0/XI45/XI12/MM2_g N_VSS_XI0/XI45/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM3 N_XI0/XI45/XI12/NET33_XI0/XI45/XI12/MM3_d
+ N_WL<86>_XI0/XI45/XI12/MM3_g N_BLN<3>_XI0/XI45/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM0 N_XI0/XI45/XI12/NET34_XI0/XI45/XI12/MM0_d
+ N_WL<86>_XI0/XI45/XI12/MM0_g N_BL<3>_XI0/XI45/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM1 N_XI0/XI45/XI12/NET33_XI0/XI45/XI12/MM1_d
+ N_XI0/XI45/XI12/NET34_XI0/XI45/XI12/MM1_g N_VSS_XI0/XI45/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM9 N_XI0/XI45/XI12/NET36_XI0/XI45/XI12/MM9_d
+ N_WL<87>_XI0/XI45/XI12/MM9_g N_BL<3>_XI0/XI45/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM6 N_XI0/XI45/XI12/NET35_XI0/XI45/XI12/MM6_d
+ N_XI0/XI45/XI12/NET36_XI0/XI45/XI12/MM6_g N_VSS_XI0/XI45/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM7 N_XI0/XI45/XI12/NET36_XI0/XI45/XI12/MM7_d
+ N_XI0/XI45/XI12/NET35_XI0/XI45/XI12/MM7_g N_VSS_XI0/XI45/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM8 N_XI0/XI45/XI12/NET35_XI0/XI45/XI12/MM8_d
+ N_WL<87>_XI0/XI45/XI12/MM8_g N_BLN<3>_XI0/XI45/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI12/MM5 N_XI0/XI45/XI12/NET34_XI0/XI45/XI12/MM5_d
+ N_XI0/XI45/XI12/NET33_XI0/XI45/XI12/MM5_g N_VDD_XI0/XI45/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI12/MM4 N_XI0/XI45/XI12/NET33_XI0/XI45/XI12/MM4_d
+ N_XI0/XI45/XI12/NET34_XI0/XI45/XI12/MM4_g N_VDD_XI0/XI45/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI12/MM10 N_XI0/XI45/XI12/NET35_XI0/XI45/XI12/MM10_d
+ N_XI0/XI45/XI12/NET36_XI0/XI45/XI12/MM10_g N_VDD_XI0/XI45/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI12/MM11 N_XI0/XI45/XI12/NET36_XI0/XI45/XI12/MM11_d
+ N_XI0/XI45/XI12/NET35_XI0/XI45/XI12/MM11_g N_VDD_XI0/XI45/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI13/MM2 N_XI0/XI45/XI13/NET34_XI0/XI45/XI13/MM2_d
+ N_XI0/XI45/XI13/NET33_XI0/XI45/XI13/MM2_g N_VSS_XI0/XI45/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM3 N_XI0/XI45/XI13/NET33_XI0/XI45/XI13/MM3_d
+ N_WL<86>_XI0/XI45/XI13/MM3_g N_BLN<2>_XI0/XI45/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM0 N_XI0/XI45/XI13/NET34_XI0/XI45/XI13/MM0_d
+ N_WL<86>_XI0/XI45/XI13/MM0_g N_BL<2>_XI0/XI45/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM1 N_XI0/XI45/XI13/NET33_XI0/XI45/XI13/MM1_d
+ N_XI0/XI45/XI13/NET34_XI0/XI45/XI13/MM1_g N_VSS_XI0/XI45/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM9 N_XI0/XI45/XI13/NET36_XI0/XI45/XI13/MM9_d
+ N_WL<87>_XI0/XI45/XI13/MM9_g N_BL<2>_XI0/XI45/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM6 N_XI0/XI45/XI13/NET35_XI0/XI45/XI13/MM6_d
+ N_XI0/XI45/XI13/NET36_XI0/XI45/XI13/MM6_g N_VSS_XI0/XI45/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM7 N_XI0/XI45/XI13/NET36_XI0/XI45/XI13/MM7_d
+ N_XI0/XI45/XI13/NET35_XI0/XI45/XI13/MM7_g N_VSS_XI0/XI45/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM8 N_XI0/XI45/XI13/NET35_XI0/XI45/XI13/MM8_d
+ N_WL<87>_XI0/XI45/XI13/MM8_g N_BLN<2>_XI0/XI45/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI13/MM5 N_XI0/XI45/XI13/NET34_XI0/XI45/XI13/MM5_d
+ N_XI0/XI45/XI13/NET33_XI0/XI45/XI13/MM5_g N_VDD_XI0/XI45/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI13/MM4 N_XI0/XI45/XI13/NET33_XI0/XI45/XI13/MM4_d
+ N_XI0/XI45/XI13/NET34_XI0/XI45/XI13/MM4_g N_VDD_XI0/XI45/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI13/MM10 N_XI0/XI45/XI13/NET35_XI0/XI45/XI13/MM10_d
+ N_XI0/XI45/XI13/NET36_XI0/XI45/XI13/MM10_g N_VDD_XI0/XI45/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI13/MM11 N_XI0/XI45/XI13/NET36_XI0/XI45/XI13/MM11_d
+ N_XI0/XI45/XI13/NET35_XI0/XI45/XI13/MM11_g N_VDD_XI0/XI45/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI14/MM2 N_XI0/XI45/XI14/NET34_XI0/XI45/XI14/MM2_d
+ N_XI0/XI45/XI14/NET33_XI0/XI45/XI14/MM2_g N_VSS_XI0/XI45/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM3 N_XI0/XI45/XI14/NET33_XI0/XI45/XI14/MM3_d
+ N_WL<86>_XI0/XI45/XI14/MM3_g N_BLN<1>_XI0/XI45/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM0 N_XI0/XI45/XI14/NET34_XI0/XI45/XI14/MM0_d
+ N_WL<86>_XI0/XI45/XI14/MM0_g N_BL<1>_XI0/XI45/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM1 N_XI0/XI45/XI14/NET33_XI0/XI45/XI14/MM1_d
+ N_XI0/XI45/XI14/NET34_XI0/XI45/XI14/MM1_g N_VSS_XI0/XI45/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM9 N_XI0/XI45/XI14/NET36_XI0/XI45/XI14/MM9_d
+ N_WL<87>_XI0/XI45/XI14/MM9_g N_BL<1>_XI0/XI45/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM6 N_XI0/XI45/XI14/NET35_XI0/XI45/XI14/MM6_d
+ N_XI0/XI45/XI14/NET36_XI0/XI45/XI14/MM6_g N_VSS_XI0/XI45/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM7 N_XI0/XI45/XI14/NET36_XI0/XI45/XI14/MM7_d
+ N_XI0/XI45/XI14/NET35_XI0/XI45/XI14/MM7_g N_VSS_XI0/XI45/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM8 N_XI0/XI45/XI14/NET35_XI0/XI45/XI14/MM8_d
+ N_WL<87>_XI0/XI45/XI14/MM8_g N_BLN<1>_XI0/XI45/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI14/MM5 N_XI0/XI45/XI14/NET34_XI0/XI45/XI14/MM5_d
+ N_XI0/XI45/XI14/NET33_XI0/XI45/XI14/MM5_g N_VDD_XI0/XI45/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI14/MM4 N_XI0/XI45/XI14/NET33_XI0/XI45/XI14/MM4_d
+ N_XI0/XI45/XI14/NET34_XI0/XI45/XI14/MM4_g N_VDD_XI0/XI45/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI14/MM10 N_XI0/XI45/XI14/NET35_XI0/XI45/XI14/MM10_d
+ N_XI0/XI45/XI14/NET36_XI0/XI45/XI14/MM10_g N_VDD_XI0/XI45/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI14/MM11 N_XI0/XI45/XI14/NET36_XI0/XI45/XI14/MM11_d
+ N_XI0/XI45/XI14/NET35_XI0/XI45/XI14/MM11_g N_VDD_XI0/XI45/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI15/MM2 N_XI0/XI45/XI15/NET34_XI0/XI45/XI15/MM2_d
+ N_XI0/XI45/XI15/NET33_XI0/XI45/XI15/MM2_g N_VSS_XI0/XI45/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM3 N_XI0/XI45/XI15/NET33_XI0/XI45/XI15/MM3_d
+ N_WL<86>_XI0/XI45/XI15/MM3_g N_BLN<0>_XI0/XI45/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM0 N_XI0/XI45/XI15/NET34_XI0/XI45/XI15/MM0_d
+ N_WL<86>_XI0/XI45/XI15/MM0_g N_BL<0>_XI0/XI45/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM1 N_XI0/XI45/XI15/NET33_XI0/XI45/XI15/MM1_d
+ N_XI0/XI45/XI15/NET34_XI0/XI45/XI15/MM1_g N_VSS_XI0/XI45/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM9 N_XI0/XI45/XI15/NET36_XI0/XI45/XI15/MM9_d
+ N_WL<87>_XI0/XI45/XI15/MM9_g N_BL<0>_XI0/XI45/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM6 N_XI0/XI45/XI15/NET35_XI0/XI45/XI15/MM6_d
+ N_XI0/XI45/XI15/NET36_XI0/XI45/XI15/MM6_g N_VSS_XI0/XI45/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM7 N_XI0/XI45/XI15/NET36_XI0/XI45/XI15/MM7_d
+ N_XI0/XI45/XI15/NET35_XI0/XI45/XI15/MM7_g N_VSS_XI0/XI45/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM8 N_XI0/XI45/XI15/NET35_XI0/XI45/XI15/MM8_d
+ N_WL<87>_XI0/XI45/XI15/MM8_g N_BLN<0>_XI0/XI45/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI45/XI15/MM5 N_XI0/XI45/XI15/NET34_XI0/XI45/XI15/MM5_d
+ N_XI0/XI45/XI15/NET33_XI0/XI45/XI15/MM5_g N_VDD_XI0/XI45/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI15/MM4 N_XI0/XI45/XI15/NET33_XI0/XI45/XI15/MM4_d
+ N_XI0/XI45/XI15/NET34_XI0/XI45/XI15/MM4_g N_VDD_XI0/XI45/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI15/MM10 N_XI0/XI45/XI15/NET35_XI0/XI45/XI15/MM10_d
+ N_XI0/XI45/XI15/NET36_XI0/XI45/XI15/MM10_g N_VDD_XI0/XI45/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI45/XI15/MM11 N_XI0/XI45/XI15/NET36_XI0/XI45/XI15/MM11_d
+ N_XI0/XI45/XI15/NET35_XI0/XI45/XI15/MM11_g N_VDD_XI0/XI45/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI0/MM2 N_XI0/XI46/XI0/NET34_XI0/XI46/XI0/MM2_d
+ N_XI0/XI46/XI0/NET33_XI0/XI46/XI0/MM2_g N_VSS_XI0/XI46/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM3 N_XI0/XI46/XI0/NET33_XI0/XI46/XI0/MM3_d
+ N_WL<88>_XI0/XI46/XI0/MM3_g N_BLN<15>_XI0/XI46/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM0 N_XI0/XI46/XI0/NET34_XI0/XI46/XI0/MM0_d
+ N_WL<88>_XI0/XI46/XI0/MM0_g N_BL<15>_XI0/XI46/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM1 N_XI0/XI46/XI0/NET33_XI0/XI46/XI0/MM1_d
+ N_XI0/XI46/XI0/NET34_XI0/XI46/XI0/MM1_g N_VSS_XI0/XI46/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM9 N_XI0/XI46/XI0/NET36_XI0/XI46/XI0/MM9_d
+ N_WL<89>_XI0/XI46/XI0/MM9_g N_BL<15>_XI0/XI46/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM6 N_XI0/XI46/XI0/NET35_XI0/XI46/XI0/MM6_d
+ N_XI0/XI46/XI0/NET36_XI0/XI46/XI0/MM6_g N_VSS_XI0/XI46/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM7 N_XI0/XI46/XI0/NET36_XI0/XI46/XI0/MM7_d
+ N_XI0/XI46/XI0/NET35_XI0/XI46/XI0/MM7_g N_VSS_XI0/XI46/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM8 N_XI0/XI46/XI0/NET35_XI0/XI46/XI0/MM8_d
+ N_WL<89>_XI0/XI46/XI0/MM8_g N_BLN<15>_XI0/XI46/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI0/MM5 N_XI0/XI46/XI0/NET34_XI0/XI46/XI0/MM5_d
+ N_XI0/XI46/XI0/NET33_XI0/XI46/XI0/MM5_g N_VDD_XI0/XI46/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI0/MM4 N_XI0/XI46/XI0/NET33_XI0/XI46/XI0/MM4_d
+ N_XI0/XI46/XI0/NET34_XI0/XI46/XI0/MM4_g N_VDD_XI0/XI46/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI0/MM10 N_XI0/XI46/XI0/NET35_XI0/XI46/XI0/MM10_d
+ N_XI0/XI46/XI0/NET36_XI0/XI46/XI0/MM10_g N_VDD_XI0/XI46/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI0/MM11 N_XI0/XI46/XI0/NET36_XI0/XI46/XI0/MM11_d
+ N_XI0/XI46/XI0/NET35_XI0/XI46/XI0/MM11_g N_VDD_XI0/XI46/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI1/MM2 N_XI0/XI46/XI1/NET34_XI0/XI46/XI1/MM2_d
+ N_XI0/XI46/XI1/NET33_XI0/XI46/XI1/MM2_g N_VSS_XI0/XI46/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM3 N_XI0/XI46/XI1/NET33_XI0/XI46/XI1/MM3_d
+ N_WL<88>_XI0/XI46/XI1/MM3_g N_BLN<14>_XI0/XI46/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM0 N_XI0/XI46/XI1/NET34_XI0/XI46/XI1/MM0_d
+ N_WL<88>_XI0/XI46/XI1/MM0_g N_BL<14>_XI0/XI46/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM1 N_XI0/XI46/XI1/NET33_XI0/XI46/XI1/MM1_d
+ N_XI0/XI46/XI1/NET34_XI0/XI46/XI1/MM1_g N_VSS_XI0/XI46/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM9 N_XI0/XI46/XI1/NET36_XI0/XI46/XI1/MM9_d
+ N_WL<89>_XI0/XI46/XI1/MM9_g N_BL<14>_XI0/XI46/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM6 N_XI0/XI46/XI1/NET35_XI0/XI46/XI1/MM6_d
+ N_XI0/XI46/XI1/NET36_XI0/XI46/XI1/MM6_g N_VSS_XI0/XI46/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM7 N_XI0/XI46/XI1/NET36_XI0/XI46/XI1/MM7_d
+ N_XI0/XI46/XI1/NET35_XI0/XI46/XI1/MM7_g N_VSS_XI0/XI46/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM8 N_XI0/XI46/XI1/NET35_XI0/XI46/XI1/MM8_d
+ N_WL<89>_XI0/XI46/XI1/MM8_g N_BLN<14>_XI0/XI46/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI1/MM5 N_XI0/XI46/XI1/NET34_XI0/XI46/XI1/MM5_d
+ N_XI0/XI46/XI1/NET33_XI0/XI46/XI1/MM5_g N_VDD_XI0/XI46/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI1/MM4 N_XI0/XI46/XI1/NET33_XI0/XI46/XI1/MM4_d
+ N_XI0/XI46/XI1/NET34_XI0/XI46/XI1/MM4_g N_VDD_XI0/XI46/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI1/MM10 N_XI0/XI46/XI1/NET35_XI0/XI46/XI1/MM10_d
+ N_XI0/XI46/XI1/NET36_XI0/XI46/XI1/MM10_g N_VDD_XI0/XI46/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI1/MM11 N_XI0/XI46/XI1/NET36_XI0/XI46/XI1/MM11_d
+ N_XI0/XI46/XI1/NET35_XI0/XI46/XI1/MM11_g N_VDD_XI0/XI46/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI2/MM2 N_XI0/XI46/XI2/NET34_XI0/XI46/XI2/MM2_d
+ N_XI0/XI46/XI2/NET33_XI0/XI46/XI2/MM2_g N_VSS_XI0/XI46/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM3 N_XI0/XI46/XI2/NET33_XI0/XI46/XI2/MM3_d
+ N_WL<88>_XI0/XI46/XI2/MM3_g N_BLN<13>_XI0/XI46/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM0 N_XI0/XI46/XI2/NET34_XI0/XI46/XI2/MM0_d
+ N_WL<88>_XI0/XI46/XI2/MM0_g N_BL<13>_XI0/XI46/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM1 N_XI0/XI46/XI2/NET33_XI0/XI46/XI2/MM1_d
+ N_XI0/XI46/XI2/NET34_XI0/XI46/XI2/MM1_g N_VSS_XI0/XI46/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM9 N_XI0/XI46/XI2/NET36_XI0/XI46/XI2/MM9_d
+ N_WL<89>_XI0/XI46/XI2/MM9_g N_BL<13>_XI0/XI46/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM6 N_XI0/XI46/XI2/NET35_XI0/XI46/XI2/MM6_d
+ N_XI0/XI46/XI2/NET36_XI0/XI46/XI2/MM6_g N_VSS_XI0/XI46/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM7 N_XI0/XI46/XI2/NET36_XI0/XI46/XI2/MM7_d
+ N_XI0/XI46/XI2/NET35_XI0/XI46/XI2/MM7_g N_VSS_XI0/XI46/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM8 N_XI0/XI46/XI2/NET35_XI0/XI46/XI2/MM8_d
+ N_WL<89>_XI0/XI46/XI2/MM8_g N_BLN<13>_XI0/XI46/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI2/MM5 N_XI0/XI46/XI2/NET34_XI0/XI46/XI2/MM5_d
+ N_XI0/XI46/XI2/NET33_XI0/XI46/XI2/MM5_g N_VDD_XI0/XI46/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI2/MM4 N_XI0/XI46/XI2/NET33_XI0/XI46/XI2/MM4_d
+ N_XI0/XI46/XI2/NET34_XI0/XI46/XI2/MM4_g N_VDD_XI0/XI46/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI2/MM10 N_XI0/XI46/XI2/NET35_XI0/XI46/XI2/MM10_d
+ N_XI0/XI46/XI2/NET36_XI0/XI46/XI2/MM10_g N_VDD_XI0/XI46/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI2/MM11 N_XI0/XI46/XI2/NET36_XI0/XI46/XI2/MM11_d
+ N_XI0/XI46/XI2/NET35_XI0/XI46/XI2/MM11_g N_VDD_XI0/XI46/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI3/MM2 N_XI0/XI46/XI3/NET34_XI0/XI46/XI3/MM2_d
+ N_XI0/XI46/XI3/NET33_XI0/XI46/XI3/MM2_g N_VSS_XI0/XI46/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM3 N_XI0/XI46/XI3/NET33_XI0/XI46/XI3/MM3_d
+ N_WL<88>_XI0/XI46/XI3/MM3_g N_BLN<12>_XI0/XI46/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM0 N_XI0/XI46/XI3/NET34_XI0/XI46/XI3/MM0_d
+ N_WL<88>_XI0/XI46/XI3/MM0_g N_BL<12>_XI0/XI46/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM1 N_XI0/XI46/XI3/NET33_XI0/XI46/XI3/MM1_d
+ N_XI0/XI46/XI3/NET34_XI0/XI46/XI3/MM1_g N_VSS_XI0/XI46/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM9 N_XI0/XI46/XI3/NET36_XI0/XI46/XI3/MM9_d
+ N_WL<89>_XI0/XI46/XI3/MM9_g N_BL<12>_XI0/XI46/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM6 N_XI0/XI46/XI3/NET35_XI0/XI46/XI3/MM6_d
+ N_XI0/XI46/XI3/NET36_XI0/XI46/XI3/MM6_g N_VSS_XI0/XI46/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM7 N_XI0/XI46/XI3/NET36_XI0/XI46/XI3/MM7_d
+ N_XI0/XI46/XI3/NET35_XI0/XI46/XI3/MM7_g N_VSS_XI0/XI46/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM8 N_XI0/XI46/XI3/NET35_XI0/XI46/XI3/MM8_d
+ N_WL<89>_XI0/XI46/XI3/MM8_g N_BLN<12>_XI0/XI46/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI3/MM5 N_XI0/XI46/XI3/NET34_XI0/XI46/XI3/MM5_d
+ N_XI0/XI46/XI3/NET33_XI0/XI46/XI3/MM5_g N_VDD_XI0/XI46/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI3/MM4 N_XI0/XI46/XI3/NET33_XI0/XI46/XI3/MM4_d
+ N_XI0/XI46/XI3/NET34_XI0/XI46/XI3/MM4_g N_VDD_XI0/XI46/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI3/MM10 N_XI0/XI46/XI3/NET35_XI0/XI46/XI3/MM10_d
+ N_XI0/XI46/XI3/NET36_XI0/XI46/XI3/MM10_g N_VDD_XI0/XI46/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI3/MM11 N_XI0/XI46/XI3/NET36_XI0/XI46/XI3/MM11_d
+ N_XI0/XI46/XI3/NET35_XI0/XI46/XI3/MM11_g N_VDD_XI0/XI46/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI4/MM2 N_XI0/XI46/XI4/NET34_XI0/XI46/XI4/MM2_d
+ N_XI0/XI46/XI4/NET33_XI0/XI46/XI4/MM2_g N_VSS_XI0/XI46/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM3 N_XI0/XI46/XI4/NET33_XI0/XI46/XI4/MM3_d
+ N_WL<88>_XI0/XI46/XI4/MM3_g N_BLN<11>_XI0/XI46/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM0 N_XI0/XI46/XI4/NET34_XI0/XI46/XI4/MM0_d
+ N_WL<88>_XI0/XI46/XI4/MM0_g N_BL<11>_XI0/XI46/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM1 N_XI0/XI46/XI4/NET33_XI0/XI46/XI4/MM1_d
+ N_XI0/XI46/XI4/NET34_XI0/XI46/XI4/MM1_g N_VSS_XI0/XI46/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM9 N_XI0/XI46/XI4/NET36_XI0/XI46/XI4/MM9_d
+ N_WL<89>_XI0/XI46/XI4/MM9_g N_BL<11>_XI0/XI46/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM6 N_XI0/XI46/XI4/NET35_XI0/XI46/XI4/MM6_d
+ N_XI0/XI46/XI4/NET36_XI0/XI46/XI4/MM6_g N_VSS_XI0/XI46/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM7 N_XI0/XI46/XI4/NET36_XI0/XI46/XI4/MM7_d
+ N_XI0/XI46/XI4/NET35_XI0/XI46/XI4/MM7_g N_VSS_XI0/XI46/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM8 N_XI0/XI46/XI4/NET35_XI0/XI46/XI4/MM8_d
+ N_WL<89>_XI0/XI46/XI4/MM8_g N_BLN<11>_XI0/XI46/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI4/MM5 N_XI0/XI46/XI4/NET34_XI0/XI46/XI4/MM5_d
+ N_XI0/XI46/XI4/NET33_XI0/XI46/XI4/MM5_g N_VDD_XI0/XI46/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI4/MM4 N_XI0/XI46/XI4/NET33_XI0/XI46/XI4/MM4_d
+ N_XI0/XI46/XI4/NET34_XI0/XI46/XI4/MM4_g N_VDD_XI0/XI46/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI4/MM10 N_XI0/XI46/XI4/NET35_XI0/XI46/XI4/MM10_d
+ N_XI0/XI46/XI4/NET36_XI0/XI46/XI4/MM10_g N_VDD_XI0/XI46/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI4/MM11 N_XI0/XI46/XI4/NET36_XI0/XI46/XI4/MM11_d
+ N_XI0/XI46/XI4/NET35_XI0/XI46/XI4/MM11_g N_VDD_XI0/XI46/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI5/MM2 N_XI0/XI46/XI5/NET34_XI0/XI46/XI5/MM2_d
+ N_XI0/XI46/XI5/NET33_XI0/XI46/XI5/MM2_g N_VSS_XI0/XI46/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM3 N_XI0/XI46/XI5/NET33_XI0/XI46/XI5/MM3_d
+ N_WL<88>_XI0/XI46/XI5/MM3_g N_BLN<10>_XI0/XI46/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM0 N_XI0/XI46/XI5/NET34_XI0/XI46/XI5/MM0_d
+ N_WL<88>_XI0/XI46/XI5/MM0_g N_BL<10>_XI0/XI46/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM1 N_XI0/XI46/XI5/NET33_XI0/XI46/XI5/MM1_d
+ N_XI0/XI46/XI5/NET34_XI0/XI46/XI5/MM1_g N_VSS_XI0/XI46/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM9 N_XI0/XI46/XI5/NET36_XI0/XI46/XI5/MM9_d
+ N_WL<89>_XI0/XI46/XI5/MM9_g N_BL<10>_XI0/XI46/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM6 N_XI0/XI46/XI5/NET35_XI0/XI46/XI5/MM6_d
+ N_XI0/XI46/XI5/NET36_XI0/XI46/XI5/MM6_g N_VSS_XI0/XI46/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM7 N_XI0/XI46/XI5/NET36_XI0/XI46/XI5/MM7_d
+ N_XI0/XI46/XI5/NET35_XI0/XI46/XI5/MM7_g N_VSS_XI0/XI46/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM8 N_XI0/XI46/XI5/NET35_XI0/XI46/XI5/MM8_d
+ N_WL<89>_XI0/XI46/XI5/MM8_g N_BLN<10>_XI0/XI46/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI5/MM5 N_XI0/XI46/XI5/NET34_XI0/XI46/XI5/MM5_d
+ N_XI0/XI46/XI5/NET33_XI0/XI46/XI5/MM5_g N_VDD_XI0/XI46/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI5/MM4 N_XI0/XI46/XI5/NET33_XI0/XI46/XI5/MM4_d
+ N_XI0/XI46/XI5/NET34_XI0/XI46/XI5/MM4_g N_VDD_XI0/XI46/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI5/MM10 N_XI0/XI46/XI5/NET35_XI0/XI46/XI5/MM10_d
+ N_XI0/XI46/XI5/NET36_XI0/XI46/XI5/MM10_g N_VDD_XI0/XI46/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI5/MM11 N_XI0/XI46/XI5/NET36_XI0/XI46/XI5/MM11_d
+ N_XI0/XI46/XI5/NET35_XI0/XI46/XI5/MM11_g N_VDD_XI0/XI46/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI6/MM2 N_XI0/XI46/XI6/NET34_XI0/XI46/XI6/MM2_d
+ N_XI0/XI46/XI6/NET33_XI0/XI46/XI6/MM2_g N_VSS_XI0/XI46/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM3 N_XI0/XI46/XI6/NET33_XI0/XI46/XI6/MM3_d
+ N_WL<88>_XI0/XI46/XI6/MM3_g N_BLN<9>_XI0/XI46/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM0 N_XI0/XI46/XI6/NET34_XI0/XI46/XI6/MM0_d
+ N_WL<88>_XI0/XI46/XI6/MM0_g N_BL<9>_XI0/XI46/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM1 N_XI0/XI46/XI6/NET33_XI0/XI46/XI6/MM1_d
+ N_XI0/XI46/XI6/NET34_XI0/XI46/XI6/MM1_g N_VSS_XI0/XI46/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM9 N_XI0/XI46/XI6/NET36_XI0/XI46/XI6/MM9_d
+ N_WL<89>_XI0/XI46/XI6/MM9_g N_BL<9>_XI0/XI46/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM6 N_XI0/XI46/XI6/NET35_XI0/XI46/XI6/MM6_d
+ N_XI0/XI46/XI6/NET36_XI0/XI46/XI6/MM6_g N_VSS_XI0/XI46/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM7 N_XI0/XI46/XI6/NET36_XI0/XI46/XI6/MM7_d
+ N_XI0/XI46/XI6/NET35_XI0/XI46/XI6/MM7_g N_VSS_XI0/XI46/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM8 N_XI0/XI46/XI6/NET35_XI0/XI46/XI6/MM8_d
+ N_WL<89>_XI0/XI46/XI6/MM8_g N_BLN<9>_XI0/XI46/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI6/MM5 N_XI0/XI46/XI6/NET34_XI0/XI46/XI6/MM5_d
+ N_XI0/XI46/XI6/NET33_XI0/XI46/XI6/MM5_g N_VDD_XI0/XI46/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI6/MM4 N_XI0/XI46/XI6/NET33_XI0/XI46/XI6/MM4_d
+ N_XI0/XI46/XI6/NET34_XI0/XI46/XI6/MM4_g N_VDD_XI0/XI46/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI6/MM10 N_XI0/XI46/XI6/NET35_XI0/XI46/XI6/MM10_d
+ N_XI0/XI46/XI6/NET36_XI0/XI46/XI6/MM10_g N_VDD_XI0/XI46/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI6/MM11 N_XI0/XI46/XI6/NET36_XI0/XI46/XI6/MM11_d
+ N_XI0/XI46/XI6/NET35_XI0/XI46/XI6/MM11_g N_VDD_XI0/XI46/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI7/MM2 N_XI0/XI46/XI7/NET34_XI0/XI46/XI7/MM2_d
+ N_XI0/XI46/XI7/NET33_XI0/XI46/XI7/MM2_g N_VSS_XI0/XI46/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM3 N_XI0/XI46/XI7/NET33_XI0/XI46/XI7/MM3_d
+ N_WL<88>_XI0/XI46/XI7/MM3_g N_BLN<8>_XI0/XI46/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM0 N_XI0/XI46/XI7/NET34_XI0/XI46/XI7/MM0_d
+ N_WL<88>_XI0/XI46/XI7/MM0_g N_BL<8>_XI0/XI46/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM1 N_XI0/XI46/XI7/NET33_XI0/XI46/XI7/MM1_d
+ N_XI0/XI46/XI7/NET34_XI0/XI46/XI7/MM1_g N_VSS_XI0/XI46/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM9 N_XI0/XI46/XI7/NET36_XI0/XI46/XI7/MM9_d
+ N_WL<89>_XI0/XI46/XI7/MM9_g N_BL<8>_XI0/XI46/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM6 N_XI0/XI46/XI7/NET35_XI0/XI46/XI7/MM6_d
+ N_XI0/XI46/XI7/NET36_XI0/XI46/XI7/MM6_g N_VSS_XI0/XI46/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM7 N_XI0/XI46/XI7/NET36_XI0/XI46/XI7/MM7_d
+ N_XI0/XI46/XI7/NET35_XI0/XI46/XI7/MM7_g N_VSS_XI0/XI46/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM8 N_XI0/XI46/XI7/NET35_XI0/XI46/XI7/MM8_d
+ N_WL<89>_XI0/XI46/XI7/MM8_g N_BLN<8>_XI0/XI46/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI7/MM5 N_XI0/XI46/XI7/NET34_XI0/XI46/XI7/MM5_d
+ N_XI0/XI46/XI7/NET33_XI0/XI46/XI7/MM5_g N_VDD_XI0/XI46/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI7/MM4 N_XI0/XI46/XI7/NET33_XI0/XI46/XI7/MM4_d
+ N_XI0/XI46/XI7/NET34_XI0/XI46/XI7/MM4_g N_VDD_XI0/XI46/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI7/MM10 N_XI0/XI46/XI7/NET35_XI0/XI46/XI7/MM10_d
+ N_XI0/XI46/XI7/NET36_XI0/XI46/XI7/MM10_g N_VDD_XI0/XI46/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI7/MM11 N_XI0/XI46/XI7/NET36_XI0/XI46/XI7/MM11_d
+ N_XI0/XI46/XI7/NET35_XI0/XI46/XI7/MM11_g N_VDD_XI0/XI46/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI8/MM2 N_XI0/XI46/XI8/NET34_XI0/XI46/XI8/MM2_d
+ N_XI0/XI46/XI8/NET33_XI0/XI46/XI8/MM2_g N_VSS_XI0/XI46/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM3 N_XI0/XI46/XI8/NET33_XI0/XI46/XI8/MM3_d
+ N_WL<88>_XI0/XI46/XI8/MM3_g N_BLN<7>_XI0/XI46/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM0 N_XI0/XI46/XI8/NET34_XI0/XI46/XI8/MM0_d
+ N_WL<88>_XI0/XI46/XI8/MM0_g N_BL<7>_XI0/XI46/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM1 N_XI0/XI46/XI8/NET33_XI0/XI46/XI8/MM1_d
+ N_XI0/XI46/XI8/NET34_XI0/XI46/XI8/MM1_g N_VSS_XI0/XI46/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM9 N_XI0/XI46/XI8/NET36_XI0/XI46/XI8/MM9_d
+ N_WL<89>_XI0/XI46/XI8/MM9_g N_BL<7>_XI0/XI46/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM6 N_XI0/XI46/XI8/NET35_XI0/XI46/XI8/MM6_d
+ N_XI0/XI46/XI8/NET36_XI0/XI46/XI8/MM6_g N_VSS_XI0/XI46/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM7 N_XI0/XI46/XI8/NET36_XI0/XI46/XI8/MM7_d
+ N_XI0/XI46/XI8/NET35_XI0/XI46/XI8/MM7_g N_VSS_XI0/XI46/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM8 N_XI0/XI46/XI8/NET35_XI0/XI46/XI8/MM8_d
+ N_WL<89>_XI0/XI46/XI8/MM8_g N_BLN<7>_XI0/XI46/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI8/MM5 N_XI0/XI46/XI8/NET34_XI0/XI46/XI8/MM5_d
+ N_XI0/XI46/XI8/NET33_XI0/XI46/XI8/MM5_g N_VDD_XI0/XI46/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI8/MM4 N_XI0/XI46/XI8/NET33_XI0/XI46/XI8/MM4_d
+ N_XI0/XI46/XI8/NET34_XI0/XI46/XI8/MM4_g N_VDD_XI0/XI46/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI8/MM10 N_XI0/XI46/XI8/NET35_XI0/XI46/XI8/MM10_d
+ N_XI0/XI46/XI8/NET36_XI0/XI46/XI8/MM10_g N_VDD_XI0/XI46/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI8/MM11 N_XI0/XI46/XI8/NET36_XI0/XI46/XI8/MM11_d
+ N_XI0/XI46/XI8/NET35_XI0/XI46/XI8/MM11_g N_VDD_XI0/XI46/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI9/MM2 N_XI0/XI46/XI9/NET34_XI0/XI46/XI9/MM2_d
+ N_XI0/XI46/XI9/NET33_XI0/XI46/XI9/MM2_g N_VSS_XI0/XI46/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM3 N_XI0/XI46/XI9/NET33_XI0/XI46/XI9/MM3_d
+ N_WL<88>_XI0/XI46/XI9/MM3_g N_BLN<6>_XI0/XI46/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM0 N_XI0/XI46/XI9/NET34_XI0/XI46/XI9/MM0_d
+ N_WL<88>_XI0/XI46/XI9/MM0_g N_BL<6>_XI0/XI46/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM1 N_XI0/XI46/XI9/NET33_XI0/XI46/XI9/MM1_d
+ N_XI0/XI46/XI9/NET34_XI0/XI46/XI9/MM1_g N_VSS_XI0/XI46/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM9 N_XI0/XI46/XI9/NET36_XI0/XI46/XI9/MM9_d
+ N_WL<89>_XI0/XI46/XI9/MM9_g N_BL<6>_XI0/XI46/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM6 N_XI0/XI46/XI9/NET35_XI0/XI46/XI9/MM6_d
+ N_XI0/XI46/XI9/NET36_XI0/XI46/XI9/MM6_g N_VSS_XI0/XI46/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM7 N_XI0/XI46/XI9/NET36_XI0/XI46/XI9/MM7_d
+ N_XI0/XI46/XI9/NET35_XI0/XI46/XI9/MM7_g N_VSS_XI0/XI46/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM8 N_XI0/XI46/XI9/NET35_XI0/XI46/XI9/MM8_d
+ N_WL<89>_XI0/XI46/XI9/MM8_g N_BLN<6>_XI0/XI46/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI9/MM5 N_XI0/XI46/XI9/NET34_XI0/XI46/XI9/MM5_d
+ N_XI0/XI46/XI9/NET33_XI0/XI46/XI9/MM5_g N_VDD_XI0/XI46/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI9/MM4 N_XI0/XI46/XI9/NET33_XI0/XI46/XI9/MM4_d
+ N_XI0/XI46/XI9/NET34_XI0/XI46/XI9/MM4_g N_VDD_XI0/XI46/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI9/MM10 N_XI0/XI46/XI9/NET35_XI0/XI46/XI9/MM10_d
+ N_XI0/XI46/XI9/NET36_XI0/XI46/XI9/MM10_g N_VDD_XI0/XI46/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI9/MM11 N_XI0/XI46/XI9/NET36_XI0/XI46/XI9/MM11_d
+ N_XI0/XI46/XI9/NET35_XI0/XI46/XI9/MM11_g N_VDD_XI0/XI46/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI10/MM2 N_XI0/XI46/XI10/NET34_XI0/XI46/XI10/MM2_d
+ N_XI0/XI46/XI10/NET33_XI0/XI46/XI10/MM2_g N_VSS_XI0/XI46/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM3 N_XI0/XI46/XI10/NET33_XI0/XI46/XI10/MM3_d
+ N_WL<88>_XI0/XI46/XI10/MM3_g N_BLN<5>_XI0/XI46/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM0 N_XI0/XI46/XI10/NET34_XI0/XI46/XI10/MM0_d
+ N_WL<88>_XI0/XI46/XI10/MM0_g N_BL<5>_XI0/XI46/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM1 N_XI0/XI46/XI10/NET33_XI0/XI46/XI10/MM1_d
+ N_XI0/XI46/XI10/NET34_XI0/XI46/XI10/MM1_g N_VSS_XI0/XI46/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM9 N_XI0/XI46/XI10/NET36_XI0/XI46/XI10/MM9_d
+ N_WL<89>_XI0/XI46/XI10/MM9_g N_BL<5>_XI0/XI46/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM6 N_XI0/XI46/XI10/NET35_XI0/XI46/XI10/MM6_d
+ N_XI0/XI46/XI10/NET36_XI0/XI46/XI10/MM6_g N_VSS_XI0/XI46/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM7 N_XI0/XI46/XI10/NET36_XI0/XI46/XI10/MM7_d
+ N_XI0/XI46/XI10/NET35_XI0/XI46/XI10/MM7_g N_VSS_XI0/XI46/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM8 N_XI0/XI46/XI10/NET35_XI0/XI46/XI10/MM8_d
+ N_WL<89>_XI0/XI46/XI10/MM8_g N_BLN<5>_XI0/XI46/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI10/MM5 N_XI0/XI46/XI10/NET34_XI0/XI46/XI10/MM5_d
+ N_XI0/XI46/XI10/NET33_XI0/XI46/XI10/MM5_g N_VDD_XI0/XI46/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI10/MM4 N_XI0/XI46/XI10/NET33_XI0/XI46/XI10/MM4_d
+ N_XI0/XI46/XI10/NET34_XI0/XI46/XI10/MM4_g N_VDD_XI0/XI46/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI10/MM10 N_XI0/XI46/XI10/NET35_XI0/XI46/XI10/MM10_d
+ N_XI0/XI46/XI10/NET36_XI0/XI46/XI10/MM10_g N_VDD_XI0/XI46/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI10/MM11 N_XI0/XI46/XI10/NET36_XI0/XI46/XI10/MM11_d
+ N_XI0/XI46/XI10/NET35_XI0/XI46/XI10/MM11_g N_VDD_XI0/XI46/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI11/MM2 N_XI0/XI46/XI11/NET34_XI0/XI46/XI11/MM2_d
+ N_XI0/XI46/XI11/NET33_XI0/XI46/XI11/MM2_g N_VSS_XI0/XI46/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM3 N_XI0/XI46/XI11/NET33_XI0/XI46/XI11/MM3_d
+ N_WL<88>_XI0/XI46/XI11/MM3_g N_BLN<4>_XI0/XI46/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM0 N_XI0/XI46/XI11/NET34_XI0/XI46/XI11/MM0_d
+ N_WL<88>_XI0/XI46/XI11/MM0_g N_BL<4>_XI0/XI46/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM1 N_XI0/XI46/XI11/NET33_XI0/XI46/XI11/MM1_d
+ N_XI0/XI46/XI11/NET34_XI0/XI46/XI11/MM1_g N_VSS_XI0/XI46/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM9 N_XI0/XI46/XI11/NET36_XI0/XI46/XI11/MM9_d
+ N_WL<89>_XI0/XI46/XI11/MM9_g N_BL<4>_XI0/XI46/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM6 N_XI0/XI46/XI11/NET35_XI0/XI46/XI11/MM6_d
+ N_XI0/XI46/XI11/NET36_XI0/XI46/XI11/MM6_g N_VSS_XI0/XI46/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM7 N_XI0/XI46/XI11/NET36_XI0/XI46/XI11/MM7_d
+ N_XI0/XI46/XI11/NET35_XI0/XI46/XI11/MM7_g N_VSS_XI0/XI46/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM8 N_XI0/XI46/XI11/NET35_XI0/XI46/XI11/MM8_d
+ N_WL<89>_XI0/XI46/XI11/MM8_g N_BLN<4>_XI0/XI46/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI11/MM5 N_XI0/XI46/XI11/NET34_XI0/XI46/XI11/MM5_d
+ N_XI0/XI46/XI11/NET33_XI0/XI46/XI11/MM5_g N_VDD_XI0/XI46/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI11/MM4 N_XI0/XI46/XI11/NET33_XI0/XI46/XI11/MM4_d
+ N_XI0/XI46/XI11/NET34_XI0/XI46/XI11/MM4_g N_VDD_XI0/XI46/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI11/MM10 N_XI0/XI46/XI11/NET35_XI0/XI46/XI11/MM10_d
+ N_XI0/XI46/XI11/NET36_XI0/XI46/XI11/MM10_g N_VDD_XI0/XI46/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI11/MM11 N_XI0/XI46/XI11/NET36_XI0/XI46/XI11/MM11_d
+ N_XI0/XI46/XI11/NET35_XI0/XI46/XI11/MM11_g N_VDD_XI0/XI46/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI12/MM2 N_XI0/XI46/XI12/NET34_XI0/XI46/XI12/MM2_d
+ N_XI0/XI46/XI12/NET33_XI0/XI46/XI12/MM2_g N_VSS_XI0/XI46/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM3 N_XI0/XI46/XI12/NET33_XI0/XI46/XI12/MM3_d
+ N_WL<88>_XI0/XI46/XI12/MM3_g N_BLN<3>_XI0/XI46/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM0 N_XI0/XI46/XI12/NET34_XI0/XI46/XI12/MM0_d
+ N_WL<88>_XI0/XI46/XI12/MM0_g N_BL<3>_XI0/XI46/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM1 N_XI0/XI46/XI12/NET33_XI0/XI46/XI12/MM1_d
+ N_XI0/XI46/XI12/NET34_XI0/XI46/XI12/MM1_g N_VSS_XI0/XI46/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM9 N_XI0/XI46/XI12/NET36_XI0/XI46/XI12/MM9_d
+ N_WL<89>_XI0/XI46/XI12/MM9_g N_BL<3>_XI0/XI46/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM6 N_XI0/XI46/XI12/NET35_XI0/XI46/XI12/MM6_d
+ N_XI0/XI46/XI12/NET36_XI0/XI46/XI12/MM6_g N_VSS_XI0/XI46/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM7 N_XI0/XI46/XI12/NET36_XI0/XI46/XI12/MM7_d
+ N_XI0/XI46/XI12/NET35_XI0/XI46/XI12/MM7_g N_VSS_XI0/XI46/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM8 N_XI0/XI46/XI12/NET35_XI0/XI46/XI12/MM8_d
+ N_WL<89>_XI0/XI46/XI12/MM8_g N_BLN<3>_XI0/XI46/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI12/MM5 N_XI0/XI46/XI12/NET34_XI0/XI46/XI12/MM5_d
+ N_XI0/XI46/XI12/NET33_XI0/XI46/XI12/MM5_g N_VDD_XI0/XI46/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI12/MM4 N_XI0/XI46/XI12/NET33_XI0/XI46/XI12/MM4_d
+ N_XI0/XI46/XI12/NET34_XI0/XI46/XI12/MM4_g N_VDD_XI0/XI46/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI12/MM10 N_XI0/XI46/XI12/NET35_XI0/XI46/XI12/MM10_d
+ N_XI0/XI46/XI12/NET36_XI0/XI46/XI12/MM10_g N_VDD_XI0/XI46/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI12/MM11 N_XI0/XI46/XI12/NET36_XI0/XI46/XI12/MM11_d
+ N_XI0/XI46/XI12/NET35_XI0/XI46/XI12/MM11_g N_VDD_XI0/XI46/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI13/MM2 N_XI0/XI46/XI13/NET34_XI0/XI46/XI13/MM2_d
+ N_XI0/XI46/XI13/NET33_XI0/XI46/XI13/MM2_g N_VSS_XI0/XI46/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM3 N_XI0/XI46/XI13/NET33_XI0/XI46/XI13/MM3_d
+ N_WL<88>_XI0/XI46/XI13/MM3_g N_BLN<2>_XI0/XI46/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM0 N_XI0/XI46/XI13/NET34_XI0/XI46/XI13/MM0_d
+ N_WL<88>_XI0/XI46/XI13/MM0_g N_BL<2>_XI0/XI46/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM1 N_XI0/XI46/XI13/NET33_XI0/XI46/XI13/MM1_d
+ N_XI0/XI46/XI13/NET34_XI0/XI46/XI13/MM1_g N_VSS_XI0/XI46/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM9 N_XI0/XI46/XI13/NET36_XI0/XI46/XI13/MM9_d
+ N_WL<89>_XI0/XI46/XI13/MM9_g N_BL<2>_XI0/XI46/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM6 N_XI0/XI46/XI13/NET35_XI0/XI46/XI13/MM6_d
+ N_XI0/XI46/XI13/NET36_XI0/XI46/XI13/MM6_g N_VSS_XI0/XI46/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM7 N_XI0/XI46/XI13/NET36_XI0/XI46/XI13/MM7_d
+ N_XI0/XI46/XI13/NET35_XI0/XI46/XI13/MM7_g N_VSS_XI0/XI46/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM8 N_XI0/XI46/XI13/NET35_XI0/XI46/XI13/MM8_d
+ N_WL<89>_XI0/XI46/XI13/MM8_g N_BLN<2>_XI0/XI46/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI13/MM5 N_XI0/XI46/XI13/NET34_XI0/XI46/XI13/MM5_d
+ N_XI0/XI46/XI13/NET33_XI0/XI46/XI13/MM5_g N_VDD_XI0/XI46/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI13/MM4 N_XI0/XI46/XI13/NET33_XI0/XI46/XI13/MM4_d
+ N_XI0/XI46/XI13/NET34_XI0/XI46/XI13/MM4_g N_VDD_XI0/XI46/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI13/MM10 N_XI0/XI46/XI13/NET35_XI0/XI46/XI13/MM10_d
+ N_XI0/XI46/XI13/NET36_XI0/XI46/XI13/MM10_g N_VDD_XI0/XI46/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI13/MM11 N_XI0/XI46/XI13/NET36_XI0/XI46/XI13/MM11_d
+ N_XI0/XI46/XI13/NET35_XI0/XI46/XI13/MM11_g N_VDD_XI0/XI46/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI14/MM2 N_XI0/XI46/XI14/NET34_XI0/XI46/XI14/MM2_d
+ N_XI0/XI46/XI14/NET33_XI0/XI46/XI14/MM2_g N_VSS_XI0/XI46/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM3 N_XI0/XI46/XI14/NET33_XI0/XI46/XI14/MM3_d
+ N_WL<88>_XI0/XI46/XI14/MM3_g N_BLN<1>_XI0/XI46/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM0 N_XI0/XI46/XI14/NET34_XI0/XI46/XI14/MM0_d
+ N_WL<88>_XI0/XI46/XI14/MM0_g N_BL<1>_XI0/XI46/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM1 N_XI0/XI46/XI14/NET33_XI0/XI46/XI14/MM1_d
+ N_XI0/XI46/XI14/NET34_XI0/XI46/XI14/MM1_g N_VSS_XI0/XI46/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM9 N_XI0/XI46/XI14/NET36_XI0/XI46/XI14/MM9_d
+ N_WL<89>_XI0/XI46/XI14/MM9_g N_BL<1>_XI0/XI46/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM6 N_XI0/XI46/XI14/NET35_XI0/XI46/XI14/MM6_d
+ N_XI0/XI46/XI14/NET36_XI0/XI46/XI14/MM6_g N_VSS_XI0/XI46/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM7 N_XI0/XI46/XI14/NET36_XI0/XI46/XI14/MM7_d
+ N_XI0/XI46/XI14/NET35_XI0/XI46/XI14/MM7_g N_VSS_XI0/XI46/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM8 N_XI0/XI46/XI14/NET35_XI0/XI46/XI14/MM8_d
+ N_WL<89>_XI0/XI46/XI14/MM8_g N_BLN<1>_XI0/XI46/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI14/MM5 N_XI0/XI46/XI14/NET34_XI0/XI46/XI14/MM5_d
+ N_XI0/XI46/XI14/NET33_XI0/XI46/XI14/MM5_g N_VDD_XI0/XI46/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI14/MM4 N_XI0/XI46/XI14/NET33_XI0/XI46/XI14/MM4_d
+ N_XI0/XI46/XI14/NET34_XI0/XI46/XI14/MM4_g N_VDD_XI0/XI46/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI14/MM10 N_XI0/XI46/XI14/NET35_XI0/XI46/XI14/MM10_d
+ N_XI0/XI46/XI14/NET36_XI0/XI46/XI14/MM10_g N_VDD_XI0/XI46/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI14/MM11 N_XI0/XI46/XI14/NET36_XI0/XI46/XI14/MM11_d
+ N_XI0/XI46/XI14/NET35_XI0/XI46/XI14/MM11_g N_VDD_XI0/XI46/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI15/MM2 N_XI0/XI46/XI15/NET34_XI0/XI46/XI15/MM2_d
+ N_XI0/XI46/XI15/NET33_XI0/XI46/XI15/MM2_g N_VSS_XI0/XI46/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM3 N_XI0/XI46/XI15/NET33_XI0/XI46/XI15/MM3_d
+ N_WL<88>_XI0/XI46/XI15/MM3_g N_BLN<0>_XI0/XI46/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM0 N_XI0/XI46/XI15/NET34_XI0/XI46/XI15/MM0_d
+ N_WL<88>_XI0/XI46/XI15/MM0_g N_BL<0>_XI0/XI46/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM1 N_XI0/XI46/XI15/NET33_XI0/XI46/XI15/MM1_d
+ N_XI0/XI46/XI15/NET34_XI0/XI46/XI15/MM1_g N_VSS_XI0/XI46/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM9 N_XI0/XI46/XI15/NET36_XI0/XI46/XI15/MM9_d
+ N_WL<89>_XI0/XI46/XI15/MM9_g N_BL<0>_XI0/XI46/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM6 N_XI0/XI46/XI15/NET35_XI0/XI46/XI15/MM6_d
+ N_XI0/XI46/XI15/NET36_XI0/XI46/XI15/MM6_g N_VSS_XI0/XI46/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM7 N_XI0/XI46/XI15/NET36_XI0/XI46/XI15/MM7_d
+ N_XI0/XI46/XI15/NET35_XI0/XI46/XI15/MM7_g N_VSS_XI0/XI46/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM8 N_XI0/XI46/XI15/NET35_XI0/XI46/XI15/MM8_d
+ N_WL<89>_XI0/XI46/XI15/MM8_g N_BLN<0>_XI0/XI46/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI46/XI15/MM5 N_XI0/XI46/XI15/NET34_XI0/XI46/XI15/MM5_d
+ N_XI0/XI46/XI15/NET33_XI0/XI46/XI15/MM5_g N_VDD_XI0/XI46/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI15/MM4 N_XI0/XI46/XI15/NET33_XI0/XI46/XI15/MM4_d
+ N_XI0/XI46/XI15/NET34_XI0/XI46/XI15/MM4_g N_VDD_XI0/XI46/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI15/MM10 N_XI0/XI46/XI15/NET35_XI0/XI46/XI15/MM10_d
+ N_XI0/XI46/XI15/NET36_XI0/XI46/XI15/MM10_g N_VDD_XI0/XI46/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI46/XI15/MM11 N_XI0/XI46/XI15/NET36_XI0/XI46/XI15/MM11_d
+ N_XI0/XI46/XI15/NET35_XI0/XI46/XI15/MM11_g N_VDD_XI0/XI46/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI0/MM2 N_XI0/XI47/XI0/NET34_XI0/XI47/XI0/MM2_d
+ N_XI0/XI47/XI0/NET33_XI0/XI47/XI0/MM2_g N_VSS_XI0/XI47/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM3 N_XI0/XI47/XI0/NET33_XI0/XI47/XI0/MM3_d
+ N_WL<90>_XI0/XI47/XI0/MM3_g N_BLN<15>_XI0/XI47/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM0 N_XI0/XI47/XI0/NET34_XI0/XI47/XI0/MM0_d
+ N_WL<90>_XI0/XI47/XI0/MM0_g N_BL<15>_XI0/XI47/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM1 N_XI0/XI47/XI0/NET33_XI0/XI47/XI0/MM1_d
+ N_XI0/XI47/XI0/NET34_XI0/XI47/XI0/MM1_g N_VSS_XI0/XI47/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM9 N_XI0/XI47/XI0/NET36_XI0/XI47/XI0/MM9_d
+ N_WL<91>_XI0/XI47/XI0/MM9_g N_BL<15>_XI0/XI47/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM6 N_XI0/XI47/XI0/NET35_XI0/XI47/XI0/MM6_d
+ N_XI0/XI47/XI0/NET36_XI0/XI47/XI0/MM6_g N_VSS_XI0/XI47/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM7 N_XI0/XI47/XI0/NET36_XI0/XI47/XI0/MM7_d
+ N_XI0/XI47/XI0/NET35_XI0/XI47/XI0/MM7_g N_VSS_XI0/XI47/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM8 N_XI0/XI47/XI0/NET35_XI0/XI47/XI0/MM8_d
+ N_WL<91>_XI0/XI47/XI0/MM8_g N_BLN<15>_XI0/XI47/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI0/MM5 N_XI0/XI47/XI0/NET34_XI0/XI47/XI0/MM5_d
+ N_XI0/XI47/XI0/NET33_XI0/XI47/XI0/MM5_g N_VDD_XI0/XI47/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI0/MM4 N_XI0/XI47/XI0/NET33_XI0/XI47/XI0/MM4_d
+ N_XI0/XI47/XI0/NET34_XI0/XI47/XI0/MM4_g N_VDD_XI0/XI47/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI0/MM10 N_XI0/XI47/XI0/NET35_XI0/XI47/XI0/MM10_d
+ N_XI0/XI47/XI0/NET36_XI0/XI47/XI0/MM10_g N_VDD_XI0/XI47/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI0/MM11 N_XI0/XI47/XI0/NET36_XI0/XI47/XI0/MM11_d
+ N_XI0/XI47/XI0/NET35_XI0/XI47/XI0/MM11_g N_VDD_XI0/XI47/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI1/MM2 N_XI0/XI47/XI1/NET34_XI0/XI47/XI1/MM2_d
+ N_XI0/XI47/XI1/NET33_XI0/XI47/XI1/MM2_g N_VSS_XI0/XI47/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM3 N_XI0/XI47/XI1/NET33_XI0/XI47/XI1/MM3_d
+ N_WL<90>_XI0/XI47/XI1/MM3_g N_BLN<14>_XI0/XI47/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM0 N_XI0/XI47/XI1/NET34_XI0/XI47/XI1/MM0_d
+ N_WL<90>_XI0/XI47/XI1/MM0_g N_BL<14>_XI0/XI47/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM1 N_XI0/XI47/XI1/NET33_XI0/XI47/XI1/MM1_d
+ N_XI0/XI47/XI1/NET34_XI0/XI47/XI1/MM1_g N_VSS_XI0/XI47/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM9 N_XI0/XI47/XI1/NET36_XI0/XI47/XI1/MM9_d
+ N_WL<91>_XI0/XI47/XI1/MM9_g N_BL<14>_XI0/XI47/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM6 N_XI0/XI47/XI1/NET35_XI0/XI47/XI1/MM6_d
+ N_XI0/XI47/XI1/NET36_XI0/XI47/XI1/MM6_g N_VSS_XI0/XI47/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM7 N_XI0/XI47/XI1/NET36_XI0/XI47/XI1/MM7_d
+ N_XI0/XI47/XI1/NET35_XI0/XI47/XI1/MM7_g N_VSS_XI0/XI47/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM8 N_XI0/XI47/XI1/NET35_XI0/XI47/XI1/MM8_d
+ N_WL<91>_XI0/XI47/XI1/MM8_g N_BLN<14>_XI0/XI47/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI1/MM5 N_XI0/XI47/XI1/NET34_XI0/XI47/XI1/MM5_d
+ N_XI0/XI47/XI1/NET33_XI0/XI47/XI1/MM5_g N_VDD_XI0/XI47/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI1/MM4 N_XI0/XI47/XI1/NET33_XI0/XI47/XI1/MM4_d
+ N_XI0/XI47/XI1/NET34_XI0/XI47/XI1/MM4_g N_VDD_XI0/XI47/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI1/MM10 N_XI0/XI47/XI1/NET35_XI0/XI47/XI1/MM10_d
+ N_XI0/XI47/XI1/NET36_XI0/XI47/XI1/MM10_g N_VDD_XI0/XI47/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI1/MM11 N_XI0/XI47/XI1/NET36_XI0/XI47/XI1/MM11_d
+ N_XI0/XI47/XI1/NET35_XI0/XI47/XI1/MM11_g N_VDD_XI0/XI47/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI2/MM2 N_XI0/XI47/XI2/NET34_XI0/XI47/XI2/MM2_d
+ N_XI0/XI47/XI2/NET33_XI0/XI47/XI2/MM2_g N_VSS_XI0/XI47/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM3 N_XI0/XI47/XI2/NET33_XI0/XI47/XI2/MM3_d
+ N_WL<90>_XI0/XI47/XI2/MM3_g N_BLN<13>_XI0/XI47/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM0 N_XI0/XI47/XI2/NET34_XI0/XI47/XI2/MM0_d
+ N_WL<90>_XI0/XI47/XI2/MM0_g N_BL<13>_XI0/XI47/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM1 N_XI0/XI47/XI2/NET33_XI0/XI47/XI2/MM1_d
+ N_XI0/XI47/XI2/NET34_XI0/XI47/XI2/MM1_g N_VSS_XI0/XI47/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM9 N_XI0/XI47/XI2/NET36_XI0/XI47/XI2/MM9_d
+ N_WL<91>_XI0/XI47/XI2/MM9_g N_BL<13>_XI0/XI47/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM6 N_XI0/XI47/XI2/NET35_XI0/XI47/XI2/MM6_d
+ N_XI0/XI47/XI2/NET36_XI0/XI47/XI2/MM6_g N_VSS_XI0/XI47/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM7 N_XI0/XI47/XI2/NET36_XI0/XI47/XI2/MM7_d
+ N_XI0/XI47/XI2/NET35_XI0/XI47/XI2/MM7_g N_VSS_XI0/XI47/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM8 N_XI0/XI47/XI2/NET35_XI0/XI47/XI2/MM8_d
+ N_WL<91>_XI0/XI47/XI2/MM8_g N_BLN<13>_XI0/XI47/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI2/MM5 N_XI0/XI47/XI2/NET34_XI0/XI47/XI2/MM5_d
+ N_XI0/XI47/XI2/NET33_XI0/XI47/XI2/MM5_g N_VDD_XI0/XI47/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI2/MM4 N_XI0/XI47/XI2/NET33_XI0/XI47/XI2/MM4_d
+ N_XI0/XI47/XI2/NET34_XI0/XI47/XI2/MM4_g N_VDD_XI0/XI47/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI2/MM10 N_XI0/XI47/XI2/NET35_XI0/XI47/XI2/MM10_d
+ N_XI0/XI47/XI2/NET36_XI0/XI47/XI2/MM10_g N_VDD_XI0/XI47/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI2/MM11 N_XI0/XI47/XI2/NET36_XI0/XI47/XI2/MM11_d
+ N_XI0/XI47/XI2/NET35_XI0/XI47/XI2/MM11_g N_VDD_XI0/XI47/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI3/MM2 N_XI0/XI47/XI3/NET34_XI0/XI47/XI3/MM2_d
+ N_XI0/XI47/XI3/NET33_XI0/XI47/XI3/MM2_g N_VSS_XI0/XI47/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM3 N_XI0/XI47/XI3/NET33_XI0/XI47/XI3/MM3_d
+ N_WL<90>_XI0/XI47/XI3/MM3_g N_BLN<12>_XI0/XI47/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM0 N_XI0/XI47/XI3/NET34_XI0/XI47/XI3/MM0_d
+ N_WL<90>_XI0/XI47/XI3/MM0_g N_BL<12>_XI0/XI47/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM1 N_XI0/XI47/XI3/NET33_XI0/XI47/XI3/MM1_d
+ N_XI0/XI47/XI3/NET34_XI0/XI47/XI3/MM1_g N_VSS_XI0/XI47/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM9 N_XI0/XI47/XI3/NET36_XI0/XI47/XI3/MM9_d
+ N_WL<91>_XI0/XI47/XI3/MM9_g N_BL<12>_XI0/XI47/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM6 N_XI0/XI47/XI3/NET35_XI0/XI47/XI3/MM6_d
+ N_XI0/XI47/XI3/NET36_XI0/XI47/XI3/MM6_g N_VSS_XI0/XI47/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM7 N_XI0/XI47/XI3/NET36_XI0/XI47/XI3/MM7_d
+ N_XI0/XI47/XI3/NET35_XI0/XI47/XI3/MM7_g N_VSS_XI0/XI47/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM8 N_XI0/XI47/XI3/NET35_XI0/XI47/XI3/MM8_d
+ N_WL<91>_XI0/XI47/XI3/MM8_g N_BLN<12>_XI0/XI47/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI3/MM5 N_XI0/XI47/XI3/NET34_XI0/XI47/XI3/MM5_d
+ N_XI0/XI47/XI3/NET33_XI0/XI47/XI3/MM5_g N_VDD_XI0/XI47/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI3/MM4 N_XI0/XI47/XI3/NET33_XI0/XI47/XI3/MM4_d
+ N_XI0/XI47/XI3/NET34_XI0/XI47/XI3/MM4_g N_VDD_XI0/XI47/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI3/MM10 N_XI0/XI47/XI3/NET35_XI0/XI47/XI3/MM10_d
+ N_XI0/XI47/XI3/NET36_XI0/XI47/XI3/MM10_g N_VDD_XI0/XI47/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI3/MM11 N_XI0/XI47/XI3/NET36_XI0/XI47/XI3/MM11_d
+ N_XI0/XI47/XI3/NET35_XI0/XI47/XI3/MM11_g N_VDD_XI0/XI47/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI4/MM2 N_XI0/XI47/XI4/NET34_XI0/XI47/XI4/MM2_d
+ N_XI0/XI47/XI4/NET33_XI0/XI47/XI4/MM2_g N_VSS_XI0/XI47/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM3 N_XI0/XI47/XI4/NET33_XI0/XI47/XI4/MM3_d
+ N_WL<90>_XI0/XI47/XI4/MM3_g N_BLN<11>_XI0/XI47/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM0 N_XI0/XI47/XI4/NET34_XI0/XI47/XI4/MM0_d
+ N_WL<90>_XI0/XI47/XI4/MM0_g N_BL<11>_XI0/XI47/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM1 N_XI0/XI47/XI4/NET33_XI0/XI47/XI4/MM1_d
+ N_XI0/XI47/XI4/NET34_XI0/XI47/XI4/MM1_g N_VSS_XI0/XI47/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM9 N_XI0/XI47/XI4/NET36_XI0/XI47/XI4/MM9_d
+ N_WL<91>_XI0/XI47/XI4/MM9_g N_BL<11>_XI0/XI47/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM6 N_XI0/XI47/XI4/NET35_XI0/XI47/XI4/MM6_d
+ N_XI0/XI47/XI4/NET36_XI0/XI47/XI4/MM6_g N_VSS_XI0/XI47/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM7 N_XI0/XI47/XI4/NET36_XI0/XI47/XI4/MM7_d
+ N_XI0/XI47/XI4/NET35_XI0/XI47/XI4/MM7_g N_VSS_XI0/XI47/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM8 N_XI0/XI47/XI4/NET35_XI0/XI47/XI4/MM8_d
+ N_WL<91>_XI0/XI47/XI4/MM8_g N_BLN<11>_XI0/XI47/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI4/MM5 N_XI0/XI47/XI4/NET34_XI0/XI47/XI4/MM5_d
+ N_XI0/XI47/XI4/NET33_XI0/XI47/XI4/MM5_g N_VDD_XI0/XI47/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI4/MM4 N_XI0/XI47/XI4/NET33_XI0/XI47/XI4/MM4_d
+ N_XI0/XI47/XI4/NET34_XI0/XI47/XI4/MM4_g N_VDD_XI0/XI47/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI4/MM10 N_XI0/XI47/XI4/NET35_XI0/XI47/XI4/MM10_d
+ N_XI0/XI47/XI4/NET36_XI0/XI47/XI4/MM10_g N_VDD_XI0/XI47/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI4/MM11 N_XI0/XI47/XI4/NET36_XI0/XI47/XI4/MM11_d
+ N_XI0/XI47/XI4/NET35_XI0/XI47/XI4/MM11_g N_VDD_XI0/XI47/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI5/MM2 N_XI0/XI47/XI5/NET34_XI0/XI47/XI5/MM2_d
+ N_XI0/XI47/XI5/NET33_XI0/XI47/XI5/MM2_g N_VSS_XI0/XI47/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM3 N_XI0/XI47/XI5/NET33_XI0/XI47/XI5/MM3_d
+ N_WL<90>_XI0/XI47/XI5/MM3_g N_BLN<10>_XI0/XI47/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM0 N_XI0/XI47/XI5/NET34_XI0/XI47/XI5/MM0_d
+ N_WL<90>_XI0/XI47/XI5/MM0_g N_BL<10>_XI0/XI47/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM1 N_XI0/XI47/XI5/NET33_XI0/XI47/XI5/MM1_d
+ N_XI0/XI47/XI5/NET34_XI0/XI47/XI5/MM1_g N_VSS_XI0/XI47/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM9 N_XI0/XI47/XI5/NET36_XI0/XI47/XI5/MM9_d
+ N_WL<91>_XI0/XI47/XI5/MM9_g N_BL<10>_XI0/XI47/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM6 N_XI0/XI47/XI5/NET35_XI0/XI47/XI5/MM6_d
+ N_XI0/XI47/XI5/NET36_XI0/XI47/XI5/MM6_g N_VSS_XI0/XI47/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM7 N_XI0/XI47/XI5/NET36_XI0/XI47/XI5/MM7_d
+ N_XI0/XI47/XI5/NET35_XI0/XI47/XI5/MM7_g N_VSS_XI0/XI47/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM8 N_XI0/XI47/XI5/NET35_XI0/XI47/XI5/MM8_d
+ N_WL<91>_XI0/XI47/XI5/MM8_g N_BLN<10>_XI0/XI47/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI5/MM5 N_XI0/XI47/XI5/NET34_XI0/XI47/XI5/MM5_d
+ N_XI0/XI47/XI5/NET33_XI0/XI47/XI5/MM5_g N_VDD_XI0/XI47/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI5/MM4 N_XI0/XI47/XI5/NET33_XI0/XI47/XI5/MM4_d
+ N_XI0/XI47/XI5/NET34_XI0/XI47/XI5/MM4_g N_VDD_XI0/XI47/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI5/MM10 N_XI0/XI47/XI5/NET35_XI0/XI47/XI5/MM10_d
+ N_XI0/XI47/XI5/NET36_XI0/XI47/XI5/MM10_g N_VDD_XI0/XI47/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI5/MM11 N_XI0/XI47/XI5/NET36_XI0/XI47/XI5/MM11_d
+ N_XI0/XI47/XI5/NET35_XI0/XI47/XI5/MM11_g N_VDD_XI0/XI47/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI6/MM2 N_XI0/XI47/XI6/NET34_XI0/XI47/XI6/MM2_d
+ N_XI0/XI47/XI6/NET33_XI0/XI47/XI6/MM2_g N_VSS_XI0/XI47/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM3 N_XI0/XI47/XI6/NET33_XI0/XI47/XI6/MM3_d
+ N_WL<90>_XI0/XI47/XI6/MM3_g N_BLN<9>_XI0/XI47/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM0 N_XI0/XI47/XI6/NET34_XI0/XI47/XI6/MM0_d
+ N_WL<90>_XI0/XI47/XI6/MM0_g N_BL<9>_XI0/XI47/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM1 N_XI0/XI47/XI6/NET33_XI0/XI47/XI6/MM1_d
+ N_XI0/XI47/XI6/NET34_XI0/XI47/XI6/MM1_g N_VSS_XI0/XI47/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM9 N_XI0/XI47/XI6/NET36_XI0/XI47/XI6/MM9_d
+ N_WL<91>_XI0/XI47/XI6/MM9_g N_BL<9>_XI0/XI47/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM6 N_XI0/XI47/XI6/NET35_XI0/XI47/XI6/MM6_d
+ N_XI0/XI47/XI6/NET36_XI0/XI47/XI6/MM6_g N_VSS_XI0/XI47/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM7 N_XI0/XI47/XI6/NET36_XI0/XI47/XI6/MM7_d
+ N_XI0/XI47/XI6/NET35_XI0/XI47/XI6/MM7_g N_VSS_XI0/XI47/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM8 N_XI0/XI47/XI6/NET35_XI0/XI47/XI6/MM8_d
+ N_WL<91>_XI0/XI47/XI6/MM8_g N_BLN<9>_XI0/XI47/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI6/MM5 N_XI0/XI47/XI6/NET34_XI0/XI47/XI6/MM5_d
+ N_XI0/XI47/XI6/NET33_XI0/XI47/XI6/MM5_g N_VDD_XI0/XI47/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI6/MM4 N_XI0/XI47/XI6/NET33_XI0/XI47/XI6/MM4_d
+ N_XI0/XI47/XI6/NET34_XI0/XI47/XI6/MM4_g N_VDD_XI0/XI47/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI6/MM10 N_XI0/XI47/XI6/NET35_XI0/XI47/XI6/MM10_d
+ N_XI0/XI47/XI6/NET36_XI0/XI47/XI6/MM10_g N_VDD_XI0/XI47/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI6/MM11 N_XI0/XI47/XI6/NET36_XI0/XI47/XI6/MM11_d
+ N_XI0/XI47/XI6/NET35_XI0/XI47/XI6/MM11_g N_VDD_XI0/XI47/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI7/MM2 N_XI0/XI47/XI7/NET34_XI0/XI47/XI7/MM2_d
+ N_XI0/XI47/XI7/NET33_XI0/XI47/XI7/MM2_g N_VSS_XI0/XI47/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM3 N_XI0/XI47/XI7/NET33_XI0/XI47/XI7/MM3_d
+ N_WL<90>_XI0/XI47/XI7/MM3_g N_BLN<8>_XI0/XI47/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM0 N_XI0/XI47/XI7/NET34_XI0/XI47/XI7/MM0_d
+ N_WL<90>_XI0/XI47/XI7/MM0_g N_BL<8>_XI0/XI47/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM1 N_XI0/XI47/XI7/NET33_XI0/XI47/XI7/MM1_d
+ N_XI0/XI47/XI7/NET34_XI0/XI47/XI7/MM1_g N_VSS_XI0/XI47/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM9 N_XI0/XI47/XI7/NET36_XI0/XI47/XI7/MM9_d
+ N_WL<91>_XI0/XI47/XI7/MM9_g N_BL<8>_XI0/XI47/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM6 N_XI0/XI47/XI7/NET35_XI0/XI47/XI7/MM6_d
+ N_XI0/XI47/XI7/NET36_XI0/XI47/XI7/MM6_g N_VSS_XI0/XI47/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM7 N_XI0/XI47/XI7/NET36_XI0/XI47/XI7/MM7_d
+ N_XI0/XI47/XI7/NET35_XI0/XI47/XI7/MM7_g N_VSS_XI0/XI47/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM8 N_XI0/XI47/XI7/NET35_XI0/XI47/XI7/MM8_d
+ N_WL<91>_XI0/XI47/XI7/MM8_g N_BLN<8>_XI0/XI47/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI7/MM5 N_XI0/XI47/XI7/NET34_XI0/XI47/XI7/MM5_d
+ N_XI0/XI47/XI7/NET33_XI0/XI47/XI7/MM5_g N_VDD_XI0/XI47/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI7/MM4 N_XI0/XI47/XI7/NET33_XI0/XI47/XI7/MM4_d
+ N_XI0/XI47/XI7/NET34_XI0/XI47/XI7/MM4_g N_VDD_XI0/XI47/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI7/MM10 N_XI0/XI47/XI7/NET35_XI0/XI47/XI7/MM10_d
+ N_XI0/XI47/XI7/NET36_XI0/XI47/XI7/MM10_g N_VDD_XI0/XI47/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI7/MM11 N_XI0/XI47/XI7/NET36_XI0/XI47/XI7/MM11_d
+ N_XI0/XI47/XI7/NET35_XI0/XI47/XI7/MM11_g N_VDD_XI0/XI47/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI8/MM2 N_XI0/XI47/XI8/NET34_XI0/XI47/XI8/MM2_d
+ N_XI0/XI47/XI8/NET33_XI0/XI47/XI8/MM2_g N_VSS_XI0/XI47/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM3 N_XI0/XI47/XI8/NET33_XI0/XI47/XI8/MM3_d
+ N_WL<90>_XI0/XI47/XI8/MM3_g N_BLN<7>_XI0/XI47/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM0 N_XI0/XI47/XI8/NET34_XI0/XI47/XI8/MM0_d
+ N_WL<90>_XI0/XI47/XI8/MM0_g N_BL<7>_XI0/XI47/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM1 N_XI0/XI47/XI8/NET33_XI0/XI47/XI8/MM1_d
+ N_XI0/XI47/XI8/NET34_XI0/XI47/XI8/MM1_g N_VSS_XI0/XI47/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM9 N_XI0/XI47/XI8/NET36_XI0/XI47/XI8/MM9_d
+ N_WL<91>_XI0/XI47/XI8/MM9_g N_BL<7>_XI0/XI47/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM6 N_XI0/XI47/XI8/NET35_XI0/XI47/XI8/MM6_d
+ N_XI0/XI47/XI8/NET36_XI0/XI47/XI8/MM6_g N_VSS_XI0/XI47/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM7 N_XI0/XI47/XI8/NET36_XI0/XI47/XI8/MM7_d
+ N_XI0/XI47/XI8/NET35_XI0/XI47/XI8/MM7_g N_VSS_XI0/XI47/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM8 N_XI0/XI47/XI8/NET35_XI0/XI47/XI8/MM8_d
+ N_WL<91>_XI0/XI47/XI8/MM8_g N_BLN<7>_XI0/XI47/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI8/MM5 N_XI0/XI47/XI8/NET34_XI0/XI47/XI8/MM5_d
+ N_XI0/XI47/XI8/NET33_XI0/XI47/XI8/MM5_g N_VDD_XI0/XI47/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI8/MM4 N_XI0/XI47/XI8/NET33_XI0/XI47/XI8/MM4_d
+ N_XI0/XI47/XI8/NET34_XI0/XI47/XI8/MM4_g N_VDD_XI0/XI47/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI8/MM10 N_XI0/XI47/XI8/NET35_XI0/XI47/XI8/MM10_d
+ N_XI0/XI47/XI8/NET36_XI0/XI47/XI8/MM10_g N_VDD_XI0/XI47/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI8/MM11 N_XI0/XI47/XI8/NET36_XI0/XI47/XI8/MM11_d
+ N_XI0/XI47/XI8/NET35_XI0/XI47/XI8/MM11_g N_VDD_XI0/XI47/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI9/MM2 N_XI0/XI47/XI9/NET34_XI0/XI47/XI9/MM2_d
+ N_XI0/XI47/XI9/NET33_XI0/XI47/XI9/MM2_g N_VSS_XI0/XI47/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM3 N_XI0/XI47/XI9/NET33_XI0/XI47/XI9/MM3_d
+ N_WL<90>_XI0/XI47/XI9/MM3_g N_BLN<6>_XI0/XI47/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM0 N_XI0/XI47/XI9/NET34_XI0/XI47/XI9/MM0_d
+ N_WL<90>_XI0/XI47/XI9/MM0_g N_BL<6>_XI0/XI47/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM1 N_XI0/XI47/XI9/NET33_XI0/XI47/XI9/MM1_d
+ N_XI0/XI47/XI9/NET34_XI0/XI47/XI9/MM1_g N_VSS_XI0/XI47/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM9 N_XI0/XI47/XI9/NET36_XI0/XI47/XI9/MM9_d
+ N_WL<91>_XI0/XI47/XI9/MM9_g N_BL<6>_XI0/XI47/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM6 N_XI0/XI47/XI9/NET35_XI0/XI47/XI9/MM6_d
+ N_XI0/XI47/XI9/NET36_XI0/XI47/XI9/MM6_g N_VSS_XI0/XI47/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM7 N_XI0/XI47/XI9/NET36_XI0/XI47/XI9/MM7_d
+ N_XI0/XI47/XI9/NET35_XI0/XI47/XI9/MM7_g N_VSS_XI0/XI47/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM8 N_XI0/XI47/XI9/NET35_XI0/XI47/XI9/MM8_d
+ N_WL<91>_XI0/XI47/XI9/MM8_g N_BLN<6>_XI0/XI47/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI9/MM5 N_XI0/XI47/XI9/NET34_XI0/XI47/XI9/MM5_d
+ N_XI0/XI47/XI9/NET33_XI0/XI47/XI9/MM5_g N_VDD_XI0/XI47/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI9/MM4 N_XI0/XI47/XI9/NET33_XI0/XI47/XI9/MM4_d
+ N_XI0/XI47/XI9/NET34_XI0/XI47/XI9/MM4_g N_VDD_XI0/XI47/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI9/MM10 N_XI0/XI47/XI9/NET35_XI0/XI47/XI9/MM10_d
+ N_XI0/XI47/XI9/NET36_XI0/XI47/XI9/MM10_g N_VDD_XI0/XI47/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI9/MM11 N_XI0/XI47/XI9/NET36_XI0/XI47/XI9/MM11_d
+ N_XI0/XI47/XI9/NET35_XI0/XI47/XI9/MM11_g N_VDD_XI0/XI47/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI10/MM2 N_XI0/XI47/XI10/NET34_XI0/XI47/XI10/MM2_d
+ N_XI0/XI47/XI10/NET33_XI0/XI47/XI10/MM2_g N_VSS_XI0/XI47/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM3 N_XI0/XI47/XI10/NET33_XI0/XI47/XI10/MM3_d
+ N_WL<90>_XI0/XI47/XI10/MM3_g N_BLN<5>_XI0/XI47/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM0 N_XI0/XI47/XI10/NET34_XI0/XI47/XI10/MM0_d
+ N_WL<90>_XI0/XI47/XI10/MM0_g N_BL<5>_XI0/XI47/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM1 N_XI0/XI47/XI10/NET33_XI0/XI47/XI10/MM1_d
+ N_XI0/XI47/XI10/NET34_XI0/XI47/XI10/MM1_g N_VSS_XI0/XI47/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM9 N_XI0/XI47/XI10/NET36_XI0/XI47/XI10/MM9_d
+ N_WL<91>_XI0/XI47/XI10/MM9_g N_BL<5>_XI0/XI47/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM6 N_XI0/XI47/XI10/NET35_XI0/XI47/XI10/MM6_d
+ N_XI0/XI47/XI10/NET36_XI0/XI47/XI10/MM6_g N_VSS_XI0/XI47/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM7 N_XI0/XI47/XI10/NET36_XI0/XI47/XI10/MM7_d
+ N_XI0/XI47/XI10/NET35_XI0/XI47/XI10/MM7_g N_VSS_XI0/XI47/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM8 N_XI0/XI47/XI10/NET35_XI0/XI47/XI10/MM8_d
+ N_WL<91>_XI0/XI47/XI10/MM8_g N_BLN<5>_XI0/XI47/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI10/MM5 N_XI0/XI47/XI10/NET34_XI0/XI47/XI10/MM5_d
+ N_XI0/XI47/XI10/NET33_XI0/XI47/XI10/MM5_g N_VDD_XI0/XI47/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI10/MM4 N_XI0/XI47/XI10/NET33_XI0/XI47/XI10/MM4_d
+ N_XI0/XI47/XI10/NET34_XI0/XI47/XI10/MM4_g N_VDD_XI0/XI47/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI10/MM10 N_XI0/XI47/XI10/NET35_XI0/XI47/XI10/MM10_d
+ N_XI0/XI47/XI10/NET36_XI0/XI47/XI10/MM10_g N_VDD_XI0/XI47/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI10/MM11 N_XI0/XI47/XI10/NET36_XI0/XI47/XI10/MM11_d
+ N_XI0/XI47/XI10/NET35_XI0/XI47/XI10/MM11_g N_VDD_XI0/XI47/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI11/MM2 N_XI0/XI47/XI11/NET34_XI0/XI47/XI11/MM2_d
+ N_XI0/XI47/XI11/NET33_XI0/XI47/XI11/MM2_g N_VSS_XI0/XI47/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM3 N_XI0/XI47/XI11/NET33_XI0/XI47/XI11/MM3_d
+ N_WL<90>_XI0/XI47/XI11/MM3_g N_BLN<4>_XI0/XI47/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM0 N_XI0/XI47/XI11/NET34_XI0/XI47/XI11/MM0_d
+ N_WL<90>_XI0/XI47/XI11/MM0_g N_BL<4>_XI0/XI47/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM1 N_XI0/XI47/XI11/NET33_XI0/XI47/XI11/MM1_d
+ N_XI0/XI47/XI11/NET34_XI0/XI47/XI11/MM1_g N_VSS_XI0/XI47/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM9 N_XI0/XI47/XI11/NET36_XI0/XI47/XI11/MM9_d
+ N_WL<91>_XI0/XI47/XI11/MM9_g N_BL<4>_XI0/XI47/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM6 N_XI0/XI47/XI11/NET35_XI0/XI47/XI11/MM6_d
+ N_XI0/XI47/XI11/NET36_XI0/XI47/XI11/MM6_g N_VSS_XI0/XI47/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM7 N_XI0/XI47/XI11/NET36_XI0/XI47/XI11/MM7_d
+ N_XI0/XI47/XI11/NET35_XI0/XI47/XI11/MM7_g N_VSS_XI0/XI47/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM8 N_XI0/XI47/XI11/NET35_XI0/XI47/XI11/MM8_d
+ N_WL<91>_XI0/XI47/XI11/MM8_g N_BLN<4>_XI0/XI47/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI11/MM5 N_XI0/XI47/XI11/NET34_XI0/XI47/XI11/MM5_d
+ N_XI0/XI47/XI11/NET33_XI0/XI47/XI11/MM5_g N_VDD_XI0/XI47/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI11/MM4 N_XI0/XI47/XI11/NET33_XI0/XI47/XI11/MM4_d
+ N_XI0/XI47/XI11/NET34_XI0/XI47/XI11/MM4_g N_VDD_XI0/XI47/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI11/MM10 N_XI0/XI47/XI11/NET35_XI0/XI47/XI11/MM10_d
+ N_XI0/XI47/XI11/NET36_XI0/XI47/XI11/MM10_g N_VDD_XI0/XI47/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI11/MM11 N_XI0/XI47/XI11/NET36_XI0/XI47/XI11/MM11_d
+ N_XI0/XI47/XI11/NET35_XI0/XI47/XI11/MM11_g N_VDD_XI0/XI47/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI12/MM2 N_XI0/XI47/XI12/NET34_XI0/XI47/XI12/MM2_d
+ N_XI0/XI47/XI12/NET33_XI0/XI47/XI12/MM2_g N_VSS_XI0/XI47/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM3 N_XI0/XI47/XI12/NET33_XI0/XI47/XI12/MM3_d
+ N_WL<90>_XI0/XI47/XI12/MM3_g N_BLN<3>_XI0/XI47/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM0 N_XI0/XI47/XI12/NET34_XI0/XI47/XI12/MM0_d
+ N_WL<90>_XI0/XI47/XI12/MM0_g N_BL<3>_XI0/XI47/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM1 N_XI0/XI47/XI12/NET33_XI0/XI47/XI12/MM1_d
+ N_XI0/XI47/XI12/NET34_XI0/XI47/XI12/MM1_g N_VSS_XI0/XI47/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM9 N_XI0/XI47/XI12/NET36_XI0/XI47/XI12/MM9_d
+ N_WL<91>_XI0/XI47/XI12/MM9_g N_BL<3>_XI0/XI47/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM6 N_XI0/XI47/XI12/NET35_XI0/XI47/XI12/MM6_d
+ N_XI0/XI47/XI12/NET36_XI0/XI47/XI12/MM6_g N_VSS_XI0/XI47/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM7 N_XI0/XI47/XI12/NET36_XI0/XI47/XI12/MM7_d
+ N_XI0/XI47/XI12/NET35_XI0/XI47/XI12/MM7_g N_VSS_XI0/XI47/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM8 N_XI0/XI47/XI12/NET35_XI0/XI47/XI12/MM8_d
+ N_WL<91>_XI0/XI47/XI12/MM8_g N_BLN<3>_XI0/XI47/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI12/MM5 N_XI0/XI47/XI12/NET34_XI0/XI47/XI12/MM5_d
+ N_XI0/XI47/XI12/NET33_XI0/XI47/XI12/MM5_g N_VDD_XI0/XI47/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI12/MM4 N_XI0/XI47/XI12/NET33_XI0/XI47/XI12/MM4_d
+ N_XI0/XI47/XI12/NET34_XI0/XI47/XI12/MM4_g N_VDD_XI0/XI47/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI12/MM10 N_XI0/XI47/XI12/NET35_XI0/XI47/XI12/MM10_d
+ N_XI0/XI47/XI12/NET36_XI0/XI47/XI12/MM10_g N_VDD_XI0/XI47/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI12/MM11 N_XI0/XI47/XI12/NET36_XI0/XI47/XI12/MM11_d
+ N_XI0/XI47/XI12/NET35_XI0/XI47/XI12/MM11_g N_VDD_XI0/XI47/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI13/MM2 N_XI0/XI47/XI13/NET34_XI0/XI47/XI13/MM2_d
+ N_XI0/XI47/XI13/NET33_XI0/XI47/XI13/MM2_g N_VSS_XI0/XI47/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM3 N_XI0/XI47/XI13/NET33_XI0/XI47/XI13/MM3_d
+ N_WL<90>_XI0/XI47/XI13/MM3_g N_BLN<2>_XI0/XI47/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM0 N_XI0/XI47/XI13/NET34_XI0/XI47/XI13/MM0_d
+ N_WL<90>_XI0/XI47/XI13/MM0_g N_BL<2>_XI0/XI47/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM1 N_XI0/XI47/XI13/NET33_XI0/XI47/XI13/MM1_d
+ N_XI0/XI47/XI13/NET34_XI0/XI47/XI13/MM1_g N_VSS_XI0/XI47/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM9 N_XI0/XI47/XI13/NET36_XI0/XI47/XI13/MM9_d
+ N_WL<91>_XI0/XI47/XI13/MM9_g N_BL<2>_XI0/XI47/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM6 N_XI0/XI47/XI13/NET35_XI0/XI47/XI13/MM6_d
+ N_XI0/XI47/XI13/NET36_XI0/XI47/XI13/MM6_g N_VSS_XI0/XI47/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM7 N_XI0/XI47/XI13/NET36_XI0/XI47/XI13/MM7_d
+ N_XI0/XI47/XI13/NET35_XI0/XI47/XI13/MM7_g N_VSS_XI0/XI47/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM8 N_XI0/XI47/XI13/NET35_XI0/XI47/XI13/MM8_d
+ N_WL<91>_XI0/XI47/XI13/MM8_g N_BLN<2>_XI0/XI47/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI13/MM5 N_XI0/XI47/XI13/NET34_XI0/XI47/XI13/MM5_d
+ N_XI0/XI47/XI13/NET33_XI0/XI47/XI13/MM5_g N_VDD_XI0/XI47/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI13/MM4 N_XI0/XI47/XI13/NET33_XI0/XI47/XI13/MM4_d
+ N_XI0/XI47/XI13/NET34_XI0/XI47/XI13/MM4_g N_VDD_XI0/XI47/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI13/MM10 N_XI0/XI47/XI13/NET35_XI0/XI47/XI13/MM10_d
+ N_XI0/XI47/XI13/NET36_XI0/XI47/XI13/MM10_g N_VDD_XI0/XI47/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI13/MM11 N_XI0/XI47/XI13/NET36_XI0/XI47/XI13/MM11_d
+ N_XI0/XI47/XI13/NET35_XI0/XI47/XI13/MM11_g N_VDD_XI0/XI47/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI14/MM2 N_XI0/XI47/XI14/NET34_XI0/XI47/XI14/MM2_d
+ N_XI0/XI47/XI14/NET33_XI0/XI47/XI14/MM2_g N_VSS_XI0/XI47/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM3 N_XI0/XI47/XI14/NET33_XI0/XI47/XI14/MM3_d
+ N_WL<90>_XI0/XI47/XI14/MM3_g N_BLN<1>_XI0/XI47/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM0 N_XI0/XI47/XI14/NET34_XI0/XI47/XI14/MM0_d
+ N_WL<90>_XI0/XI47/XI14/MM0_g N_BL<1>_XI0/XI47/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM1 N_XI0/XI47/XI14/NET33_XI0/XI47/XI14/MM1_d
+ N_XI0/XI47/XI14/NET34_XI0/XI47/XI14/MM1_g N_VSS_XI0/XI47/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM9 N_XI0/XI47/XI14/NET36_XI0/XI47/XI14/MM9_d
+ N_WL<91>_XI0/XI47/XI14/MM9_g N_BL<1>_XI0/XI47/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM6 N_XI0/XI47/XI14/NET35_XI0/XI47/XI14/MM6_d
+ N_XI0/XI47/XI14/NET36_XI0/XI47/XI14/MM6_g N_VSS_XI0/XI47/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM7 N_XI0/XI47/XI14/NET36_XI0/XI47/XI14/MM7_d
+ N_XI0/XI47/XI14/NET35_XI0/XI47/XI14/MM7_g N_VSS_XI0/XI47/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM8 N_XI0/XI47/XI14/NET35_XI0/XI47/XI14/MM8_d
+ N_WL<91>_XI0/XI47/XI14/MM8_g N_BLN<1>_XI0/XI47/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI14/MM5 N_XI0/XI47/XI14/NET34_XI0/XI47/XI14/MM5_d
+ N_XI0/XI47/XI14/NET33_XI0/XI47/XI14/MM5_g N_VDD_XI0/XI47/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI14/MM4 N_XI0/XI47/XI14/NET33_XI0/XI47/XI14/MM4_d
+ N_XI0/XI47/XI14/NET34_XI0/XI47/XI14/MM4_g N_VDD_XI0/XI47/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI14/MM10 N_XI0/XI47/XI14/NET35_XI0/XI47/XI14/MM10_d
+ N_XI0/XI47/XI14/NET36_XI0/XI47/XI14/MM10_g N_VDD_XI0/XI47/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI14/MM11 N_XI0/XI47/XI14/NET36_XI0/XI47/XI14/MM11_d
+ N_XI0/XI47/XI14/NET35_XI0/XI47/XI14/MM11_g N_VDD_XI0/XI47/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI15/MM2 N_XI0/XI47/XI15/NET34_XI0/XI47/XI15/MM2_d
+ N_XI0/XI47/XI15/NET33_XI0/XI47/XI15/MM2_g N_VSS_XI0/XI47/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM3 N_XI0/XI47/XI15/NET33_XI0/XI47/XI15/MM3_d
+ N_WL<90>_XI0/XI47/XI15/MM3_g N_BLN<0>_XI0/XI47/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM0 N_XI0/XI47/XI15/NET34_XI0/XI47/XI15/MM0_d
+ N_WL<90>_XI0/XI47/XI15/MM0_g N_BL<0>_XI0/XI47/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM1 N_XI0/XI47/XI15/NET33_XI0/XI47/XI15/MM1_d
+ N_XI0/XI47/XI15/NET34_XI0/XI47/XI15/MM1_g N_VSS_XI0/XI47/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM9 N_XI0/XI47/XI15/NET36_XI0/XI47/XI15/MM9_d
+ N_WL<91>_XI0/XI47/XI15/MM9_g N_BL<0>_XI0/XI47/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM6 N_XI0/XI47/XI15/NET35_XI0/XI47/XI15/MM6_d
+ N_XI0/XI47/XI15/NET36_XI0/XI47/XI15/MM6_g N_VSS_XI0/XI47/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM7 N_XI0/XI47/XI15/NET36_XI0/XI47/XI15/MM7_d
+ N_XI0/XI47/XI15/NET35_XI0/XI47/XI15/MM7_g N_VSS_XI0/XI47/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM8 N_XI0/XI47/XI15/NET35_XI0/XI47/XI15/MM8_d
+ N_WL<91>_XI0/XI47/XI15/MM8_g N_BLN<0>_XI0/XI47/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI47/XI15/MM5 N_XI0/XI47/XI15/NET34_XI0/XI47/XI15/MM5_d
+ N_XI0/XI47/XI15/NET33_XI0/XI47/XI15/MM5_g N_VDD_XI0/XI47/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI15/MM4 N_XI0/XI47/XI15/NET33_XI0/XI47/XI15/MM4_d
+ N_XI0/XI47/XI15/NET34_XI0/XI47/XI15/MM4_g N_VDD_XI0/XI47/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI15/MM10 N_XI0/XI47/XI15/NET35_XI0/XI47/XI15/MM10_d
+ N_XI0/XI47/XI15/NET36_XI0/XI47/XI15/MM10_g N_VDD_XI0/XI47/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI47/XI15/MM11 N_XI0/XI47/XI15/NET36_XI0/XI47/XI15/MM11_d
+ N_XI0/XI47/XI15/NET35_XI0/XI47/XI15/MM11_g N_VDD_XI0/XI47/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI0/MM2 N_XI0/XI48/XI0/NET34_XI0/XI48/XI0/MM2_d
+ N_XI0/XI48/XI0/NET33_XI0/XI48/XI0/MM2_g N_VSS_XI0/XI48/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM3 N_XI0/XI48/XI0/NET33_XI0/XI48/XI0/MM3_d
+ N_WL<92>_XI0/XI48/XI0/MM3_g N_BLN<15>_XI0/XI48/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM0 N_XI0/XI48/XI0/NET34_XI0/XI48/XI0/MM0_d
+ N_WL<92>_XI0/XI48/XI0/MM0_g N_BL<15>_XI0/XI48/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM1 N_XI0/XI48/XI0/NET33_XI0/XI48/XI0/MM1_d
+ N_XI0/XI48/XI0/NET34_XI0/XI48/XI0/MM1_g N_VSS_XI0/XI48/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM9 N_XI0/XI48/XI0/NET36_XI0/XI48/XI0/MM9_d
+ N_WL<93>_XI0/XI48/XI0/MM9_g N_BL<15>_XI0/XI48/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM6 N_XI0/XI48/XI0/NET35_XI0/XI48/XI0/MM6_d
+ N_XI0/XI48/XI0/NET36_XI0/XI48/XI0/MM6_g N_VSS_XI0/XI48/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM7 N_XI0/XI48/XI0/NET36_XI0/XI48/XI0/MM7_d
+ N_XI0/XI48/XI0/NET35_XI0/XI48/XI0/MM7_g N_VSS_XI0/XI48/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM8 N_XI0/XI48/XI0/NET35_XI0/XI48/XI0/MM8_d
+ N_WL<93>_XI0/XI48/XI0/MM8_g N_BLN<15>_XI0/XI48/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI0/MM5 N_XI0/XI48/XI0/NET34_XI0/XI48/XI0/MM5_d
+ N_XI0/XI48/XI0/NET33_XI0/XI48/XI0/MM5_g N_VDD_XI0/XI48/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI0/MM4 N_XI0/XI48/XI0/NET33_XI0/XI48/XI0/MM4_d
+ N_XI0/XI48/XI0/NET34_XI0/XI48/XI0/MM4_g N_VDD_XI0/XI48/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI0/MM10 N_XI0/XI48/XI0/NET35_XI0/XI48/XI0/MM10_d
+ N_XI0/XI48/XI0/NET36_XI0/XI48/XI0/MM10_g N_VDD_XI0/XI48/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI0/MM11 N_XI0/XI48/XI0/NET36_XI0/XI48/XI0/MM11_d
+ N_XI0/XI48/XI0/NET35_XI0/XI48/XI0/MM11_g N_VDD_XI0/XI48/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI1/MM2 N_XI0/XI48/XI1/NET34_XI0/XI48/XI1/MM2_d
+ N_XI0/XI48/XI1/NET33_XI0/XI48/XI1/MM2_g N_VSS_XI0/XI48/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM3 N_XI0/XI48/XI1/NET33_XI0/XI48/XI1/MM3_d
+ N_WL<92>_XI0/XI48/XI1/MM3_g N_BLN<14>_XI0/XI48/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM0 N_XI0/XI48/XI1/NET34_XI0/XI48/XI1/MM0_d
+ N_WL<92>_XI0/XI48/XI1/MM0_g N_BL<14>_XI0/XI48/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM1 N_XI0/XI48/XI1/NET33_XI0/XI48/XI1/MM1_d
+ N_XI0/XI48/XI1/NET34_XI0/XI48/XI1/MM1_g N_VSS_XI0/XI48/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM9 N_XI0/XI48/XI1/NET36_XI0/XI48/XI1/MM9_d
+ N_WL<93>_XI0/XI48/XI1/MM9_g N_BL<14>_XI0/XI48/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM6 N_XI0/XI48/XI1/NET35_XI0/XI48/XI1/MM6_d
+ N_XI0/XI48/XI1/NET36_XI0/XI48/XI1/MM6_g N_VSS_XI0/XI48/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM7 N_XI0/XI48/XI1/NET36_XI0/XI48/XI1/MM7_d
+ N_XI0/XI48/XI1/NET35_XI0/XI48/XI1/MM7_g N_VSS_XI0/XI48/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM8 N_XI0/XI48/XI1/NET35_XI0/XI48/XI1/MM8_d
+ N_WL<93>_XI0/XI48/XI1/MM8_g N_BLN<14>_XI0/XI48/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI1/MM5 N_XI0/XI48/XI1/NET34_XI0/XI48/XI1/MM5_d
+ N_XI0/XI48/XI1/NET33_XI0/XI48/XI1/MM5_g N_VDD_XI0/XI48/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI1/MM4 N_XI0/XI48/XI1/NET33_XI0/XI48/XI1/MM4_d
+ N_XI0/XI48/XI1/NET34_XI0/XI48/XI1/MM4_g N_VDD_XI0/XI48/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI1/MM10 N_XI0/XI48/XI1/NET35_XI0/XI48/XI1/MM10_d
+ N_XI0/XI48/XI1/NET36_XI0/XI48/XI1/MM10_g N_VDD_XI0/XI48/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI1/MM11 N_XI0/XI48/XI1/NET36_XI0/XI48/XI1/MM11_d
+ N_XI0/XI48/XI1/NET35_XI0/XI48/XI1/MM11_g N_VDD_XI0/XI48/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI2/MM2 N_XI0/XI48/XI2/NET34_XI0/XI48/XI2/MM2_d
+ N_XI0/XI48/XI2/NET33_XI0/XI48/XI2/MM2_g N_VSS_XI0/XI48/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM3 N_XI0/XI48/XI2/NET33_XI0/XI48/XI2/MM3_d
+ N_WL<92>_XI0/XI48/XI2/MM3_g N_BLN<13>_XI0/XI48/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM0 N_XI0/XI48/XI2/NET34_XI0/XI48/XI2/MM0_d
+ N_WL<92>_XI0/XI48/XI2/MM0_g N_BL<13>_XI0/XI48/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM1 N_XI0/XI48/XI2/NET33_XI0/XI48/XI2/MM1_d
+ N_XI0/XI48/XI2/NET34_XI0/XI48/XI2/MM1_g N_VSS_XI0/XI48/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM9 N_XI0/XI48/XI2/NET36_XI0/XI48/XI2/MM9_d
+ N_WL<93>_XI0/XI48/XI2/MM9_g N_BL<13>_XI0/XI48/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM6 N_XI0/XI48/XI2/NET35_XI0/XI48/XI2/MM6_d
+ N_XI0/XI48/XI2/NET36_XI0/XI48/XI2/MM6_g N_VSS_XI0/XI48/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM7 N_XI0/XI48/XI2/NET36_XI0/XI48/XI2/MM7_d
+ N_XI0/XI48/XI2/NET35_XI0/XI48/XI2/MM7_g N_VSS_XI0/XI48/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM8 N_XI0/XI48/XI2/NET35_XI0/XI48/XI2/MM8_d
+ N_WL<93>_XI0/XI48/XI2/MM8_g N_BLN<13>_XI0/XI48/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI2/MM5 N_XI0/XI48/XI2/NET34_XI0/XI48/XI2/MM5_d
+ N_XI0/XI48/XI2/NET33_XI0/XI48/XI2/MM5_g N_VDD_XI0/XI48/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI2/MM4 N_XI0/XI48/XI2/NET33_XI0/XI48/XI2/MM4_d
+ N_XI0/XI48/XI2/NET34_XI0/XI48/XI2/MM4_g N_VDD_XI0/XI48/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI2/MM10 N_XI0/XI48/XI2/NET35_XI0/XI48/XI2/MM10_d
+ N_XI0/XI48/XI2/NET36_XI0/XI48/XI2/MM10_g N_VDD_XI0/XI48/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI2/MM11 N_XI0/XI48/XI2/NET36_XI0/XI48/XI2/MM11_d
+ N_XI0/XI48/XI2/NET35_XI0/XI48/XI2/MM11_g N_VDD_XI0/XI48/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI3/MM2 N_XI0/XI48/XI3/NET34_XI0/XI48/XI3/MM2_d
+ N_XI0/XI48/XI3/NET33_XI0/XI48/XI3/MM2_g N_VSS_XI0/XI48/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM3 N_XI0/XI48/XI3/NET33_XI0/XI48/XI3/MM3_d
+ N_WL<92>_XI0/XI48/XI3/MM3_g N_BLN<12>_XI0/XI48/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM0 N_XI0/XI48/XI3/NET34_XI0/XI48/XI3/MM0_d
+ N_WL<92>_XI0/XI48/XI3/MM0_g N_BL<12>_XI0/XI48/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM1 N_XI0/XI48/XI3/NET33_XI0/XI48/XI3/MM1_d
+ N_XI0/XI48/XI3/NET34_XI0/XI48/XI3/MM1_g N_VSS_XI0/XI48/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM9 N_XI0/XI48/XI3/NET36_XI0/XI48/XI3/MM9_d
+ N_WL<93>_XI0/XI48/XI3/MM9_g N_BL<12>_XI0/XI48/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM6 N_XI0/XI48/XI3/NET35_XI0/XI48/XI3/MM6_d
+ N_XI0/XI48/XI3/NET36_XI0/XI48/XI3/MM6_g N_VSS_XI0/XI48/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM7 N_XI0/XI48/XI3/NET36_XI0/XI48/XI3/MM7_d
+ N_XI0/XI48/XI3/NET35_XI0/XI48/XI3/MM7_g N_VSS_XI0/XI48/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM8 N_XI0/XI48/XI3/NET35_XI0/XI48/XI3/MM8_d
+ N_WL<93>_XI0/XI48/XI3/MM8_g N_BLN<12>_XI0/XI48/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI3/MM5 N_XI0/XI48/XI3/NET34_XI0/XI48/XI3/MM5_d
+ N_XI0/XI48/XI3/NET33_XI0/XI48/XI3/MM5_g N_VDD_XI0/XI48/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI3/MM4 N_XI0/XI48/XI3/NET33_XI0/XI48/XI3/MM4_d
+ N_XI0/XI48/XI3/NET34_XI0/XI48/XI3/MM4_g N_VDD_XI0/XI48/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI3/MM10 N_XI0/XI48/XI3/NET35_XI0/XI48/XI3/MM10_d
+ N_XI0/XI48/XI3/NET36_XI0/XI48/XI3/MM10_g N_VDD_XI0/XI48/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI3/MM11 N_XI0/XI48/XI3/NET36_XI0/XI48/XI3/MM11_d
+ N_XI0/XI48/XI3/NET35_XI0/XI48/XI3/MM11_g N_VDD_XI0/XI48/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI4/MM2 N_XI0/XI48/XI4/NET34_XI0/XI48/XI4/MM2_d
+ N_XI0/XI48/XI4/NET33_XI0/XI48/XI4/MM2_g N_VSS_XI0/XI48/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM3 N_XI0/XI48/XI4/NET33_XI0/XI48/XI4/MM3_d
+ N_WL<92>_XI0/XI48/XI4/MM3_g N_BLN<11>_XI0/XI48/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM0 N_XI0/XI48/XI4/NET34_XI0/XI48/XI4/MM0_d
+ N_WL<92>_XI0/XI48/XI4/MM0_g N_BL<11>_XI0/XI48/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM1 N_XI0/XI48/XI4/NET33_XI0/XI48/XI4/MM1_d
+ N_XI0/XI48/XI4/NET34_XI0/XI48/XI4/MM1_g N_VSS_XI0/XI48/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM9 N_XI0/XI48/XI4/NET36_XI0/XI48/XI4/MM9_d
+ N_WL<93>_XI0/XI48/XI4/MM9_g N_BL<11>_XI0/XI48/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM6 N_XI0/XI48/XI4/NET35_XI0/XI48/XI4/MM6_d
+ N_XI0/XI48/XI4/NET36_XI0/XI48/XI4/MM6_g N_VSS_XI0/XI48/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM7 N_XI0/XI48/XI4/NET36_XI0/XI48/XI4/MM7_d
+ N_XI0/XI48/XI4/NET35_XI0/XI48/XI4/MM7_g N_VSS_XI0/XI48/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM8 N_XI0/XI48/XI4/NET35_XI0/XI48/XI4/MM8_d
+ N_WL<93>_XI0/XI48/XI4/MM8_g N_BLN<11>_XI0/XI48/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI4/MM5 N_XI0/XI48/XI4/NET34_XI0/XI48/XI4/MM5_d
+ N_XI0/XI48/XI4/NET33_XI0/XI48/XI4/MM5_g N_VDD_XI0/XI48/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI4/MM4 N_XI0/XI48/XI4/NET33_XI0/XI48/XI4/MM4_d
+ N_XI0/XI48/XI4/NET34_XI0/XI48/XI4/MM4_g N_VDD_XI0/XI48/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI4/MM10 N_XI0/XI48/XI4/NET35_XI0/XI48/XI4/MM10_d
+ N_XI0/XI48/XI4/NET36_XI0/XI48/XI4/MM10_g N_VDD_XI0/XI48/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI4/MM11 N_XI0/XI48/XI4/NET36_XI0/XI48/XI4/MM11_d
+ N_XI0/XI48/XI4/NET35_XI0/XI48/XI4/MM11_g N_VDD_XI0/XI48/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI5/MM2 N_XI0/XI48/XI5/NET34_XI0/XI48/XI5/MM2_d
+ N_XI0/XI48/XI5/NET33_XI0/XI48/XI5/MM2_g N_VSS_XI0/XI48/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM3 N_XI0/XI48/XI5/NET33_XI0/XI48/XI5/MM3_d
+ N_WL<92>_XI0/XI48/XI5/MM3_g N_BLN<10>_XI0/XI48/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM0 N_XI0/XI48/XI5/NET34_XI0/XI48/XI5/MM0_d
+ N_WL<92>_XI0/XI48/XI5/MM0_g N_BL<10>_XI0/XI48/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM1 N_XI0/XI48/XI5/NET33_XI0/XI48/XI5/MM1_d
+ N_XI0/XI48/XI5/NET34_XI0/XI48/XI5/MM1_g N_VSS_XI0/XI48/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM9 N_XI0/XI48/XI5/NET36_XI0/XI48/XI5/MM9_d
+ N_WL<93>_XI0/XI48/XI5/MM9_g N_BL<10>_XI0/XI48/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM6 N_XI0/XI48/XI5/NET35_XI0/XI48/XI5/MM6_d
+ N_XI0/XI48/XI5/NET36_XI0/XI48/XI5/MM6_g N_VSS_XI0/XI48/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM7 N_XI0/XI48/XI5/NET36_XI0/XI48/XI5/MM7_d
+ N_XI0/XI48/XI5/NET35_XI0/XI48/XI5/MM7_g N_VSS_XI0/XI48/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM8 N_XI0/XI48/XI5/NET35_XI0/XI48/XI5/MM8_d
+ N_WL<93>_XI0/XI48/XI5/MM8_g N_BLN<10>_XI0/XI48/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI5/MM5 N_XI0/XI48/XI5/NET34_XI0/XI48/XI5/MM5_d
+ N_XI0/XI48/XI5/NET33_XI0/XI48/XI5/MM5_g N_VDD_XI0/XI48/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI5/MM4 N_XI0/XI48/XI5/NET33_XI0/XI48/XI5/MM4_d
+ N_XI0/XI48/XI5/NET34_XI0/XI48/XI5/MM4_g N_VDD_XI0/XI48/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI5/MM10 N_XI0/XI48/XI5/NET35_XI0/XI48/XI5/MM10_d
+ N_XI0/XI48/XI5/NET36_XI0/XI48/XI5/MM10_g N_VDD_XI0/XI48/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI5/MM11 N_XI0/XI48/XI5/NET36_XI0/XI48/XI5/MM11_d
+ N_XI0/XI48/XI5/NET35_XI0/XI48/XI5/MM11_g N_VDD_XI0/XI48/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI6/MM2 N_XI0/XI48/XI6/NET34_XI0/XI48/XI6/MM2_d
+ N_XI0/XI48/XI6/NET33_XI0/XI48/XI6/MM2_g N_VSS_XI0/XI48/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM3 N_XI0/XI48/XI6/NET33_XI0/XI48/XI6/MM3_d
+ N_WL<92>_XI0/XI48/XI6/MM3_g N_BLN<9>_XI0/XI48/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM0 N_XI0/XI48/XI6/NET34_XI0/XI48/XI6/MM0_d
+ N_WL<92>_XI0/XI48/XI6/MM0_g N_BL<9>_XI0/XI48/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM1 N_XI0/XI48/XI6/NET33_XI0/XI48/XI6/MM1_d
+ N_XI0/XI48/XI6/NET34_XI0/XI48/XI6/MM1_g N_VSS_XI0/XI48/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM9 N_XI0/XI48/XI6/NET36_XI0/XI48/XI6/MM9_d
+ N_WL<93>_XI0/XI48/XI6/MM9_g N_BL<9>_XI0/XI48/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM6 N_XI0/XI48/XI6/NET35_XI0/XI48/XI6/MM6_d
+ N_XI0/XI48/XI6/NET36_XI0/XI48/XI6/MM6_g N_VSS_XI0/XI48/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM7 N_XI0/XI48/XI6/NET36_XI0/XI48/XI6/MM7_d
+ N_XI0/XI48/XI6/NET35_XI0/XI48/XI6/MM7_g N_VSS_XI0/XI48/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM8 N_XI0/XI48/XI6/NET35_XI0/XI48/XI6/MM8_d
+ N_WL<93>_XI0/XI48/XI6/MM8_g N_BLN<9>_XI0/XI48/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI6/MM5 N_XI0/XI48/XI6/NET34_XI0/XI48/XI6/MM5_d
+ N_XI0/XI48/XI6/NET33_XI0/XI48/XI6/MM5_g N_VDD_XI0/XI48/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI6/MM4 N_XI0/XI48/XI6/NET33_XI0/XI48/XI6/MM4_d
+ N_XI0/XI48/XI6/NET34_XI0/XI48/XI6/MM4_g N_VDD_XI0/XI48/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI6/MM10 N_XI0/XI48/XI6/NET35_XI0/XI48/XI6/MM10_d
+ N_XI0/XI48/XI6/NET36_XI0/XI48/XI6/MM10_g N_VDD_XI0/XI48/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI6/MM11 N_XI0/XI48/XI6/NET36_XI0/XI48/XI6/MM11_d
+ N_XI0/XI48/XI6/NET35_XI0/XI48/XI6/MM11_g N_VDD_XI0/XI48/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI7/MM2 N_XI0/XI48/XI7/NET34_XI0/XI48/XI7/MM2_d
+ N_XI0/XI48/XI7/NET33_XI0/XI48/XI7/MM2_g N_VSS_XI0/XI48/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM3 N_XI0/XI48/XI7/NET33_XI0/XI48/XI7/MM3_d
+ N_WL<92>_XI0/XI48/XI7/MM3_g N_BLN<8>_XI0/XI48/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM0 N_XI0/XI48/XI7/NET34_XI0/XI48/XI7/MM0_d
+ N_WL<92>_XI0/XI48/XI7/MM0_g N_BL<8>_XI0/XI48/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM1 N_XI0/XI48/XI7/NET33_XI0/XI48/XI7/MM1_d
+ N_XI0/XI48/XI7/NET34_XI0/XI48/XI7/MM1_g N_VSS_XI0/XI48/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM9 N_XI0/XI48/XI7/NET36_XI0/XI48/XI7/MM9_d
+ N_WL<93>_XI0/XI48/XI7/MM9_g N_BL<8>_XI0/XI48/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM6 N_XI0/XI48/XI7/NET35_XI0/XI48/XI7/MM6_d
+ N_XI0/XI48/XI7/NET36_XI0/XI48/XI7/MM6_g N_VSS_XI0/XI48/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM7 N_XI0/XI48/XI7/NET36_XI0/XI48/XI7/MM7_d
+ N_XI0/XI48/XI7/NET35_XI0/XI48/XI7/MM7_g N_VSS_XI0/XI48/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM8 N_XI0/XI48/XI7/NET35_XI0/XI48/XI7/MM8_d
+ N_WL<93>_XI0/XI48/XI7/MM8_g N_BLN<8>_XI0/XI48/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI7/MM5 N_XI0/XI48/XI7/NET34_XI0/XI48/XI7/MM5_d
+ N_XI0/XI48/XI7/NET33_XI0/XI48/XI7/MM5_g N_VDD_XI0/XI48/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI7/MM4 N_XI0/XI48/XI7/NET33_XI0/XI48/XI7/MM4_d
+ N_XI0/XI48/XI7/NET34_XI0/XI48/XI7/MM4_g N_VDD_XI0/XI48/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI7/MM10 N_XI0/XI48/XI7/NET35_XI0/XI48/XI7/MM10_d
+ N_XI0/XI48/XI7/NET36_XI0/XI48/XI7/MM10_g N_VDD_XI0/XI48/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI7/MM11 N_XI0/XI48/XI7/NET36_XI0/XI48/XI7/MM11_d
+ N_XI0/XI48/XI7/NET35_XI0/XI48/XI7/MM11_g N_VDD_XI0/XI48/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI8/MM2 N_XI0/XI48/XI8/NET34_XI0/XI48/XI8/MM2_d
+ N_XI0/XI48/XI8/NET33_XI0/XI48/XI8/MM2_g N_VSS_XI0/XI48/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM3 N_XI0/XI48/XI8/NET33_XI0/XI48/XI8/MM3_d
+ N_WL<92>_XI0/XI48/XI8/MM3_g N_BLN<7>_XI0/XI48/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM0 N_XI0/XI48/XI8/NET34_XI0/XI48/XI8/MM0_d
+ N_WL<92>_XI0/XI48/XI8/MM0_g N_BL<7>_XI0/XI48/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM1 N_XI0/XI48/XI8/NET33_XI0/XI48/XI8/MM1_d
+ N_XI0/XI48/XI8/NET34_XI0/XI48/XI8/MM1_g N_VSS_XI0/XI48/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM9 N_XI0/XI48/XI8/NET36_XI0/XI48/XI8/MM9_d
+ N_WL<93>_XI0/XI48/XI8/MM9_g N_BL<7>_XI0/XI48/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM6 N_XI0/XI48/XI8/NET35_XI0/XI48/XI8/MM6_d
+ N_XI0/XI48/XI8/NET36_XI0/XI48/XI8/MM6_g N_VSS_XI0/XI48/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM7 N_XI0/XI48/XI8/NET36_XI0/XI48/XI8/MM7_d
+ N_XI0/XI48/XI8/NET35_XI0/XI48/XI8/MM7_g N_VSS_XI0/XI48/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM8 N_XI0/XI48/XI8/NET35_XI0/XI48/XI8/MM8_d
+ N_WL<93>_XI0/XI48/XI8/MM8_g N_BLN<7>_XI0/XI48/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI8/MM5 N_XI0/XI48/XI8/NET34_XI0/XI48/XI8/MM5_d
+ N_XI0/XI48/XI8/NET33_XI0/XI48/XI8/MM5_g N_VDD_XI0/XI48/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI8/MM4 N_XI0/XI48/XI8/NET33_XI0/XI48/XI8/MM4_d
+ N_XI0/XI48/XI8/NET34_XI0/XI48/XI8/MM4_g N_VDD_XI0/XI48/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI8/MM10 N_XI0/XI48/XI8/NET35_XI0/XI48/XI8/MM10_d
+ N_XI0/XI48/XI8/NET36_XI0/XI48/XI8/MM10_g N_VDD_XI0/XI48/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI8/MM11 N_XI0/XI48/XI8/NET36_XI0/XI48/XI8/MM11_d
+ N_XI0/XI48/XI8/NET35_XI0/XI48/XI8/MM11_g N_VDD_XI0/XI48/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI9/MM2 N_XI0/XI48/XI9/NET34_XI0/XI48/XI9/MM2_d
+ N_XI0/XI48/XI9/NET33_XI0/XI48/XI9/MM2_g N_VSS_XI0/XI48/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM3 N_XI0/XI48/XI9/NET33_XI0/XI48/XI9/MM3_d
+ N_WL<92>_XI0/XI48/XI9/MM3_g N_BLN<6>_XI0/XI48/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM0 N_XI0/XI48/XI9/NET34_XI0/XI48/XI9/MM0_d
+ N_WL<92>_XI0/XI48/XI9/MM0_g N_BL<6>_XI0/XI48/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM1 N_XI0/XI48/XI9/NET33_XI0/XI48/XI9/MM1_d
+ N_XI0/XI48/XI9/NET34_XI0/XI48/XI9/MM1_g N_VSS_XI0/XI48/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM9 N_XI0/XI48/XI9/NET36_XI0/XI48/XI9/MM9_d
+ N_WL<93>_XI0/XI48/XI9/MM9_g N_BL<6>_XI0/XI48/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM6 N_XI0/XI48/XI9/NET35_XI0/XI48/XI9/MM6_d
+ N_XI0/XI48/XI9/NET36_XI0/XI48/XI9/MM6_g N_VSS_XI0/XI48/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM7 N_XI0/XI48/XI9/NET36_XI0/XI48/XI9/MM7_d
+ N_XI0/XI48/XI9/NET35_XI0/XI48/XI9/MM7_g N_VSS_XI0/XI48/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM8 N_XI0/XI48/XI9/NET35_XI0/XI48/XI9/MM8_d
+ N_WL<93>_XI0/XI48/XI9/MM8_g N_BLN<6>_XI0/XI48/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI9/MM5 N_XI0/XI48/XI9/NET34_XI0/XI48/XI9/MM5_d
+ N_XI0/XI48/XI9/NET33_XI0/XI48/XI9/MM5_g N_VDD_XI0/XI48/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI9/MM4 N_XI0/XI48/XI9/NET33_XI0/XI48/XI9/MM4_d
+ N_XI0/XI48/XI9/NET34_XI0/XI48/XI9/MM4_g N_VDD_XI0/XI48/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI9/MM10 N_XI0/XI48/XI9/NET35_XI0/XI48/XI9/MM10_d
+ N_XI0/XI48/XI9/NET36_XI0/XI48/XI9/MM10_g N_VDD_XI0/XI48/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI9/MM11 N_XI0/XI48/XI9/NET36_XI0/XI48/XI9/MM11_d
+ N_XI0/XI48/XI9/NET35_XI0/XI48/XI9/MM11_g N_VDD_XI0/XI48/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI10/MM2 N_XI0/XI48/XI10/NET34_XI0/XI48/XI10/MM2_d
+ N_XI0/XI48/XI10/NET33_XI0/XI48/XI10/MM2_g N_VSS_XI0/XI48/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM3 N_XI0/XI48/XI10/NET33_XI0/XI48/XI10/MM3_d
+ N_WL<92>_XI0/XI48/XI10/MM3_g N_BLN<5>_XI0/XI48/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM0 N_XI0/XI48/XI10/NET34_XI0/XI48/XI10/MM0_d
+ N_WL<92>_XI0/XI48/XI10/MM0_g N_BL<5>_XI0/XI48/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM1 N_XI0/XI48/XI10/NET33_XI0/XI48/XI10/MM1_d
+ N_XI0/XI48/XI10/NET34_XI0/XI48/XI10/MM1_g N_VSS_XI0/XI48/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM9 N_XI0/XI48/XI10/NET36_XI0/XI48/XI10/MM9_d
+ N_WL<93>_XI0/XI48/XI10/MM9_g N_BL<5>_XI0/XI48/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM6 N_XI0/XI48/XI10/NET35_XI0/XI48/XI10/MM6_d
+ N_XI0/XI48/XI10/NET36_XI0/XI48/XI10/MM6_g N_VSS_XI0/XI48/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM7 N_XI0/XI48/XI10/NET36_XI0/XI48/XI10/MM7_d
+ N_XI0/XI48/XI10/NET35_XI0/XI48/XI10/MM7_g N_VSS_XI0/XI48/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM8 N_XI0/XI48/XI10/NET35_XI0/XI48/XI10/MM8_d
+ N_WL<93>_XI0/XI48/XI10/MM8_g N_BLN<5>_XI0/XI48/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI10/MM5 N_XI0/XI48/XI10/NET34_XI0/XI48/XI10/MM5_d
+ N_XI0/XI48/XI10/NET33_XI0/XI48/XI10/MM5_g N_VDD_XI0/XI48/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI10/MM4 N_XI0/XI48/XI10/NET33_XI0/XI48/XI10/MM4_d
+ N_XI0/XI48/XI10/NET34_XI0/XI48/XI10/MM4_g N_VDD_XI0/XI48/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI10/MM10 N_XI0/XI48/XI10/NET35_XI0/XI48/XI10/MM10_d
+ N_XI0/XI48/XI10/NET36_XI0/XI48/XI10/MM10_g N_VDD_XI0/XI48/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI10/MM11 N_XI0/XI48/XI10/NET36_XI0/XI48/XI10/MM11_d
+ N_XI0/XI48/XI10/NET35_XI0/XI48/XI10/MM11_g N_VDD_XI0/XI48/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI11/MM2 N_XI0/XI48/XI11/NET34_XI0/XI48/XI11/MM2_d
+ N_XI0/XI48/XI11/NET33_XI0/XI48/XI11/MM2_g N_VSS_XI0/XI48/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM3 N_XI0/XI48/XI11/NET33_XI0/XI48/XI11/MM3_d
+ N_WL<92>_XI0/XI48/XI11/MM3_g N_BLN<4>_XI0/XI48/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM0 N_XI0/XI48/XI11/NET34_XI0/XI48/XI11/MM0_d
+ N_WL<92>_XI0/XI48/XI11/MM0_g N_BL<4>_XI0/XI48/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM1 N_XI0/XI48/XI11/NET33_XI0/XI48/XI11/MM1_d
+ N_XI0/XI48/XI11/NET34_XI0/XI48/XI11/MM1_g N_VSS_XI0/XI48/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM9 N_XI0/XI48/XI11/NET36_XI0/XI48/XI11/MM9_d
+ N_WL<93>_XI0/XI48/XI11/MM9_g N_BL<4>_XI0/XI48/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM6 N_XI0/XI48/XI11/NET35_XI0/XI48/XI11/MM6_d
+ N_XI0/XI48/XI11/NET36_XI0/XI48/XI11/MM6_g N_VSS_XI0/XI48/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM7 N_XI0/XI48/XI11/NET36_XI0/XI48/XI11/MM7_d
+ N_XI0/XI48/XI11/NET35_XI0/XI48/XI11/MM7_g N_VSS_XI0/XI48/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM8 N_XI0/XI48/XI11/NET35_XI0/XI48/XI11/MM8_d
+ N_WL<93>_XI0/XI48/XI11/MM8_g N_BLN<4>_XI0/XI48/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI11/MM5 N_XI0/XI48/XI11/NET34_XI0/XI48/XI11/MM5_d
+ N_XI0/XI48/XI11/NET33_XI0/XI48/XI11/MM5_g N_VDD_XI0/XI48/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI11/MM4 N_XI0/XI48/XI11/NET33_XI0/XI48/XI11/MM4_d
+ N_XI0/XI48/XI11/NET34_XI0/XI48/XI11/MM4_g N_VDD_XI0/XI48/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI11/MM10 N_XI0/XI48/XI11/NET35_XI0/XI48/XI11/MM10_d
+ N_XI0/XI48/XI11/NET36_XI0/XI48/XI11/MM10_g N_VDD_XI0/XI48/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI11/MM11 N_XI0/XI48/XI11/NET36_XI0/XI48/XI11/MM11_d
+ N_XI0/XI48/XI11/NET35_XI0/XI48/XI11/MM11_g N_VDD_XI0/XI48/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI12/MM2 N_XI0/XI48/XI12/NET34_XI0/XI48/XI12/MM2_d
+ N_XI0/XI48/XI12/NET33_XI0/XI48/XI12/MM2_g N_VSS_XI0/XI48/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM3 N_XI0/XI48/XI12/NET33_XI0/XI48/XI12/MM3_d
+ N_WL<92>_XI0/XI48/XI12/MM3_g N_BLN<3>_XI0/XI48/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM0 N_XI0/XI48/XI12/NET34_XI0/XI48/XI12/MM0_d
+ N_WL<92>_XI0/XI48/XI12/MM0_g N_BL<3>_XI0/XI48/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM1 N_XI0/XI48/XI12/NET33_XI0/XI48/XI12/MM1_d
+ N_XI0/XI48/XI12/NET34_XI0/XI48/XI12/MM1_g N_VSS_XI0/XI48/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM9 N_XI0/XI48/XI12/NET36_XI0/XI48/XI12/MM9_d
+ N_WL<93>_XI0/XI48/XI12/MM9_g N_BL<3>_XI0/XI48/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM6 N_XI0/XI48/XI12/NET35_XI0/XI48/XI12/MM6_d
+ N_XI0/XI48/XI12/NET36_XI0/XI48/XI12/MM6_g N_VSS_XI0/XI48/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM7 N_XI0/XI48/XI12/NET36_XI0/XI48/XI12/MM7_d
+ N_XI0/XI48/XI12/NET35_XI0/XI48/XI12/MM7_g N_VSS_XI0/XI48/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM8 N_XI0/XI48/XI12/NET35_XI0/XI48/XI12/MM8_d
+ N_WL<93>_XI0/XI48/XI12/MM8_g N_BLN<3>_XI0/XI48/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI12/MM5 N_XI0/XI48/XI12/NET34_XI0/XI48/XI12/MM5_d
+ N_XI0/XI48/XI12/NET33_XI0/XI48/XI12/MM5_g N_VDD_XI0/XI48/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI12/MM4 N_XI0/XI48/XI12/NET33_XI0/XI48/XI12/MM4_d
+ N_XI0/XI48/XI12/NET34_XI0/XI48/XI12/MM4_g N_VDD_XI0/XI48/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI12/MM10 N_XI0/XI48/XI12/NET35_XI0/XI48/XI12/MM10_d
+ N_XI0/XI48/XI12/NET36_XI0/XI48/XI12/MM10_g N_VDD_XI0/XI48/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI12/MM11 N_XI0/XI48/XI12/NET36_XI0/XI48/XI12/MM11_d
+ N_XI0/XI48/XI12/NET35_XI0/XI48/XI12/MM11_g N_VDD_XI0/XI48/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI13/MM2 N_XI0/XI48/XI13/NET34_XI0/XI48/XI13/MM2_d
+ N_XI0/XI48/XI13/NET33_XI0/XI48/XI13/MM2_g N_VSS_XI0/XI48/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM3 N_XI0/XI48/XI13/NET33_XI0/XI48/XI13/MM3_d
+ N_WL<92>_XI0/XI48/XI13/MM3_g N_BLN<2>_XI0/XI48/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM0 N_XI0/XI48/XI13/NET34_XI0/XI48/XI13/MM0_d
+ N_WL<92>_XI0/XI48/XI13/MM0_g N_BL<2>_XI0/XI48/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM1 N_XI0/XI48/XI13/NET33_XI0/XI48/XI13/MM1_d
+ N_XI0/XI48/XI13/NET34_XI0/XI48/XI13/MM1_g N_VSS_XI0/XI48/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM9 N_XI0/XI48/XI13/NET36_XI0/XI48/XI13/MM9_d
+ N_WL<93>_XI0/XI48/XI13/MM9_g N_BL<2>_XI0/XI48/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM6 N_XI0/XI48/XI13/NET35_XI0/XI48/XI13/MM6_d
+ N_XI0/XI48/XI13/NET36_XI0/XI48/XI13/MM6_g N_VSS_XI0/XI48/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM7 N_XI0/XI48/XI13/NET36_XI0/XI48/XI13/MM7_d
+ N_XI0/XI48/XI13/NET35_XI0/XI48/XI13/MM7_g N_VSS_XI0/XI48/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM8 N_XI0/XI48/XI13/NET35_XI0/XI48/XI13/MM8_d
+ N_WL<93>_XI0/XI48/XI13/MM8_g N_BLN<2>_XI0/XI48/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI13/MM5 N_XI0/XI48/XI13/NET34_XI0/XI48/XI13/MM5_d
+ N_XI0/XI48/XI13/NET33_XI0/XI48/XI13/MM5_g N_VDD_XI0/XI48/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI13/MM4 N_XI0/XI48/XI13/NET33_XI0/XI48/XI13/MM4_d
+ N_XI0/XI48/XI13/NET34_XI0/XI48/XI13/MM4_g N_VDD_XI0/XI48/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI13/MM10 N_XI0/XI48/XI13/NET35_XI0/XI48/XI13/MM10_d
+ N_XI0/XI48/XI13/NET36_XI0/XI48/XI13/MM10_g N_VDD_XI0/XI48/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI13/MM11 N_XI0/XI48/XI13/NET36_XI0/XI48/XI13/MM11_d
+ N_XI0/XI48/XI13/NET35_XI0/XI48/XI13/MM11_g N_VDD_XI0/XI48/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI14/MM2 N_XI0/XI48/XI14/NET34_XI0/XI48/XI14/MM2_d
+ N_XI0/XI48/XI14/NET33_XI0/XI48/XI14/MM2_g N_VSS_XI0/XI48/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM3 N_XI0/XI48/XI14/NET33_XI0/XI48/XI14/MM3_d
+ N_WL<92>_XI0/XI48/XI14/MM3_g N_BLN<1>_XI0/XI48/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM0 N_XI0/XI48/XI14/NET34_XI0/XI48/XI14/MM0_d
+ N_WL<92>_XI0/XI48/XI14/MM0_g N_BL<1>_XI0/XI48/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM1 N_XI0/XI48/XI14/NET33_XI0/XI48/XI14/MM1_d
+ N_XI0/XI48/XI14/NET34_XI0/XI48/XI14/MM1_g N_VSS_XI0/XI48/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM9 N_XI0/XI48/XI14/NET36_XI0/XI48/XI14/MM9_d
+ N_WL<93>_XI0/XI48/XI14/MM9_g N_BL<1>_XI0/XI48/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM6 N_XI0/XI48/XI14/NET35_XI0/XI48/XI14/MM6_d
+ N_XI0/XI48/XI14/NET36_XI0/XI48/XI14/MM6_g N_VSS_XI0/XI48/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM7 N_XI0/XI48/XI14/NET36_XI0/XI48/XI14/MM7_d
+ N_XI0/XI48/XI14/NET35_XI0/XI48/XI14/MM7_g N_VSS_XI0/XI48/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM8 N_XI0/XI48/XI14/NET35_XI0/XI48/XI14/MM8_d
+ N_WL<93>_XI0/XI48/XI14/MM8_g N_BLN<1>_XI0/XI48/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI14/MM5 N_XI0/XI48/XI14/NET34_XI0/XI48/XI14/MM5_d
+ N_XI0/XI48/XI14/NET33_XI0/XI48/XI14/MM5_g N_VDD_XI0/XI48/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI14/MM4 N_XI0/XI48/XI14/NET33_XI0/XI48/XI14/MM4_d
+ N_XI0/XI48/XI14/NET34_XI0/XI48/XI14/MM4_g N_VDD_XI0/XI48/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI14/MM10 N_XI0/XI48/XI14/NET35_XI0/XI48/XI14/MM10_d
+ N_XI0/XI48/XI14/NET36_XI0/XI48/XI14/MM10_g N_VDD_XI0/XI48/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI14/MM11 N_XI0/XI48/XI14/NET36_XI0/XI48/XI14/MM11_d
+ N_XI0/XI48/XI14/NET35_XI0/XI48/XI14/MM11_g N_VDD_XI0/XI48/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI15/MM2 N_XI0/XI48/XI15/NET34_XI0/XI48/XI15/MM2_d
+ N_XI0/XI48/XI15/NET33_XI0/XI48/XI15/MM2_g N_VSS_XI0/XI48/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM3 N_XI0/XI48/XI15/NET33_XI0/XI48/XI15/MM3_d
+ N_WL<92>_XI0/XI48/XI15/MM3_g N_BLN<0>_XI0/XI48/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM0 N_XI0/XI48/XI15/NET34_XI0/XI48/XI15/MM0_d
+ N_WL<92>_XI0/XI48/XI15/MM0_g N_BL<0>_XI0/XI48/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM1 N_XI0/XI48/XI15/NET33_XI0/XI48/XI15/MM1_d
+ N_XI0/XI48/XI15/NET34_XI0/XI48/XI15/MM1_g N_VSS_XI0/XI48/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM9 N_XI0/XI48/XI15/NET36_XI0/XI48/XI15/MM9_d
+ N_WL<93>_XI0/XI48/XI15/MM9_g N_BL<0>_XI0/XI48/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM6 N_XI0/XI48/XI15/NET35_XI0/XI48/XI15/MM6_d
+ N_XI0/XI48/XI15/NET36_XI0/XI48/XI15/MM6_g N_VSS_XI0/XI48/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM7 N_XI0/XI48/XI15/NET36_XI0/XI48/XI15/MM7_d
+ N_XI0/XI48/XI15/NET35_XI0/XI48/XI15/MM7_g N_VSS_XI0/XI48/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM8 N_XI0/XI48/XI15/NET35_XI0/XI48/XI15/MM8_d
+ N_WL<93>_XI0/XI48/XI15/MM8_g N_BLN<0>_XI0/XI48/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI48/XI15/MM5 N_XI0/XI48/XI15/NET34_XI0/XI48/XI15/MM5_d
+ N_XI0/XI48/XI15/NET33_XI0/XI48/XI15/MM5_g N_VDD_XI0/XI48/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI15/MM4 N_XI0/XI48/XI15/NET33_XI0/XI48/XI15/MM4_d
+ N_XI0/XI48/XI15/NET34_XI0/XI48/XI15/MM4_g N_VDD_XI0/XI48/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI15/MM10 N_XI0/XI48/XI15/NET35_XI0/XI48/XI15/MM10_d
+ N_XI0/XI48/XI15/NET36_XI0/XI48/XI15/MM10_g N_VDD_XI0/XI48/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI48/XI15/MM11 N_XI0/XI48/XI15/NET36_XI0/XI48/XI15/MM11_d
+ N_XI0/XI48/XI15/NET35_XI0/XI48/XI15/MM11_g N_VDD_XI0/XI48/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI0/MM2 N_XI0/XI49/XI0/NET34_XI0/XI49/XI0/MM2_d
+ N_XI0/XI49/XI0/NET33_XI0/XI49/XI0/MM2_g N_VSS_XI0/XI49/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM3 N_XI0/XI49/XI0/NET33_XI0/XI49/XI0/MM3_d
+ N_WL<94>_XI0/XI49/XI0/MM3_g N_BLN<15>_XI0/XI49/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM0 N_XI0/XI49/XI0/NET34_XI0/XI49/XI0/MM0_d
+ N_WL<94>_XI0/XI49/XI0/MM0_g N_BL<15>_XI0/XI49/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM1 N_XI0/XI49/XI0/NET33_XI0/XI49/XI0/MM1_d
+ N_XI0/XI49/XI0/NET34_XI0/XI49/XI0/MM1_g N_VSS_XI0/XI49/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM9 N_XI0/XI49/XI0/NET36_XI0/XI49/XI0/MM9_d
+ N_WL<95>_XI0/XI49/XI0/MM9_g N_BL<15>_XI0/XI49/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM6 N_XI0/XI49/XI0/NET35_XI0/XI49/XI0/MM6_d
+ N_XI0/XI49/XI0/NET36_XI0/XI49/XI0/MM6_g N_VSS_XI0/XI49/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM7 N_XI0/XI49/XI0/NET36_XI0/XI49/XI0/MM7_d
+ N_XI0/XI49/XI0/NET35_XI0/XI49/XI0/MM7_g N_VSS_XI0/XI49/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM8 N_XI0/XI49/XI0/NET35_XI0/XI49/XI0/MM8_d
+ N_WL<95>_XI0/XI49/XI0/MM8_g N_BLN<15>_XI0/XI49/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI0/MM5 N_XI0/XI49/XI0/NET34_XI0/XI49/XI0/MM5_d
+ N_XI0/XI49/XI0/NET33_XI0/XI49/XI0/MM5_g N_VDD_XI0/XI49/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI0/MM4 N_XI0/XI49/XI0/NET33_XI0/XI49/XI0/MM4_d
+ N_XI0/XI49/XI0/NET34_XI0/XI49/XI0/MM4_g N_VDD_XI0/XI49/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI0/MM10 N_XI0/XI49/XI0/NET35_XI0/XI49/XI0/MM10_d
+ N_XI0/XI49/XI0/NET36_XI0/XI49/XI0/MM10_g N_VDD_XI0/XI49/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI0/MM11 N_XI0/XI49/XI0/NET36_XI0/XI49/XI0/MM11_d
+ N_XI0/XI49/XI0/NET35_XI0/XI49/XI0/MM11_g N_VDD_XI0/XI49/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI1/MM2 N_XI0/XI49/XI1/NET34_XI0/XI49/XI1/MM2_d
+ N_XI0/XI49/XI1/NET33_XI0/XI49/XI1/MM2_g N_VSS_XI0/XI49/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM3 N_XI0/XI49/XI1/NET33_XI0/XI49/XI1/MM3_d
+ N_WL<94>_XI0/XI49/XI1/MM3_g N_BLN<14>_XI0/XI49/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM0 N_XI0/XI49/XI1/NET34_XI0/XI49/XI1/MM0_d
+ N_WL<94>_XI0/XI49/XI1/MM0_g N_BL<14>_XI0/XI49/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM1 N_XI0/XI49/XI1/NET33_XI0/XI49/XI1/MM1_d
+ N_XI0/XI49/XI1/NET34_XI0/XI49/XI1/MM1_g N_VSS_XI0/XI49/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM9 N_XI0/XI49/XI1/NET36_XI0/XI49/XI1/MM9_d
+ N_WL<95>_XI0/XI49/XI1/MM9_g N_BL<14>_XI0/XI49/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM6 N_XI0/XI49/XI1/NET35_XI0/XI49/XI1/MM6_d
+ N_XI0/XI49/XI1/NET36_XI0/XI49/XI1/MM6_g N_VSS_XI0/XI49/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM7 N_XI0/XI49/XI1/NET36_XI0/XI49/XI1/MM7_d
+ N_XI0/XI49/XI1/NET35_XI0/XI49/XI1/MM7_g N_VSS_XI0/XI49/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM8 N_XI0/XI49/XI1/NET35_XI0/XI49/XI1/MM8_d
+ N_WL<95>_XI0/XI49/XI1/MM8_g N_BLN<14>_XI0/XI49/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI1/MM5 N_XI0/XI49/XI1/NET34_XI0/XI49/XI1/MM5_d
+ N_XI0/XI49/XI1/NET33_XI0/XI49/XI1/MM5_g N_VDD_XI0/XI49/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI1/MM4 N_XI0/XI49/XI1/NET33_XI0/XI49/XI1/MM4_d
+ N_XI0/XI49/XI1/NET34_XI0/XI49/XI1/MM4_g N_VDD_XI0/XI49/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI1/MM10 N_XI0/XI49/XI1/NET35_XI0/XI49/XI1/MM10_d
+ N_XI0/XI49/XI1/NET36_XI0/XI49/XI1/MM10_g N_VDD_XI0/XI49/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI1/MM11 N_XI0/XI49/XI1/NET36_XI0/XI49/XI1/MM11_d
+ N_XI0/XI49/XI1/NET35_XI0/XI49/XI1/MM11_g N_VDD_XI0/XI49/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI2/MM2 N_XI0/XI49/XI2/NET34_XI0/XI49/XI2/MM2_d
+ N_XI0/XI49/XI2/NET33_XI0/XI49/XI2/MM2_g N_VSS_XI0/XI49/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM3 N_XI0/XI49/XI2/NET33_XI0/XI49/XI2/MM3_d
+ N_WL<94>_XI0/XI49/XI2/MM3_g N_BLN<13>_XI0/XI49/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM0 N_XI0/XI49/XI2/NET34_XI0/XI49/XI2/MM0_d
+ N_WL<94>_XI0/XI49/XI2/MM0_g N_BL<13>_XI0/XI49/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM1 N_XI0/XI49/XI2/NET33_XI0/XI49/XI2/MM1_d
+ N_XI0/XI49/XI2/NET34_XI0/XI49/XI2/MM1_g N_VSS_XI0/XI49/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM9 N_XI0/XI49/XI2/NET36_XI0/XI49/XI2/MM9_d
+ N_WL<95>_XI0/XI49/XI2/MM9_g N_BL<13>_XI0/XI49/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM6 N_XI0/XI49/XI2/NET35_XI0/XI49/XI2/MM6_d
+ N_XI0/XI49/XI2/NET36_XI0/XI49/XI2/MM6_g N_VSS_XI0/XI49/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM7 N_XI0/XI49/XI2/NET36_XI0/XI49/XI2/MM7_d
+ N_XI0/XI49/XI2/NET35_XI0/XI49/XI2/MM7_g N_VSS_XI0/XI49/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM8 N_XI0/XI49/XI2/NET35_XI0/XI49/XI2/MM8_d
+ N_WL<95>_XI0/XI49/XI2/MM8_g N_BLN<13>_XI0/XI49/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI2/MM5 N_XI0/XI49/XI2/NET34_XI0/XI49/XI2/MM5_d
+ N_XI0/XI49/XI2/NET33_XI0/XI49/XI2/MM5_g N_VDD_XI0/XI49/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI2/MM4 N_XI0/XI49/XI2/NET33_XI0/XI49/XI2/MM4_d
+ N_XI0/XI49/XI2/NET34_XI0/XI49/XI2/MM4_g N_VDD_XI0/XI49/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI2/MM10 N_XI0/XI49/XI2/NET35_XI0/XI49/XI2/MM10_d
+ N_XI0/XI49/XI2/NET36_XI0/XI49/XI2/MM10_g N_VDD_XI0/XI49/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI2/MM11 N_XI0/XI49/XI2/NET36_XI0/XI49/XI2/MM11_d
+ N_XI0/XI49/XI2/NET35_XI0/XI49/XI2/MM11_g N_VDD_XI0/XI49/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI3/MM2 N_XI0/XI49/XI3/NET34_XI0/XI49/XI3/MM2_d
+ N_XI0/XI49/XI3/NET33_XI0/XI49/XI3/MM2_g N_VSS_XI0/XI49/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM3 N_XI0/XI49/XI3/NET33_XI0/XI49/XI3/MM3_d
+ N_WL<94>_XI0/XI49/XI3/MM3_g N_BLN<12>_XI0/XI49/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM0 N_XI0/XI49/XI3/NET34_XI0/XI49/XI3/MM0_d
+ N_WL<94>_XI0/XI49/XI3/MM0_g N_BL<12>_XI0/XI49/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM1 N_XI0/XI49/XI3/NET33_XI0/XI49/XI3/MM1_d
+ N_XI0/XI49/XI3/NET34_XI0/XI49/XI3/MM1_g N_VSS_XI0/XI49/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM9 N_XI0/XI49/XI3/NET36_XI0/XI49/XI3/MM9_d
+ N_WL<95>_XI0/XI49/XI3/MM9_g N_BL<12>_XI0/XI49/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM6 N_XI0/XI49/XI3/NET35_XI0/XI49/XI3/MM6_d
+ N_XI0/XI49/XI3/NET36_XI0/XI49/XI3/MM6_g N_VSS_XI0/XI49/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM7 N_XI0/XI49/XI3/NET36_XI0/XI49/XI3/MM7_d
+ N_XI0/XI49/XI3/NET35_XI0/XI49/XI3/MM7_g N_VSS_XI0/XI49/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM8 N_XI0/XI49/XI3/NET35_XI0/XI49/XI3/MM8_d
+ N_WL<95>_XI0/XI49/XI3/MM8_g N_BLN<12>_XI0/XI49/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI3/MM5 N_XI0/XI49/XI3/NET34_XI0/XI49/XI3/MM5_d
+ N_XI0/XI49/XI3/NET33_XI0/XI49/XI3/MM5_g N_VDD_XI0/XI49/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI3/MM4 N_XI0/XI49/XI3/NET33_XI0/XI49/XI3/MM4_d
+ N_XI0/XI49/XI3/NET34_XI0/XI49/XI3/MM4_g N_VDD_XI0/XI49/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI3/MM10 N_XI0/XI49/XI3/NET35_XI0/XI49/XI3/MM10_d
+ N_XI0/XI49/XI3/NET36_XI0/XI49/XI3/MM10_g N_VDD_XI0/XI49/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI3/MM11 N_XI0/XI49/XI3/NET36_XI0/XI49/XI3/MM11_d
+ N_XI0/XI49/XI3/NET35_XI0/XI49/XI3/MM11_g N_VDD_XI0/XI49/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI4/MM2 N_XI0/XI49/XI4/NET34_XI0/XI49/XI4/MM2_d
+ N_XI0/XI49/XI4/NET33_XI0/XI49/XI4/MM2_g N_VSS_XI0/XI49/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM3 N_XI0/XI49/XI4/NET33_XI0/XI49/XI4/MM3_d
+ N_WL<94>_XI0/XI49/XI4/MM3_g N_BLN<11>_XI0/XI49/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM0 N_XI0/XI49/XI4/NET34_XI0/XI49/XI4/MM0_d
+ N_WL<94>_XI0/XI49/XI4/MM0_g N_BL<11>_XI0/XI49/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM1 N_XI0/XI49/XI4/NET33_XI0/XI49/XI4/MM1_d
+ N_XI0/XI49/XI4/NET34_XI0/XI49/XI4/MM1_g N_VSS_XI0/XI49/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM9 N_XI0/XI49/XI4/NET36_XI0/XI49/XI4/MM9_d
+ N_WL<95>_XI0/XI49/XI4/MM9_g N_BL<11>_XI0/XI49/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM6 N_XI0/XI49/XI4/NET35_XI0/XI49/XI4/MM6_d
+ N_XI0/XI49/XI4/NET36_XI0/XI49/XI4/MM6_g N_VSS_XI0/XI49/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM7 N_XI0/XI49/XI4/NET36_XI0/XI49/XI4/MM7_d
+ N_XI0/XI49/XI4/NET35_XI0/XI49/XI4/MM7_g N_VSS_XI0/XI49/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM8 N_XI0/XI49/XI4/NET35_XI0/XI49/XI4/MM8_d
+ N_WL<95>_XI0/XI49/XI4/MM8_g N_BLN<11>_XI0/XI49/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI4/MM5 N_XI0/XI49/XI4/NET34_XI0/XI49/XI4/MM5_d
+ N_XI0/XI49/XI4/NET33_XI0/XI49/XI4/MM5_g N_VDD_XI0/XI49/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI4/MM4 N_XI0/XI49/XI4/NET33_XI0/XI49/XI4/MM4_d
+ N_XI0/XI49/XI4/NET34_XI0/XI49/XI4/MM4_g N_VDD_XI0/XI49/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI4/MM10 N_XI0/XI49/XI4/NET35_XI0/XI49/XI4/MM10_d
+ N_XI0/XI49/XI4/NET36_XI0/XI49/XI4/MM10_g N_VDD_XI0/XI49/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI4/MM11 N_XI0/XI49/XI4/NET36_XI0/XI49/XI4/MM11_d
+ N_XI0/XI49/XI4/NET35_XI0/XI49/XI4/MM11_g N_VDD_XI0/XI49/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI5/MM2 N_XI0/XI49/XI5/NET34_XI0/XI49/XI5/MM2_d
+ N_XI0/XI49/XI5/NET33_XI0/XI49/XI5/MM2_g N_VSS_XI0/XI49/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM3 N_XI0/XI49/XI5/NET33_XI0/XI49/XI5/MM3_d
+ N_WL<94>_XI0/XI49/XI5/MM3_g N_BLN<10>_XI0/XI49/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM0 N_XI0/XI49/XI5/NET34_XI0/XI49/XI5/MM0_d
+ N_WL<94>_XI0/XI49/XI5/MM0_g N_BL<10>_XI0/XI49/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM1 N_XI0/XI49/XI5/NET33_XI0/XI49/XI5/MM1_d
+ N_XI0/XI49/XI5/NET34_XI0/XI49/XI5/MM1_g N_VSS_XI0/XI49/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM9 N_XI0/XI49/XI5/NET36_XI0/XI49/XI5/MM9_d
+ N_WL<95>_XI0/XI49/XI5/MM9_g N_BL<10>_XI0/XI49/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM6 N_XI0/XI49/XI5/NET35_XI0/XI49/XI5/MM6_d
+ N_XI0/XI49/XI5/NET36_XI0/XI49/XI5/MM6_g N_VSS_XI0/XI49/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM7 N_XI0/XI49/XI5/NET36_XI0/XI49/XI5/MM7_d
+ N_XI0/XI49/XI5/NET35_XI0/XI49/XI5/MM7_g N_VSS_XI0/XI49/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM8 N_XI0/XI49/XI5/NET35_XI0/XI49/XI5/MM8_d
+ N_WL<95>_XI0/XI49/XI5/MM8_g N_BLN<10>_XI0/XI49/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI5/MM5 N_XI0/XI49/XI5/NET34_XI0/XI49/XI5/MM5_d
+ N_XI0/XI49/XI5/NET33_XI0/XI49/XI5/MM5_g N_VDD_XI0/XI49/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI5/MM4 N_XI0/XI49/XI5/NET33_XI0/XI49/XI5/MM4_d
+ N_XI0/XI49/XI5/NET34_XI0/XI49/XI5/MM4_g N_VDD_XI0/XI49/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI5/MM10 N_XI0/XI49/XI5/NET35_XI0/XI49/XI5/MM10_d
+ N_XI0/XI49/XI5/NET36_XI0/XI49/XI5/MM10_g N_VDD_XI0/XI49/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI5/MM11 N_XI0/XI49/XI5/NET36_XI0/XI49/XI5/MM11_d
+ N_XI0/XI49/XI5/NET35_XI0/XI49/XI5/MM11_g N_VDD_XI0/XI49/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI6/MM2 N_XI0/XI49/XI6/NET34_XI0/XI49/XI6/MM2_d
+ N_XI0/XI49/XI6/NET33_XI0/XI49/XI6/MM2_g N_VSS_XI0/XI49/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM3 N_XI0/XI49/XI6/NET33_XI0/XI49/XI6/MM3_d
+ N_WL<94>_XI0/XI49/XI6/MM3_g N_BLN<9>_XI0/XI49/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM0 N_XI0/XI49/XI6/NET34_XI0/XI49/XI6/MM0_d
+ N_WL<94>_XI0/XI49/XI6/MM0_g N_BL<9>_XI0/XI49/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM1 N_XI0/XI49/XI6/NET33_XI0/XI49/XI6/MM1_d
+ N_XI0/XI49/XI6/NET34_XI0/XI49/XI6/MM1_g N_VSS_XI0/XI49/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM9 N_XI0/XI49/XI6/NET36_XI0/XI49/XI6/MM9_d
+ N_WL<95>_XI0/XI49/XI6/MM9_g N_BL<9>_XI0/XI49/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM6 N_XI0/XI49/XI6/NET35_XI0/XI49/XI6/MM6_d
+ N_XI0/XI49/XI6/NET36_XI0/XI49/XI6/MM6_g N_VSS_XI0/XI49/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM7 N_XI0/XI49/XI6/NET36_XI0/XI49/XI6/MM7_d
+ N_XI0/XI49/XI6/NET35_XI0/XI49/XI6/MM7_g N_VSS_XI0/XI49/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM8 N_XI0/XI49/XI6/NET35_XI0/XI49/XI6/MM8_d
+ N_WL<95>_XI0/XI49/XI6/MM8_g N_BLN<9>_XI0/XI49/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI6/MM5 N_XI0/XI49/XI6/NET34_XI0/XI49/XI6/MM5_d
+ N_XI0/XI49/XI6/NET33_XI0/XI49/XI6/MM5_g N_VDD_XI0/XI49/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI6/MM4 N_XI0/XI49/XI6/NET33_XI0/XI49/XI6/MM4_d
+ N_XI0/XI49/XI6/NET34_XI0/XI49/XI6/MM4_g N_VDD_XI0/XI49/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI6/MM10 N_XI0/XI49/XI6/NET35_XI0/XI49/XI6/MM10_d
+ N_XI0/XI49/XI6/NET36_XI0/XI49/XI6/MM10_g N_VDD_XI0/XI49/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI6/MM11 N_XI0/XI49/XI6/NET36_XI0/XI49/XI6/MM11_d
+ N_XI0/XI49/XI6/NET35_XI0/XI49/XI6/MM11_g N_VDD_XI0/XI49/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI7/MM2 N_XI0/XI49/XI7/NET34_XI0/XI49/XI7/MM2_d
+ N_XI0/XI49/XI7/NET33_XI0/XI49/XI7/MM2_g N_VSS_XI0/XI49/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM3 N_XI0/XI49/XI7/NET33_XI0/XI49/XI7/MM3_d
+ N_WL<94>_XI0/XI49/XI7/MM3_g N_BLN<8>_XI0/XI49/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM0 N_XI0/XI49/XI7/NET34_XI0/XI49/XI7/MM0_d
+ N_WL<94>_XI0/XI49/XI7/MM0_g N_BL<8>_XI0/XI49/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM1 N_XI0/XI49/XI7/NET33_XI0/XI49/XI7/MM1_d
+ N_XI0/XI49/XI7/NET34_XI0/XI49/XI7/MM1_g N_VSS_XI0/XI49/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM9 N_XI0/XI49/XI7/NET36_XI0/XI49/XI7/MM9_d
+ N_WL<95>_XI0/XI49/XI7/MM9_g N_BL<8>_XI0/XI49/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM6 N_XI0/XI49/XI7/NET35_XI0/XI49/XI7/MM6_d
+ N_XI0/XI49/XI7/NET36_XI0/XI49/XI7/MM6_g N_VSS_XI0/XI49/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM7 N_XI0/XI49/XI7/NET36_XI0/XI49/XI7/MM7_d
+ N_XI0/XI49/XI7/NET35_XI0/XI49/XI7/MM7_g N_VSS_XI0/XI49/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM8 N_XI0/XI49/XI7/NET35_XI0/XI49/XI7/MM8_d
+ N_WL<95>_XI0/XI49/XI7/MM8_g N_BLN<8>_XI0/XI49/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI7/MM5 N_XI0/XI49/XI7/NET34_XI0/XI49/XI7/MM5_d
+ N_XI0/XI49/XI7/NET33_XI0/XI49/XI7/MM5_g N_VDD_XI0/XI49/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI7/MM4 N_XI0/XI49/XI7/NET33_XI0/XI49/XI7/MM4_d
+ N_XI0/XI49/XI7/NET34_XI0/XI49/XI7/MM4_g N_VDD_XI0/XI49/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI7/MM10 N_XI0/XI49/XI7/NET35_XI0/XI49/XI7/MM10_d
+ N_XI0/XI49/XI7/NET36_XI0/XI49/XI7/MM10_g N_VDD_XI0/XI49/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI7/MM11 N_XI0/XI49/XI7/NET36_XI0/XI49/XI7/MM11_d
+ N_XI0/XI49/XI7/NET35_XI0/XI49/XI7/MM11_g N_VDD_XI0/XI49/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI8/MM2 N_XI0/XI49/XI8/NET34_XI0/XI49/XI8/MM2_d
+ N_XI0/XI49/XI8/NET33_XI0/XI49/XI8/MM2_g N_VSS_XI0/XI49/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM3 N_XI0/XI49/XI8/NET33_XI0/XI49/XI8/MM3_d
+ N_WL<94>_XI0/XI49/XI8/MM3_g N_BLN<7>_XI0/XI49/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM0 N_XI0/XI49/XI8/NET34_XI0/XI49/XI8/MM0_d
+ N_WL<94>_XI0/XI49/XI8/MM0_g N_BL<7>_XI0/XI49/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM1 N_XI0/XI49/XI8/NET33_XI0/XI49/XI8/MM1_d
+ N_XI0/XI49/XI8/NET34_XI0/XI49/XI8/MM1_g N_VSS_XI0/XI49/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM9 N_XI0/XI49/XI8/NET36_XI0/XI49/XI8/MM9_d
+ N_WL<95>_XI0/XI49/XI8/MM9_g N_BL<7>_XI0/XI49/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM6 N_XI0/XI49/XI8/NET35_XI0/XI49/XI8/MM6_d
+ N_XI0/XI49/XI8/NET36_XI0/XI49/XI8/MM6_g N_VSS_XI0/XI49/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM7 N_XI0/XI49/XI8/NET36_XI0/XI49/XI8/MM7_d
+ N_XI0/XI49/XI8/NET35_XI0/XI49/XI8/MM7_g N_VSS_XI0/XI49/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM8 N_XI0/XI49/XI8/NET35_XI0/XI49/XI8/MM8_d
+ N_WL<95>_XI0/XI49/XI8/MM8_g N_BLN<7>_XI0/XI49/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI8/MM5 N_XI0/XI49/XI8/NET34_XI0/XI49/XI8/MM5_d
+ N_XI0/XI49/XI8/NET33_XI0/XI49/XI8/MM5_g N_VDD_XI0/XI49/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI8/MM4 N_XI0/XI49/XI8/NET33_XI0/XI49/XI8/MM4_d
+ N_XI0/XI49/XI8/NET34_XI0/XI49/XI8/MM4_g N_VDD_XI0/XI49/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI8/MM10 N_XI0/XI49/XI8/NET35_XI0/XI49/XI8/MM10_d
+ N_XI0/XI49/XI8/NET36_XI0/XI49/XI8/MM10_g N_VDD_XI0/XI49/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI8/MM11 N_XI0/XI49/XI8/NET36_XI0/XI49/XI8/MM11_d
+ N_XI0/XI49/XI8/NET35_XI0/XI49/XI8/MM11_g N_VDD_XI0/XI49/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI9/MM2 N_XI0/XI49/XI9/NET34_XI0/XI49/XI9/MM2_d
+ N_XI0/XI49/XI9/NET33_XI0/XI49/XI9/MM2_g N_VSS_XI0/XI49/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM3 N_XI0/XI49/XI9/NET33_XI0/XI49/XI9/MM3_d
+ N_WL<94>_XI0/XI49/XI9/MM3_g N_BLN<6>_XI0/XI49/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM0 N_XI0/XI49/XI9/NET34_XI0/XI49/XI9/MM0_d
+ N_WL<94>_XI0/XI49/XI9/MM0_g N_BL<6>_XI0/XI49/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM1 N_XI0/XI49/XI9/NET33_XI0/XI49/XI9/MM1_d
+ N_XI0/XI49/XI9/NET34_XI0/XI49/XI9/MM1_g N_VSS_XI0/XI49/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM9 N_XI0/XI49/XI9/NET36_XI0/XI49/XI9/MM9_d
+ N_WL<95>_XI0/XI49/XI9/MM9_g N_BL<6>_XI0/XI49/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM6 N_XI0/XI49/XI9/NET35_XI0/XI49/XI9/MM6_d
+ N_XI0/XI49/XI9/NET36_XI0/XI49/XI9/MM6_g N_VSS_XI0/XI49/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM7 N_XI0/XI49/XI9/NET36_XI0/XI49/XI9/MM7_d
+ N_XI0/XI49/XI9/NET35_XI0/XI49/XI9/MM7_g N_VSS_XI0/XI49/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM8 N_XI0/XI49/XI9/NET35_XI0/XI49/XI9/MM8_d
+ N_WL<95>_XI0/XI49/XI9/MM8_g N_BLN<6>_XI0/XI49/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI9/MM5 N_XI0/XI49/XI9/NET34_XI0/XI49/XI9/MM5_d
+ N_XI0/XI49/XI9/NET33_XI0/XI49/XI9/MM5_g N_VDD_XI0/XI49/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI9/MM4 N_XI0/XI49/XI9/NET33_XI0/XI49/XI9/MM4_d
+ N_XI0/XI49/XI9/NET34_XI0/XI49/XI9/MM4_g N_VDD_XI0/XI49/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI9/MM10 N_XI0/XI49/XI9/NET35_XI0/XI49/XI9/MM10_d
+ N_XI0/XI49/XI9/NET36_XI0/XI49/XI9/MM10_g N_VDD_XI0/XI49/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI9/MM11 N_XI0/XI49/XI9/NET36_XI0/XI49/XI9/MM11_d
+ N_XI0/XI49/XI9/NET35_XI0/XI49/XI9/MM11_g N_VDD_XI0/XI49/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI10/MM2 N_XI0/XI49/XI10/NET34_XI0/XI49/XI10/MM2_d
+ N_XI0/XI49/XI10/NET33_XI0/XI49/XI10/MM2_g N_VSS_XI0/XI49/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM3 N_XI0/XI49/XI10/NET33_XI0/XI49/XI10/MM3_d
+ N_WL<94>_XI0/XI49/XI10/MM3_g N_BLN<5>_XI0/XI49/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM0 N_XI0/XI49/XI10/NET34_XI0/XI49/XI10/MM0_d
+ N_WL<94>_XI0/XI49/XI10/MM0_g N_BL<5>_XI0/XI49/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM1 N_XI0/XI49/XI10/NET33_XI0/XI49/XI10/MM1_d
+ N_XI0/XI49/XI10/NET34_XI0/XI49/XI10/MM1_g N_VSS_XI0/XI49/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM9 N_XI0/XI49/XI10/NET36_XI0/XI49/XI10/MM9_d
+ N_WL<95>_XI0/XI49/XI10/MM9_g N_BL<5>_XI0/XI49/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM6 N_XI0/XI49/XI10/NET35_XI0/XI49/XI10/MM6_d
+ N_XI0/XI49/XI10/NET36_XI0/XI49/XI10/MM6_g N_VSS_XI0/XI49/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM7 N_XI0/XI49/XI10/NET36_XI0/XI49/XI10/MM7_d
+ N_XI0/XI49/XI10/NET35_XI0/XI49/XI10/MM7_g N_VSS_XI0/XI49/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM8 N_XI0/XI49/XI10/NET35_XI0/XI49/XI10/MM8_d
+ N_WL<95>_XI0/XI49/XI10/MM8_g N_BLN<5>_XI0/XI49/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI10/MM5 N_XI0/XI49/XI10/NET34_XI0/XI49/XI10/MM5_d
+ N_XI0/XI49/XI10/NET33_XI0/XI49/XI10/MM5_g N_VDD_XI0/XI49/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI10/MM4 N_XI0/XI49/XI10/NET33_XI0/XI49/XI10/MM4_d
+ N_XI0/XI49/XI10/NET34_XI0/XI49/XI10/MM4_g N_VDD_XI0/XI49/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI10/MM10 N_XI0/XI49/XI10/NET35_XI0/XI49/XI10/MM10_d
+ N_XI0/XI49/XI10/NET36_XI0/XI49/XI10/MM10_g N_VDD_XI0/XI49/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI10/MM11 N_XI0/XI49/XI10/NET36_XI0/XI49/XI10/MM11_d
+ N_XI0/XI49/XI10/NET35_XI0/XI49/XI10/MM11_g N_VDD_XI0/XI49/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI11/MM2 N_XI0/XI49/XI11/NET34_XI0/XI49/XI11/MM2_d
+ N_XI0/XI49/XI11/NET33_XI0/XI49/XI11/MM2_g N_VSS_XI0/XI49/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM3 N_XI0/XI49/XI11/NET33_XI0/XI49/XI11/MM3_d
+ N_WL<94>_XI0/XI49/XI11/MM3_g N_BLN<4>_XI0/XI49/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM0 N_XI0/XI49/XI11/NET34_XI0/XI49/XI11/MM0_d
+ N_WL<94>_XI0/XI49/XI11/MM0_g N_BL<4>_XI0/XI49/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM1 N_XI0/XI49/XI11/NET33_XI0/XI49/XI11/MM1_d
+ N_XI0/XI49/XI11/NET34_XI0/XI49/XI11/MM1_g N_VSS_XI0/XI49/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM9 N_XI0/XI49/XI11/NET36_XI0/XI49/XI11/MM9_d
+ N_WL<95>_XI0/XI49/XI11/MM9_g N_BL<4>_XI0/XI49/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM6 N_XI0/XI49/XI11/NET35_XI0/XI49/XI11/MM6_d
+ N_XI0/XI49/XI11/NET36_XI0/XI49/XI11/MM6_g N_VSS_XI0/XI49/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM7 N_XI0/XI49/XI11/NET36_XI0/XI49/XI11/MM7_d
+ N_XI0/XI49/XI11/NET35_XI0/XI49/XI11/MM7_g N_VSS_XI0/XI49/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM8 N_XI0/XI49/XI11/NET35_XI0/XI49/XI11/MM8_d
+ N_WL<95>_XI0/XI49/XI11/MM8_g N_BLN<4>_XI0/XI49/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI11/MM5 N_XI0/XI49/XI11/NET34_XI0/XI49/XI11/MM5_d
+ N_XI0/XI49/XI11/NET33_XI0/XI49/XI11/MM5_g N_VDD_XI0/XI49/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI11/MM4 N_XI0/XI49/XI11/NET33_XI0/XI49/XI11/MM4_d
+ N_XI0/XI49/XI11/NET34_XI0/XI49/XI11/MM4_g N_VDD_XI0/XI49/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI11/MM10 N_XI0/XI49/XI11/NET35_XI0/XI49/XI11/MM10_d
+ N_XI0/XI49/XI11/NET36_XI0/XI49/XI11/MM10_g N_VDD_XI0/XI49/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI11/MM11 N_XI0/XI49/XI11/NET36_XI0/XI49/XI11/MM11_d
+ N_XI0/XI49/XI11/NET35_XI0/XI49/XI11/MM11_g N_VDD_XI0/XI49/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI12/MM2 N_XI0/XI49/XI12/NET34_XI0/XI49/XI12/MM2_d
+ N_XI0/XI49/XI12/NET33_XI0/XI49/XI12/MM2_g N_VSS_XI0/XI49/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM3 N_XI0/XI49/XI12/NET33_XI0/XI49/XI12/MM3_d
+ N_WL<94>_XI0/XI49/XI12/MM3_g N_BLN<3>_XI0/XI49/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM0 N_XI0/XI49/XI12/NET34_XI0/XI49/XI12/MM0_d
+ N_WL<94>_XI0/XI49/XI12/MM0_g N_BL<3>_XI0/XI49/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM1 N_XI0/XI49/XI12/NET33_XI0/XI49/XI12/MM1_d
+ N_XI0/XI49/XI12/NET34_XI0/XI49/XI12/MM1_g N_VSS_XI0/XI49/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM9 N_XI0/XI49/XI12/NET36_XI0/XI49/XI12/MM9_d
+ N_WL<95>_XI0/XI49/XI12/MM9_g N_BL<3>_XI0/XI49/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM6 N_XI0/XI49/XI12/NET35_XI0/XI49/XI12/MM6_d
+ N_XI0/XI49/XI12/NET36_XI0/XI49/XI12/MM6_g N_VSS_XI0/XI49/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM7 N_XI0/XI49/XI12/NET36_XI0/XI49/XI12/MM7_d
+ N_XI0/XI49/XI12/NET35_XI0/XI49/XI12/MM7_g N_VSS_XI0/XI49/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM8 N_XI0/XI49/XI12/NET35_XI0/XI49/XI12/MM8_d
+ N_WL<95>_XI0/XI49/XI12/MM8_g N_BLN<3>_XI0/XI49/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI12/MM5 N_XI0/XI49/XI12/NET34_XI0/XI49/XI12/MM5_d
+ N_XI0/XI49/XI12/NET33_XI0/XI49/XI12/MM5_g N_VDD_XI0/XI49/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI12/MM4 N_XI0/XI49/XI12/NET33_XI0/XI49/XI12/MM4_d
+ N_XI0/XI49/XI12/NET34_XI0/XI49/XI12/MM4_g N_VDD_XI0/XI49/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI12/MM10 N_XI0/XI49/XI12/NET35_XI0/XI49/XI12/MM10_d
+ N_XI0/XI49/XI12/NET36_XI0/XI49/XI12/MM10_g N_VDD_XI0/XI49/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI12/MM11 N_XI0/XI49/XI12/NET36_XI0/XI49/XI12/MM11_d
+ N_XI0/XI49/XI12/NET35_XI0/XI49/XI12/MM11_g N_VDD_XI0/XI49/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI13/MM2 N_XI0/XI49/XI13/NET34_XI0/XI49/XI13/MM2_d
+ N_XI0/XI49/XI13/NET33_XI0/XI49/XI13/MM2_g N_VSS_XI0/XI49/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM3 N_XI0/XI49/XI13/NET33_XI0/XI49/XI13/MM3_d
+ N_WL<94>_XI0/XI49/XI13/MM3_g N_BLN<2>_XI0/XI49/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM0 N_XI0/XI49/XI13/NET34_XI0/XI49/XI13/MM0_d
+ N_WL<94>_XI0/XI49/XI13/MM0_g N_BL<2>_XI0/XI49/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM1 N_XI0/XI49/XI13/NET33_XI0/XI49/XI13/MM1_d
+ N_XI0/XI49/XI13/NET34_XI0/XI49/XI13/MM1_g N_VSS_XI0/XI49/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM9 N_XI0/XI49/XI13/NET36_XI0/XI49/XI13/MM9_d
+ N_WL<95>_XI0/XI49/XI13/MM9_g N_BL<2>_XI0/XI49/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM6 N_XI0/XI49/XI13/NET35_XI0/XI49/XI13/MM6_d
+ N_XI0/XI49/XI13/NET36_XI0/XI49/XI13/MM6_g N_VSS_XI0/XI49/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM7 N_XI0/XI49/XI13/NET36_XI0/XI49/XI13/MM7_d
+ N_XI0/XI49/XI13/NET35_XI0/XI49/XI13/MM7_g N_VSS_XI0/XI49/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM8 N_XI0/XI49/XI13/NET35_XI0/XI49/XI13/MM8_d
+ N_WL<95>_XI0/XI49/XI13/MM8_g N_BLN<2>_XI0/XI49/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI13/MM5 N_XI0/XI49/XI13/NET34_XI0/XI49/XI13/MM5_d
+ N_XI0/XI49/XI13/NET33_XI0/XI49/XI13/MM5_g N_VDD_XI0/XI49/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI13/MM4 N_XI0/XI49/XI13/NET33_XI0/XI49/XI13/MM4_d
+ N_XI0/XI49/XI13/NET34_XI0/XI49/XI13/MM4_g N_VDD_XI0/XI49/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI13/MM10 N_XI0/XI49/XI13/NET35_XI0/XI49/XI13/MM10_d
+ N_XI0/XI49/XI13/NET36_XI0/XI49/XI13/MM10_g N_VDD_XI0/XI49/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI13/MM11 N_XI0/XI49/XI13/NET36_XI0/XI49/XI13/MM11_d
+ N_XI0/XI49/XI13/NET35_XI0/XI49/XI13/MM11_g N_VDD_XI0/XI49/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI14/MM2 N_XI0/XI49/XI14/NET34_XI0/XI49/XI14/MM2_d
+ N_XI0/XI49/XI14/NET33_XI0/XI49/XI14/MM2_g N_VSS_XI0/XI49/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM3 N_XI0/XI49/XI14/NET33_XI0/XI49/XI14/MM3_d
+ N_WL<94>_XI0/XI49/XI14/MM3_g N_BLN<1>_XI0/XI49/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM0 N_XI0/XI49/XI14/NET34_XI0/XI49/XI14/MM0_d
+ N_WL<94>_XI0/XI49/XI14/MM0_g N_BL<1>_XI0/XI49/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM1 N_XI0/XI49/XI14/NET33_XI0/XI49/XI14/MM1_d
+ N_XI0/XI49/XI14/NET34_XI0/XI49/XI14/MM1_g N_VSS_XI0/XI49/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM9 N_XI0/XI49/XI14/NET36_XI0/XI49/XI14/MM9_d
+ N_WL<95>_XI0/XI49/XI14/MM9_g N_BL<1>_XI0/XI49/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM6 N_XI0/XI49/XI14/NET35_XI0/XI49/XI14/MM6_d
+ N_XI0/XI49/XI14/NET36_XI0/XI49/XI14/MM6_g N_VSS_XI0/XI49/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM7 N_XI0/XI49/XI14/NET36_XI0/XI49/XI14/MM7_d
+ N_XI0/XI49/XI14/NET35_XI0/XI49/XI14/MM7_g N_VSS_XI0/XI49/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM8 N_XI0/XI49/XI14/NET35_XI0/XI49/XI14/MM8_d
+ N_WL<95>_XI0/XI49/XI14/MM8_g N_BLN<1>_XI0/XI49/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI14/MM5 N_XI0/XI49/XI14/NET34_XI0/XI49/XI14/MM5_d
+ N_XI0/XI49/XI14/NET33_XI0/XI49/XI14/MM5_g N_VDD_XI0/XI49/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI14/MM4 N_XI0/XI49/XI14/NET33_XI0/XI49/XI14/MM4_d
+ N_XI0/XI49/XI14/NET34_XI0/XI49/XI14/MM4_g N_VDD_XI0/XI49/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI14/MM10 N_XI0/XI49/XI14/NET35_XI0/XI49/XI14/MM10_d
+ N_XI0/XI49/XI14/NET36_XI0/XI49/XI14/MM10_g N_VDD_XI0/XI49/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI14/MM11 N_XI0/XI49/XI14/NET36_XI0/XI49/XI14/MM11_d
+ N_XI0/XI49/XI14/NET35_XI0/XI49/XI14/MM11_g N_VDD_XI0/XI49/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI15/MM2 N_XI0/XI49/XI15/NET34_XI0/XI49/XI15/MM2_d
+ N_XI0/XI49/XI15/NET33_XI0/XI49/XI15/MM2_g N_VSS_XI0/XI49/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM3 N_XI0/XI49/XI15/NET33_XI0/XI49/XI15/MM3_d
+ N_WL<94>_XI0/XI49/XI15/MM3_g N_BLN<0>_XI0/XI49/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM0 N_XI0/XI49/XI15/NET34_XI0/XI49/XI15/MM0_d
+ N_WL<94>_XI0/XI49/XI15/MM0_g N_BL<0>_XI0/XI49/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM1 N_XI0/XI49/XI15/NET33_XI0/XI49/XI15/MM1_d
+ N_XI0/XI49/XI15/NET34_XI0/XI49/XI15/MM1_g N_VSS_XI0/XI49/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM9 N_XI0/XI49/XI15/NET36_XI0/XI49/XI15/MM9_d
+ N_WL<95>_XI0/XI49/XI15/MM9_g N_BL<0>_XI0/XI49/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM6 N_XI0/XI49/XI15/NET35_XI0/XI49/XI15/MM6_d
+ N_XI0/XI49/XI15/NET36_XI0/XI49/XI15/MM6_g N_VSS_XI0/XI49/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM7 N_XI0/XI49/XI15/NET36_XI0/XI49/XI15/MM7_d
+ N_XI0/XI49/XI15/NET35_XI0/XI49/XI15/MM7_g N_VSS_XI0/XI49/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM8 N_XI0/XI49/XI15/NET35_XI0/XI49/XI15/MM8_d
+ N_WL<95>_XI0/XI49/XI15/MM8_g N_BLN<0>_XI0/XI49/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI49/XI15/MM5 N_XI0/XI49/XI15/NET34_XI0/XI49/XI15/MM5_d
+ N_XI0/XI49/XI15/NET33_XI0/XI49/XI15/MM5_g N_VDD_XI0/XI49/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI15/MM4 N_XI0/XI49/XI15/NET33_XI0/XI49/XI15/MM4_d
+ N_XI0/XI49/XI15/NET34_XI0/XI49/XI15/MM4_g N_VDD_XI0/XI49/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI15/MM10 N_XI0/XI49/XI15/NET35_XI0/XI49/XI15/MM10_d
+ N_XI0/XI49/XI15/NET36_XI0/XI49/XI15/MM10_g N_VDD_XI0/XI49/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI49/XI15/MM11 N_XI0/XI49/XI15/NET36_XI0/XI49/XI15/MM11_d
+ N_XI0/XI49/XI15/NET35_XI0/XI49/XI15/MM11_g N_VDD_XI0/XI49/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI0/MM2 N_XI0/XI50/XI0/NET34_XI0/XI50/XI0/MM2_d
+ N_XI0/XI50/XI0/NET33_XI0/XI50/XI0/MM2_g N_VSS_XI0/XI50/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM3 N_XI0/XI50/XI0/NET33_XI0/XI50/XI0/MM3_d
+ N_WL<96>_XI0/XI50/XI0/MM3_g N_BLN<15>_XI0/XI50/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM0 N_XI0/XI50/XI0/NET34_XI0/XI50/XI0/MM0_d
+ N_WL<96>_XI0/XI50/XI0/MM0_g N_BL<15>_XI0/XI50/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM1 N_XI0/XI50/XI0/NET33_XI0/XI50/XI0/MM1_d
+ N_XI0/XI50/XI0/NET34_XI0/XI50/XI0/MM1_g N_VSS_XI0/XI50/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM9 N_XI0/XI50/XI0/NET36_XI0/XI50/XI0/MM9_d
+ N_WL<97>_XI0/XI50/XI0/MM9_g N_BL<15>_XI0/XI50/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM6 N_XI0/XI50/XI0/NET35_XI0/XI50/XI0/MM6_d
+ N_XI0/XI50/XI0/NET36_XI0/XI50/XI0/MM6_g N_VSS_XI0/XI50/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM7 N_XI0/XI50/XI0/NET36_XI0/XI50/XI0/MM7_d
+ N_XI0/XI50/XI0/NET35_XI0/XI50/XI0/MM7_g N_VSS_XI0/XI50/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM8 N_XI0/XI50/XI0/NET35_XI0/XI50/XI0/MM8_d
+ N_WL<97>_XI0/XI50/XI0/MM8_g N_BLN<15>_XI0/XI50/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI0/MM5 N_XI0/XI50/XI0/NET34_XI0/XI50/XI0/MM5_d
+ N_XI0/XI50/XI0/NET33_XI0/XI50/XI0/MM5_g N_VDD_XI0/XI50/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI0/MM4 N_XI0/XI50/XI0/NET33_XI0/XI50/XI0/MM4_d
+ N_XI0/XI50/XI0/NET34_XI0/XI50/XI0/MM4_g N_VDD_XI0/XI50/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI0/MM10 N_XI0/XI50/XI0/NET35_XI0/XI50/XI0/MM10_d
+ N_XI0/XI50/XI0/NET36_XI0/XI50/XI0/MM10_g N_VDD_XI0/XI50/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI0/MM11 N_XI0/XI50/XI0/NET36_XI0/XI50/XI0/MM11_d
+ N_XI0/XI50/XI0/NET35_XI0/XI50/XI0/MM11_g N_VDD_XI0/XI50/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI1/MM2 N_XI0/XI50/XI1/NET34_XI0/XI50/XI1/MM2_d
+ N_XI0/XI50/XI1/NET33_XI0/XI50/XI1/MM2_g N_VSS_XI0/XI50/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM3 N_XI0/XI50/XI1/NET33_XI0/XI50/XI1/MM3_d
+ N_WL<96>_XI0/XI50/XI1/MM3_g N_BLN<14>_XI0/XI50/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM0 N_XI0/XI50/XI1/NET34_XI0/XI50/XI1/MM0_d
+ N_WL<96>_XI0/XI50/XI1/MM0_g N_BL<14>_XI0/XI50/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM1 N_XI0/XI50/XI1/NET33_XI0/XI50/XI1/MM1_d
+ N_XI0/XI50/XI1/NET34_XI0/XI50/XI1/MM1_g N_VSS_XI0/XI50/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM9 N_XI0/XI50/XI1/NET36_XI0/XI50/XI1/MM9_d
+ N_WL<97>_XI0/XI50/XI1/MM9_g N_BL<14>_XI0/XI50/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM6 N_XI0/XI50/XI1/NET35_XI0/XI50/XI1/MM6_d
+ N_XI0/XI50/XI1/NET36_XI0/XI50/XI1/MM6_g N_VSS_XI0/XI50/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM7 N_XI0/XI50/XI1/NET36_XI0/XI50/XI1/MM7_d
+ N_XI0/XI50/XI1/NET35_XI0/XI50/XI1/MM7_g N_VSS_XI0/XI50/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM8 N_XI0/XI50/XI1/NET35_XI0/XI50/XI1/MM8_d
+ N_WL<97>_XI0/XI50/XI1/MM8_g N_BLN<14>_XI0/XI50/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI1/MM5 N_XI0/XI50/XI1/NET34_XI0/XI50/XI1/MM5_d
+ N_XI0/XI50/XI1/NET33_XI0/XI50/XI1/MM5_g N_VDD_XI0/XI50/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI1/MM4 N_XI0/XI50/XI1/NET33_XI0/XI50/XI1/MM4_d
+ N_XI0/XI50/XI1/NET34_XI0/XI50/XI1/MM4_g N_VDD_XI0/XI50/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI1/MM10 N_XI0/XI50/XI1/NET35_XI0/XI50/XI1/MM10_d
+ N_XI0/XI50/XI1/NET36_XI0/XI50/XI1/MM10_g N_VDD_XI0/XI50/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI1/MM11 N_XI0/XI50/XI1/NET36_XI0/XI50/XI1/MM11_d
+ N_XI0/XI50/XI1/NET35_XI0/XI50/XI1/MM11_g N_VDD_XI0/XI50/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI2/MM2 N_XI0/XI50/XI2/NET34_XI0/XI50/XI2/MM2_d
+ N_XI0/XI50/XI2/NET33_XI0/XI50/XI2/MM2_g N_VSS_XI0/XI50/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM3 N_XI0/XI50/XI2/NET33_XI0/XI50/XI2/MM3_d
+ N_WL<96>_XI0/XI50/XI2/MM3_g N_BLN<13>_XI0/XI50/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM0 N_XI0/XI50/XI2/NET34_XI0/XI50/XI2/MM0_d
+ N_WL<96>_XI0/XI50/XI2/MM0_g N_BL<13>_XI0/XI50/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM1 N_XI0/XI50/XI2/NET33_XI0/XI50/XI2/MM1_d
+ N_XI0/XI50/XI2/NET34_XI0/XI50/XI2/MM1_g N_VSS_XI0/XI50/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM9 N_XI0/XI50/XI2/NET36_XI0/XI50/XI2/MM9_d
+ N_WL<97>_XI0/XI50/XI2/MM9_g N_BL<13>_XI0/XI50/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM6 N_XI0/XI50/XI2/NET35_XI0/XI50/XI2/MM6_d
+ N_XI0/XI50/XI2/NET36_XI0/XI50/XI2/MM6_g N_VSS_XI0/XI50/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM7 N_XI0/XI50/XI2/NET36_XI0/XI50/XI2/MM7_d
+ N_XI0/XI50/XI2/NET35_XI0/XI50/XI2/MM7_g N_VSS_XI0/XI50/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM8 N_XI0/XI50/XI2/NET35_XI0/XI50/XI2/MM8_d
+ N_WL<97>_XI0/XI50/XI2/MM8_g N_BLN<13>_XI0/XI50/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI2/MM5 N_XI0/XI50/XI2/NET34_XI0/XI50/XI2/MM5_d
+ N_XI0/XI50/XI2/NET33_XI0/XI50/XI2/MM5_g N_VDD_XI0/XI50/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI2/MM4 N_XI0/XI50/XI2/NET33_XI0/XI50/XI2/MM4_d
+ N_XI0/XI50/XI2/NET34_XI0/XI50/XI2/MM4_g N_VDD_XI0/XI50/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI2/MM10 N_XI0/XI50/XI2/NET35_XI0/XI50/XI2/MM10_d
+ N_XI0/XI50/XI2/NET36_XI0/XI50/XI2/MM10_g N_VDD_XI0/XI50/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI2/MM11 N_XI0/XI50/XI2/NET36_XI0/XI50/XI2/MM11_d
+ N_XI0/XI50/XI2/NET35_XI0/XI50/XI2/MM11_g N_VDD_XI0/XI50/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI3/MM2 N_XI0/XI50/XI3/NET34_XI0/XI50/XI3/MM2_d
+ N_XI0/XI50/XI3/NET33_XI0/XI50/XI3/MM2_g N_VSS_XI0/XI50/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM3 N_XI0/XI50/XI3/NET33_XI0/XI50/XI3/MM3_d
+ N_WL<96>_XI0/XI50/XI3/MM3_g N_BLN<12>_XI0/XI50/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM0 N_XI0/XI50/XI3/NET34_XI0/XI50/XI3/MM0_d
+ N_WL<96>_XI0/XI50/XI3/MM0_g N_BL<12>_XI0/XI50/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM1 N_XI0/XI50/XI3/NET33_XI0/XI50/XI3/MM1_d
+ N_XI0/XI50/XI3/NET34_XI0/XI50/XI3/MM1_g N_VSS_XI0/XI50/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM9 N_XI0/XI50/XI3/NET36_XI0/XI50/XI3/MM9_d
+ N_WL<97>_XI0/XI50/XI3/MM9_g N_BL<12>_XI0/XI50/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM6 N_XI0/XI50/XI3/NET35_XI0/XI50/XI3/MM6_d
+ N_XI0/XI50/XI3/NET36_XI0/XI50/XI3/MM6_g N_VSS_XI0/XI50/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM7 N_XI0/XI50/XI3/NET36_XI0/XI50/XI3/MM7_d
+ N_XI0/XI50/XI3/NET35_XI0/XI50/XI3/MM7_g N_VSS_XI0/XI50/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM8 N_XI0/XI50/XI3/NET35_XI0/XI50/XI3/MM8_d
+ N_WL<97>_XI0/XI50/XI3/MM8_g N_BLN<12>_XI0/XI50/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI3/MM5 N_XI0/XI50/XI3/NET34_XI0/XI50/XI3/MM5_d
+ N_XI0/XI50/XI3/NET33_XI0/XI50/XI3/MM5_g N_VDD_XI0/XI50/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI3/MM4 N_XI0/XI50/XI3/NET33_XI0/XI50/XI3/MM4_d
+ N_XI0/XI50/XI3/NET34_XI0/XI50/XI3/MM4_g N_VDD_XI0/XI50/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI3/MM10 N_XI0/XI50/XI3/NET35_XI0/XI50/XI3/MM10_d
+ N_XI0/XI50/XI3/NET36_XI0/XI50/XI3/MM10_g N_VDD_XI0/XI50/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI3/MM11 N_XI0/XI50/XI3/NET36_XI0/XI50/XI3/MM11_d
+ N_XI0/XI50/XI3/NET35_XI0/XI50/XI3/MM11_g N_VDD_XI0/XI50/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI4/MM2 N_XI0/XI50/XI4/NET34_XI0/XI50/XI4/MM2_d
+ N_XI0/XI50/XI4/NET33_XI0/XI50/XI4/MM2_g N_VSS_XI0/XI50/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM3 N_XI0/XI50/XI4/NET33_XI0/XI50/XI4/MM3_d
+ N_WL<96>_XI0/XI50/XI4/MM3_g N_BLN<11>_XI0/XI50/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM0 N_XI0/XI50/XI4/NET34_XI0/XI50/XI4/MM0_d
+ N_WL<96>_XI0/XI50/XI4/MM0_g N_BL<11>_XI0/XI50/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM1 N_XI0/XI50/XI4/NET33_XI0/XI50/XI4/MM1_d
+ N_XI0/XI50/XI4/NET34_XI0/XI50/XI4/MM1_g N_VSS_XI0/XI50/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM9 N_XI0/XI50/XI4/NET36_XI0/XI50/XI4/MM9_d
+ N_WL<97>_XI0/XI50/XI4/MM9_g N_BL<11>_XI0/XI50/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM6 N_XI0/XI50/XI4/NET35_XI0/XI50/XI4/MM6_d
+ N_XI0/XI50/XI4/NET36_XI0/XI50/XI4/MM6_g N_VSS_XI0/XI50/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM7 N_XI0/XI50/XI4/NET36_XI0/XI50/XI4/MM7_d
+ N_XI0/XI50/XI4/NET35_XI0/XI50/XI4/MM7_g N_VSS_XI0/XI50/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM8 N_XI0/XI50/XI4/NET35_XI0/XI50/XI4/MM8_d
+ N_WL<97>_XI0/XI50/XI4/MM8_g N_BLN<11>_XI0/XI50/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI4/MM5 N_XI0/XI50/XI4/NET34_XI0/XI50/XI4/MM5_d
+ N_XI0/XI50/XI4/NET33_XI0/XI50/XI4/MM5_g N_VDD_XI0/XI50/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI4/MM4 N_XI0/XI50/XI4/NET33_XI0/XI50/XI4/MM4_d
+ N_XI0/XI50/XI4/NET34_XI0/XI50/XI4/MM4_g N_VDD_XI0/XI50/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI4/MM10 N_XI0/XI50/XI4/NET35_XI0/XI50/XI4/MM10_d
+ N_XI0/XI50/XI4/NET36_XI0/XI50/XI4/MM10_g N_VDD_XI0/XI50/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI4/MM11 N_XI0/XI50/XI4/NET36_XI0/XI50/XI4/MM11_d
+ N_XI0/XI50/XI4/NET35_XI0/XI50/XI4/MM11_g N_VDD_XI0/XI50/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI5/MM2 N_XI0/XI50/XI5/NET34_XI0/XI50/XI5/MM2_d
+ N_XI0/XI50/XI5/NET33_XI0/XI50/XI5/MM2_g N_VSS_XI0/XI50/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM3 N_XI0/XI50/XI5/NET33_XI0/XI50/XI5/MM3_d
+ N_WL<96>_XI0/XI50/XI5/MM3_g N_BLN<10>_XI0/XI50/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM0 N_XI0/XI50/XI5/NET34_XI0/XI50/XI5/MM0_d
+ N_WL<96>_XI0/XI50/XI5/MM0_g N_BL<10>_XI0/XI50/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM1 N_XI0/XI50/XI5/NET33_XI0/XI50/XI5/MM1_d
+ N_XI0/XI50/XI5/NET34_XI0/XI50/XI5/MM1_g N_VSS_XI0/XI50/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM9 N_XI0/XI50/XI5/NET36_XI0/XI50/XI5/MM9_d
+ N_WL<97>_XI0/XI50/XI5/MM9_g N_BL<10>_XI0/XI50/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM6 N_XI0/XI50/XI5/NET35_XI0/XI50/XI5/MM6_d
+ N_XI0/XI50/XI5/NET36_XI0/XI50/XI5/MM6_g N_VSS_XI0/XI50/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM7 N_XI0/XI50/XI5/NET36_XI0/XI50/XI5/MM7_d
+ N_XI0/XI50/XI5/NET35_XI0/XI50/XI5/MM7_g N_VSS_XI0/XI50/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM8 N_XI0/XI50/XI5/NET35_XI0/XI50/XI5/MM8_d
+ N_WL<97>_XI0/XI50/XI5/MM8_g N_BLN<10>_XI0/XI50/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI5/MM5 N_XI0/XI50/XI5/NET34_XI0/XI50/XI5/MM5_d
+ N_XI0/XI50/XI5/NET33_XI0/XI50/XI5/MM5_g N_VDD_XI0/XI50/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI5/MM4 N_XI0/XI50/XI5/NET33_XI0/XI50/XI5/MM4_d
+ N_XI0/XI50/XI5/NET34_XI0/XI50/XI5/MM4_g N_VDD_XI0/XI50/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI5/MM10 N_XI0/XI50/XI5/NET35_XI0/XI50/XI5/MM10_d
+ N_XI0/XI50/XI5/NET36_XI0/XI50/XI5/MM10_g N_VDD_XI0/XI50/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI5/MM11 N_XI0/XI50/XI5/NET36_XI0/XI50/XI5/MM11_d
+ N_XI0/XI50/XI5/NET35_XI0/XI50/XI5/MM11_g N_VDD_XI0/XI50/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI6/MM2 N_XI0/XI50/XI6/NET34_XI0/XI50/XI6/MM2_d
+ N_XI0/XI50/XI6/NET33_XI0/XI50/XI6/MM2_g N_VSS_XI0/XI50/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM3 N_XI0/XI50/XI6/NET33_XI0/XI50/XI6/MM3_d
+ N_WL<96>_XI0/XI50/XI6/MM3_g N_BLN<9>_XI0/XI50/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM0 N_XI0/XI50/XI6/NET34_XI0/XI50/XI6/MM0_d
+ N_WL<96>_XI0/XI50/XI6/MM0_g N_BL<9>_XI0/XI50/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM1 N_XI0/XI50/XI6/NET33_XI0/XI50/XI6/MM1_d
+ N_XI0/XI50/XI6/NET34_XI0/XI50/XI6/MM1_g N_VSS_XI0/XI50/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM9 N_XI0/XI50/XI6/NET36_XI0/XI50/XI6/MM9_d
+ N_WL<97>_XI0/XI50/XI6/MM9_g N_BL<9>_XI0/XI50/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM6 N_XI0/XI50/XI6/NET35_XI0/XI50/XI6/MM6_d
+ N_XI0/XI50/XI6/NET36_XI0/XI50/XI6/MM6_g N_VSS_XI0/XI50/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM7 N_XI0/XI50/XI6/NET36_XI0/XI50/XI6/MM7_d
+ N_XI0/XI50/XI6/NET35_XI0/XI50/XI6/MM7_g N_VSS_XI0/XI50/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM8 N_XI0/XI50/XI6/NET35_XI0/XI50/XI6/MM8_d
+ N_WL<97>_XI0/XI50/XI6/MM8_g N_BLN<9>_XI0/XI50/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI6/MM5 N_XI0/XI50/XI6/NET34_XI0/XI50/XI6/MM5_d
+ N_XI0/XI50/XI6/NET33_XI0/XI50/XI6/MM5_g N_VDD_XI0/XI50/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI6/MM4 N_XI0/XI50/XI6/NET33_XI0/XI50/XI6/MM4_d
+ N_XI0/XI50/XI6/NET34_XI0/XI50/XI6/MM4_g N_VDD_XI0/XI50/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI6/MM10 N_XI0/XI50/XI6/NET35_XI0/XI50/XI6/MM10_d
+ N_XI0/XI50/XI6/NET36_XI0/XI50/XI6/MM10_g N_VDD_XI0/XI50/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI6/MM11 N_XI0/XI50/XI6/NET36_XI0/XI50/XI6/MM11_d
+ N_XI0/XI50/XI6/NET35_XI0/XI50/XI6/MM11_g N_VDD_XI0/XI50/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI7/MM2 N_XI0/XI50/XI7/NET34_XI0/XI50/XI7/MM2_d
+ N_XI0/XI50/XI7/NET33_XI0/XI50/XI7/MM2_g N_VSS_XI0/XI50/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM3 N_XI0/XI50/XI7/NET33_XI0/XI50/XI7/MM3_d
+ N_WL<96>_XI0/XI50/XI7/MM3_g N_BLN<8>_XI0/XI50/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM0 N_XI0/XI50/XI7/NET34_XI0/XI50/XI7/MM0_d
+ N_WL<96>_XI0/XI50/XI7/MM0_g N_BL<8>_XI0/XI50/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM1 N_XI0/XI50/XI7/NET33_XI0/XI50/XI7/MM1_d
+ N_XI0/XI50/XI7/NET34_XI0/XI50/XI7/MM1_g N_VSS_XI0/XI50/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM9 N_XI0/XI50/XI7/NET36_XI0/XI50/XI7/MM9_d
+ N_WL<97>_XI0/XI50/XI7/MM9_g N_BL<8>_XI0/XI50/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM6 N_XI0/XI50/XI7/NET35_XI0/XI50/XI7/MM6_d
+ N_XI0/XI50/XI7/NET36_XI0/XI50/XI7/MM6_g N_VSS_XI0/XI50/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM7 N_XI0/XI50/XI7/NET36_XI0/XI50/XI7/MM7_d
+ N_XI0/XI50/XI7/NET35_XI0/XI50/XI7/MM7_g N_VSS_XI0/XI50/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM8 N_XI0/XI50/XI7/NET35_XI0/XI50/XI7/MM8_d
+ N_WL<97>_XI0/XI50/XI7/MM8_g N_BLN<8>_XI0/XI50/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI7/MM5 N_XI0/XI50/XI7/NET34_XI0/XI50/XI7/MM5_d
+ N_XI0/XI50/XI7/NET33_XI0/XI50/XI7/MM5_g N_VDD_XI0/XI50/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI7/MM4 N_XI0/XI50/XI7/NET33_XI0/XI50/XI7/MM4_d
+ N_XI0/XI50/XI7/NET34_XI0/XI50/XI7/MM4_g N_VDD_XI0/XI50/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI7/MM10 N_XI0/XI50/XI7/NET35_XI0/XI50/XI7/MM10_d
+ N_XI0/XI50/XI7/NET36_XI0/XI50/XI7/MM10_g N_VDD_XI0/XI50/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI7/MM11 N_XI0/XI50/XI7/NET36_XI0/XI50/XI7/MM11_d
+ N_XI0/XI50/XI7/NET35_XI0/XI50/XI7/MM11_g N_VDD_XI0/XI50/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI8/MM2 N_XI0/XI50/XI8/NET34_XI0/XI50/XI8/MM2_d
+ N_XI0/XI50/XI8/NET33_XI0/XI50/XI8/MM2_g N_VSS_XI0/XI50/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM3 N_XI0/XI50/XI8/NET33_XI0/XI50/XI8/MM3_d
+ N_WL<96>_XI0/XI50/XI8/MM3_g N_BLN<7>_XI0/XI50/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM0 N_XI0/XI50/XI8/NET34_XI0/XI50/XI8/MM0_d
+ N_WL<96>_XI0/XI50/XI8/MM0_g N_BL<7>_XI0/XI50/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM1 N_XI0/XI50/XI8/NET33_XI0/XI50/XI8/MM1_d
+ N_XI0/XI50/XI8/NET34_XI0/XI50/XI8/MM1_g N_VSS_XI0/XI50/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM9 N_XI0/XI50/XI8/NET36_XI0/XI50/XI8/MM9_d
+ N_WL<97>_XI0/XI50/XI8/MM9_g N_BL<7>_XI0/XI50/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM6 N_XI0/XI50/XI8/NET35_XI0/XI50/XI8/MM6_d
+ N_XI0/XI50/XI8/NET36_XI0/XI50/XI8/MM6_g N_VSS_XI0/XI50/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM7 N_XI0/XI50/XI8/NET36_XI0/XI50/XI8/MM7_d
+ N_XI0/XI50/XI8/NET35_XI0/XI50/XI8/MM7_g N_VSS_XI0/XI50/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM8 N_XI0/XI50/XI8/NET35_XI0/XI50/XI8/MM8_d
+ N_WL<97>_XI0/XI50/XI8/MM8_g N_BLN<7>_XI0/XI50/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI8/MM5 N_XI0/XI50/XI8/NET34_XI0/XI50/XI8/MM5_d
+ N_XI0/XI50/XI8/NET33_XI0/XI50/XI8/MM5_g N_VDD_XI0/XI50/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI8/MM4 N_XI0/XI50/XI8/NET33_XI0/XI50/XI8/MM4_d
+ N_XI0/XI50/XI8/NET34_XI0/XI50/XI8/MM4_g N_VDD_XI0/XI50/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI8/MM10 N_XI0/XI50/XI8/NET35_XI0/XI50/XI8/MM10_d
+ N_XI0/XI50/XI8/NET36_XI0/XI50/XI8/MM10_g N_VDD_XI0/XI50/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI8/MM11 N_XI0/XI50/XI8/NET36_XI0/XI50/XI8/MM11_d
+ N_XI0/XI50/XI8/NET35_XI0/XI50/XI8/MM11_g N_VDD_XI0/XI50/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI9/MM2 N_XI0/XI50/XI9/NET34_XI0/XI50/XI9/MM2_d
+ N_XI0/XI50/XI9/NET33_XI0/XI50/XI9/MM2_g N_VSS_XI0/XI50/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM3 N_XI0/XI50/XI9/NET33_XI0/XI50/XI9/MM3_d
+ N_WL<96>_XI0/XI50/XI9/MM3_g N_BLN<6>_XI0/XI50/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM0 N_XI0/XI50/XI9/NET34_XI0/XI50/XI9/MM0_d
+ N_WL<96>_XI0/XI50/XI9/MM0_g N_BL<6>_XI0/XI50/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM1 N_XI0/XI50/XI9/NET33_XI0/XI50/XI9/MM1_d
+ N_XI0/XI50/XI9/NET34_XI0/XI50/XI9/MM1_g N_VSS_XI0/XI50/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM9 N_XI0/XI50/XI9/NET36_XI0/XI50/XI9/MM9_d
+ N_WL<97>_XI0/XI50/XI9/MM9_g N_BL<6>_XI0/XI50/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM6 N_XI0/XI50/XI9/NET35_XI0/XI50/XI9/MM6_d
+ N_XI0/XI50/XI9/NET36_XI0/XI50/XI9/MM6_g N_VSS_XI0/XI50/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM7 N_XI0/XI50/XI9/NET36_XI0/XI50/XI9/MM7_d
+ N_XI0/XI50/XI9/NET35_XI0/XI50/XI9/MM7_g N_VSS_XI0/XI50/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM8 N_XI0/XI50/XI9/NET35_XI0/XI50/XI9/MM8_d
+ N_WL<97>_XI0/XI50/XI9/MM8_g N_BLN<6>_XI0/XI50/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI9/MM5 N_XI0/XI50/XI9/NET34_XI0/XI50/XI9/MM5_d
+ N_XI0/XI50/XI9/NET33_XI0/XI50/XI9/MM5_g N_VDD_XI0/XI50/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI9/MM4 N_XI0/XI50/XI9/NET33_XI0/XI50/XI9/MM4_d
+ N_XI0/XI50/XI9/NET34_XI0/XI50/XI9/MM4_g N_VDD_XI0/XI50/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI9/MM10 N_XI0/XI50/XI9/NET35_XI0/XI50/XI9/MM10_d
+ N_XI0/XI50/XI9/NET36_XI0/XI50/XI9/MM10_g N_VDD_XI0/XI50/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI9/MM11 N_XI0/XI50/XI9/NET36_XI0/XI50/XI9/MM11_d
+ N_XI0/XI50/XI9/NET35_XI0/XI50/XI9/MM11_g N_VDD_XI0/XI50/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI10/MM2 N_XI0/XI50/XI10/NET34_XI0/XI50/XI10/MM2_d
+ N_XI0/XI50/XI10/NET33_XI0/XI50/XI10/MM2_g N_VSS_XI0/XI50/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM3 N_XI0/XI50/XI10/NET33_XI0/XI50/XI10/MM3_d
+ N_WL<96>_XI0/XI50/XI10/MM3_g N_BLN<5>_XI0/XI50/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM0 N_XI0/XI50/XI10/NET34_XI0/XI50/XI10/MM0_d
+ N_WL<96>_XI0/XI50/XI10/MM0_g N_BL<5>_XI0/XI50/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM1 N_XI0/XI50/XI10/NET33_XI0/XI50/XI10/MM1_d
+ N_XI0/XI50/XI10/NET34_XI0/XI50/XI10/MM1_g N_VSS_XI0/XI50/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM9 N_XI0/XI50/XI10/NET36_XI0/XI50/XI10/MM9_d
+ N_WL<97>_XI0/XI50/XI10/MM9_g N_BL<5>_XI0/XI50/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM6 N_XI0/XI50/XI10/NET35_XI0/XI50/XI10/MM6_d
+ N_XI0/XI50/XI10/NET36_XI0/XI50/XI10/MM6_g N_VSS_XI0/XI50/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM7 N_XI0/XI50/XI10/NET36_XI0/XI50/XI10/MM7_d
+ N_XI0/XI50/XI10/NET35_XI0/XI50/XI10/MM7_g N_VSS_XI0/XI50/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM8 N_XI0/XI50/XI10/NET35_XI0/XI50/XI10/MM8_d
+ N_WL<97>_XI0/XI50/XI10/MM8_g N_BLN<5>_XI0/XI50/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI10/MM5 N_XI0/XI50/XI10/NET34_XI0/XI50/XI10/MM5_d
+ N_XI0/XI50/XI10/NET33_XI0/XI50/XI10/MM5_g N_VDD_XI0/XI50/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI10/MM4 N_XI0/XI50/XI10/NET33_XI0/XI50/XI10/MM4_d
+ N_XI0/XI50/XI10/NET34_XI0/XI50/XI10/MM4_g N_VDD_XI0/XI50/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI10/MM10 N_XI0/XI50/XI10/NET35_XI0/XI50/XI10/MM10_d
+ N_XI0/XI50/XI10/NET36_XI0/XI50/XI10/MM10_g N_VDD_XI0/XI50/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI10/MM11 N_XI0/XI50/XI10/NET36_XI0/XI50/XI10/MM11_d
+ N_XI0/XI50/XI10/NET35_XI0/XI50/XI10/MM11_g N_VDD_XI0/XI50/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI11/MM2 N_XI0/XI50/XI11/NET34_XI0/XI50/XI11/MM2_d
+ N_XI0/XI50/XI11/NET33_XI0/XI50/XI11/MM2_g N_VSS_XI0/XI50/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM3 N_XI0/XI50/XI11/NET33_XI0/XI50/XI11/MM3_d
+ N_WL<96>_XI0/XI50/XI11/MM3_g N_BLN<4>_XI0/XI50/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM0 N_XI0/XI50/XI11/NET34_XI0/XI50/XI11/MM0_d
+ N_WL<96>_XI0/XI50/XI11/MM0_g N_BL<4>_XI0/XI50/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM1 N_XI0/XI50/XI11/NET33_XI0/XI50/XI11/MM1_d
+ N_XI0/XI50/XI11/NET34_XI0/XI50/XI11/MM1_g N_VSS_XI0/XI50/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM9 N_XI0/XI50/XI11/NET36_XI0/XI50/XI11/MM9_d
+ N_WL<97>_XI0/XI50/XI11/MM9_g N_BL<4>_XI0/XI50/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM6 N_XI0/XI50/XI11/NET35_XI0/XI50/XI11/MM6_d
+ N_XI0/XI50/XI11/NET36_XI0/XI50/XI11/MM6_g N_VSS_XI0/XI50/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM7 N_XI0/XI50/XI11/NET36_XI0/XI50/XI11/MM7_d
+ N_XI0/XI50/XI11/NET35_XI0/XI50/XI11/MM7_g N_VSS_XI0/XI50/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM8 N_XI0/XI50/XI11/NET35_XI0/XI50/XI11/MM8_d
+ N_WL<97>_XI0/XI50/XI11/MM8_g N_BLN<4>_XI0/XI50/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI11/MM5 N_XI0/XI50/XI11/NET34_XI0/XI50/XI11/MM5_d
+ N_XI0/XI50/XI11/NET33_XI0/XI50/XI11/MM5_g N_VDD_XI0/XI50/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI11/MM4 N_XI0/XI50/XI11/NET33_XI0/XI50/XI11/MM4_d
+ N_XI0/XI50/XI11/NET34_XI0/XI50/XI11/MM4_g N_VDD_XI0/XI50/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI11/MM10 N_XI0/XI50/XI11/NET35_XI0/XI50/XI11/MM10_d
+ N_XI0/XI50/XI11/NET36_XI0/XI50/XI11/MM10_g N_VDD_XI0/XI50/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI11/MM11 N_XI0/XI50/XI11/NET36_XI0/XI50/XI11/MM11_d
+ N_XI0/XI50/XI11/NET35_XI0/XI50/XI11/MM11_g N_VDD_XI0/XI50/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI12/MM2 N_XI0/XI50/XI12/NET34_XI0/XI50/XI12/MM2_d
+ N_XI0/XI50/XI12/NET33_XI0/XI50/XI12/MM2_g N_VSS_XI0/XI50/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM3 N_XI0/XI50/XI12/NET33_XI0/XI50/XI12/MM3_d
+ N_WL<96>_XI0/XI50/XI12/MM3_g N_BLN<3>_XI0/XI50/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM0 N_XI0/XI50/XI12/NET34_XI0/XI50/XI12/MM0_d
+ N_WL<96>_XI0/XI50/XI12/MM0_g N_BL<3>_XI0/XI50/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM1 N_XI0/XI50/XI12/NET33_XI0/XI50/XI12/MM1_d
+ N_XI0/XI50/XI12/NET34_XI0/XI50/XI12/MM1_g N_VSS_XI0/XI50/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM9 N_XI0/XI50/XI12/NET36_XI0/XI50/XI12/MM9_d
+ N_WL<97>_XI0/XI50/XI12/MM9_g N_BL<3>_XI0/XI50/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM6 N_XI0/XI50/XI12/NET35_XI0/XI50/XI12/MM6_d
+ N_XI0/XI50/XI12/NET36_XI0/XI50/XI12/MM6_g N_VSS_XI0/XI50/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM7 N_XI0/XI50/XI12/NET36_XI0/XI50/XI12/MM7_d
+ N_XI0/XI50/XI12/NET35_XI0/XI50/XI12/MM7_g N_VSS_XI0/XI50/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM8 N_XI0/XI50/XI12/NET35_XI0/XI50/XI12/MM8_d
+ N_WL<97>_XI0/XI50/XI12/MM8_g N_BLN<3>_XI0/XI50/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI12/MM5 N_XI0/XI50/XI12/NET34_XI0/XI50/XI12/MM5_d
+ N_XI0/XI50/XI12/NET33_XI0/XI50/XI12/MM5_g N_VDD_XI0/XI50/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI12/MM4 N_XI0/XI50/XI12/NET33_XI0/XI50/XI12/MM4_d
+ N_XI0/XI50/XI12/NET34_XI0/XI50/XI12/MM4_g N_VDD_XI0/XI50/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI12/MM10 N_XI0/XI50/XI12/NET35_XI0/XI50/XI12/MM10_d
+ N_XI0/XI50/XI12/NET36_XI0/XI50/XI12/MM10_g N_VDD_XI0/XI50/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI12/MM11 N_XI0/XI50/XI12/NET36_XI0/XI50/XI12/MM11_d
+ N_XI0/XI50/XI12/NET35_XI0/XI50/XI12/MM11_g N_VDD_XI0/XI50/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI13/MM2 N_XI0/XI50/XI13/NET34_XI0/XI50/XI13/MM2_d
+ N_XI0/XI50/XI13/NET33_XI0/XI50/XI13/MM2_g N_VSS_XI0/XI50/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM3 N_XI0/XI50/XI13/NET33_XI0/XI50/XI13/MM3_d
+ N_WL<96>_XI0/XI50/XI13/MM3_g N_BLN<2>_XI0/XI50/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM0 N_XI0/XI50/XI13/NET34_XI0/XI50/XI13/MM0_d
+ N_WL<96>_XI0/XI50/XI13/MM0_g N_BL<2>_XI0/XI50/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM1 N_XI0/XI50/XI13/NET33_XI0/XI50/XI13/MM1_d
+ N_XI0/XI50/XI13/NET34_XI0/XI50/XI13/MM1_g N_VSS_XI0/XI50/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM9 N_XI0/XI50/XI13/NET36_XI0/XI50/XI13/MM9_d
+ N_WL<97>_XI0/XI50/XI13/MM9_g N_BL<2>_XI0/XI50/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM6 N_XI0/XI50/XI13/NET35_XI0/XI50/XI13/MM6_d
+ N_XI0/XI50/XI13/NET36_XI0/XI50/XI13/MM6_g N_VSS_XI0/XI50/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM7 N_XI0/XI50/XI13/NET36_XI0/XI50/XI13/MM7_d
+ N_XI0/XI50/XI13/NET35_XI0/XI50/XI13/MM7_g N_VSS_XI0/XI50/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM8 N_XI0/XI50/XI13/NET35_XI0/XI50/XI13/MM8_d
+ N_WL<97>_XI0/XI50/XI13/MM8_g N_BLN<2>_XI0/XI50/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI13/MM5 N_XI0/XI50/XI13/NET34_XI0/XI50/XI13/MM5_d
+ N_XI0/XI50/XI13/NET33_XI0/XI50/XI13/MM5_g N_VDD_XI0/XI50/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI13/MM4 N_XI0/XI50/XI13/NET33_XI0/XI50/XI13/MM4_d
+ N_XI0/XI50/XI13/NET34_XI0/XI50/XI13/MM4_g N_VDD_XI0/XI50/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI13/MM10 N_XI0/XI50/XI13/NET35_XI0/XI50/XI13/MM10_d
+ N_XI0/XI50/XI13/NET36_XI0/XI50/XI13/MM10_g N_VDD_XI0/XI50/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI13/MM11 N_XI0/XI50/XI13/NET36_XI0/XI50/XI13/MM11_d
+ N_XI0/XI50/XI13/NET35_XI0/XI50/XI13/MM11_g N_VDD_XI0/XI50/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI14/MM2 N_XI0/XI50/XI14/NET34_XI0/XI50/XI14/MM2_d
+ N_XI0/XI50/XI14/NET33_XI0/XI50/XI14/MM2_g N_VSS_XI0/XI50/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM3 N_XI0/XI50/XI14/NET33_XI0/XI50/XI14/MM3_d
+ N_WL<96>_XI0/XI50/XI14/MM3_g N_BLN<1>_XI0/XI50/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM0 N_XI0/XI50/XI14/NET34_XI0/XI50/XI14/MM0_d
+ N_WL<96>_XI0/XI50/XI14/MM0_g N_BL<1>_XI0/XI50/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM1 N_XI0/XI50/XI14/NET33_XI0/XI50/XI14/MM1_d
+ N_XI0/XI50/XI14/NET34_XI0/XI50/XI14/MM1_g N_VSS_XI0/XI50/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM9 N_XI0/XI50/XI14/NET36_XI0/XI50/XI14/MM9_d
+ N_WL<97>_XI0/XI50/XI14/MM9_g N_BL<1>_XI0/XI50/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM6 N_XI0/XI50/XI14/NET35_XI0/XI50/XI14/MM6_d
+ N_XI0/XI50/XI14/NET36_XI0/XI50/XI14/MM6_g N_VSS_XI0/XI50/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM7 N_XI0/XI50/XI14/NET36_XI0/XI50/XI14/MM7_d
+ N_XI0/XI50/XI14/NET35_XI0/XI50/XI14/MM7_g N_VSS_XI0/XI50/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM8 N_XI0/XI50/XI14/NET35_XI0/XI50/XI14/MM8_d
+ N_WL<97>_XI0/XI50/XI14/MM8_g N_BLN<1>_XI0/XI50/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI14/MM5 N_XI0/XI50/XI14/NET34_XI0/XI50/XI14/MM5_d
+ N_XI0/XI50/XI14/NET33_XI0/XI50/XI14/MM5_g N_VDD_XI0/XI50/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI14/MM4 N_XI0/XI50/XI14/NET33_XI0/XI50/XI14/MM4_d
+ N_XI0/XI50/XI14/NET34_XI0/XI50/XI14/MM4_g N_VDD_XI0/XI50/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI14/MM10 N_XI0/XI50/XI14/NET35_XI0/XI50/XI14/MM10_d
+ N_XI0/XI50/XI14/NET36_XI0/XI50/XI14/MM10_g N_VDD_XI0/XI50/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI14/MM11 N_XI0/XI50/XI14/NET36_XI0/XI50/XI14/MM11_d
+ N_XI0/XI50/XI14/NET35_XI0/XI50/XI14/MM11_g N_VDD_XI0/XI50/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI15/MM2 N_XI0/XI50/XI15/NET34_XI0/XI50/XI15/MM2_d
+ N_XI0/XI50/XI15/NET33_XI0/XI50/XI15/MM2_g N_VSS_XI0/XI50/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM3 N_XI0/XI50/XI15/NET33_XI0/XI50/XI15/MM3_d
+ N_WL<96>_XI0/XI50/XI15/MM3_g N_BLN<0>_XI0/XI50/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM0 N_XI0/XI50/XI15/NET34_XI0/XI50/XI15/MM0_d
+ N_WL<96>_XI0/XI50/XI15/MM0_g N_BL<0>_XI0/XI50/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM1 N_XI0/XI50/XI15/NET33_XI0/XI50/XI15/MM1_d
+ N_XI0/XI50/XI15/NET34_XI0/XI50/XI15/MM1_g N_VSS_XI0/XI50/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM9 N_XI0/XI50/XI15/NET36_XI0/XI50/XI15/MM9_d
+ N_WL<97>_XI0/XI50/XI15/MM9_g N_BL<0>_XI0/XI50/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM6 N_XI0/XI50/XI15/NET35_XI0/XI50/XI15/MM6_d
+ N_XI0/XI50/XI15/NET36_XI0/XI50/XI15/MM6_g N_VSS_XI0/XI50/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM7 N_XI0/XI50/XI15/NET36_XI0/XI50/XI15/MM7_d
+ N_XI0/XI50/XI15/NET35_XI0/XI50/XI15/MM7_g N_VSS_XI0/XI50/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM8 N_XI0/XI50/XI15/NET35_XI0/XI50/XI15/MM8_d
+ N_WL<97>_XI0/XI50/XI15/MM8_g N_BLN<0>_XI0/XI50/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI50/XI15/MM5 N_XI0/XI50/XI15/NET34_XI0/XI50/XI15/MM5_d
+ N_XI0/XI50/XI15/NET33_XI0/XI50/XI15/MM5_g N_VDD_XI0/XI50/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI15/MM4 N_XI0/XI50/XI15/NET33_XI0/XI50/XI15/MM4_d
+ N_XI0/XI50/XI15/NET34_XI0/XI50/XI15/MM4_g N_VDD_XI0/XI50/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI15/MM10 N_XI0/XI50/XI15/NET35_XI0/XI50/XI15/MM10_d
+ N_XI0/XI50/XI15/NET36_XI0/XI50/XI15/MM10_g N_VDD_XI0/XI50/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI50/XI15/MM11 N_XI0/XI50/XI15/NET36_XI0/XI50/XI15/MM11_d
+ N_XI0/XI50/XI15/NET35_XI0/XI50/XI15/MM11_g N_VDD_XI0/XI50/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI0/MM2 N_XI0/XI51/XI0/NET34_XI0/XI51/XI0/MM2_d
+ N_XI0/XI51/XI0/NET33_XI0/XI51/XI0/MM2_g N_VSS_XI0/XI51/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM3 N_XI0/XI51/XI0/NET33_XI0/XI51/XI0/MM3_d
+ N_WL<98>_XI0/XI51/XI0/MM3_g N_BLN<15>_XI0/XI51/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM0 N_XI0/XI51/XI0/NET34_XI0/XI51/XI0/MM0_d
+ N_WL<98>_XI0/XI51/XI0/MM0_g N_BL<15>_XI0/XI51/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM1 N_XI0/XI51/XI0/NET33_XI0/XI51/XI0/MM1_d
+ N_XI0/XI51/XI0/NET34_XI0/XI51/XI0/MM1_g N_VSS_XI0/XI51/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM9 N_XI0/XI51/XI0/NET36_XI0/XI51/XI0/MM9_d
+ N_WL<99>_XI0/XI51/XI0/MM9_g N_BL<15>_XI0/XI51/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM6 N_XI0/XI51/XI0/NET35_XI0/XI51/XI0/MM6_d
+ N_XI0/XI51/XI0/NET36_XI0/XI51/XI0/MM6_g N_VSS_XI0/XI51/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM7 N_XI0/XI51/XI0/NET36_XI0/XI51/XI0/MM7_d
+ N_XI0/XI51/XI0/NET35_XI0/XI51/XI0/MM7_g N_VSS_XI0/XI51/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM8 N_XI0/XI51/XI0/NET35_XI0/XI51/XI0/MM8_d
+ N_WL<99>_XI0/XI51/XI0/MM8_g N_BLN<15>_XI0/XI51/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI0/MM5 N_XI0/XI51/XI0/NET34_XI0/XI51/XI0/MM5_d
+ N_XI0/XI51/XI0/NET33_XI0/XI51/XI0/MM5_g N_VDD_XI0/XI51/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI0/MM4 N_XI0/XI51/XI0/NET33_XI0/XI51/XI0/MM4_d
+ N_XI0/XI51/XI0/NET34_XI0/XI51/XI0/MM4_g N_VDD_XI0/XI51/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI0/MM10 N_XI0/XI51/XI0/NET35_XI0/XI51/XI0/MM10_d
+ N_XI0/XI51/XI0/NET36_XI0/XI51/XI0/MM10_g N_VDD_XI0/XI51/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI0/MM11 N_XI0/XI51/XI0/NET36_XI0/XI51/XI0/MM11_d
+ N_XI0/XI51/XI0/NET35_XI0/XI51/XI0/MM11_g N_VDD_XI0/XI51/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI1/MM2 N_XI0/XI51/XI1/NET34_XI0/XI51/XI1/MM2_d
+ N_XI0/XI51/XI1/NET33_XI0/XI51/XI1/MM2_g N_VSS_XI0/XI51/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM3 N_XI0/XI51/XI1/NET33_XI0/XI51/XI1/MM3_d
+ N_WL<98>_XI0/XI51/XI1/MM3_g N_BLN<14>_XI0/XI51/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM0 N_XI0/XI51/XI1/NET34_XI0/XI51/XI1/MM0_d
+ N_WL<98>_XI0/XI51/XI1/MM0_g N_BL<14>_XI0/XI51/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM1 N_XI0/XI51/XI1/NET33_XI0/XI51/XI1/MM1_d
+ N_XI0/XI51/XI1/NET34_XI0/XI51/XI1/MM1_g N_VSS_XI0/XI51/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM9 N_XI0/XI51/XI1/NET36_XI0/XI51/XI1/MM9_d
+ N_WL<99>_XI0/XI51/XI1/MM9_g N_BL<14>_XI0/XI51/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM6 N_XI0/XI51/XI1/NET35_XI0/XI51/XI1/MM6_d
+ N_XI0/XI51/XI1/NET36_XI0/XI51/XI1/MM6_g N_VSS_XI0/XI51/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM7 N_XI0/XI51/XI1/NET36_XI0/XI51/XI1/MM7_d
+ N_XI0/XI51/XI1/NET35_XI0/XI51/XI1/MM7_g N_VSS_XI0/XI51/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM8 N_XI0/XI51/XI1/NET35_XI0/XI51/XI1/MM8_d
+ N_WL<99>_XI0/XI51/XI1/MM8_g N_BLN<14>_XI0/XI51/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI1/MM5 N_XI0/XI51/XI1/NET34_XI0/XI51/XI1/MM5_d
+ N_XI0/XI51/XI1/NET33_XI0/XI51/XI1/MM5_g N_VDD_XI0/XI51/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI1/MM4 N_XI0/XI51/XI1/NET33_XI0/XI51/XI1/MM4_d
+ N_XI0/XI51/XI1/NET34_XI0/XI51/XI1/MM4_g N_VDD_XI0/XI51/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI1/MM10 N_XI0/XI51/XI1/NET35_XI0/XI51/XI1/MM10_d
+ N_XI0/XI51/XI1/NET36_XI0/XI51/XI1/MM10_g N_VDD_XI0/XI51/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI1/MM11 N_XI0/XI51/XI1/NET36_XI0/XI51/XI1/MM11_d
+ N_XI0/XI51/XI1/NET35_XI0/XI51/XI1/MM11_g N_VDD_XI0/XI51/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI2/MM2 N_XI0/XI51/XI2/NET34_XI0/XI51/XI2/MM2_d
+ N_XI0/XI51/XI2/NET33_XI0/XI51/XI2/MM2_g N_VSS_XI0/XI51/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM3 N_XI0/XI51/XI2/NET33_XI0/XI51/XI2/MM3_d
+ N_WL<98>_XI0/XI51/XI2/MM3_g N_BLN<13>_XI0/XI51/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM0 N_XI0/XI51/XI2/NET34_XI0/XI51/XI2/MM0_d
+ N_WL<98>_XI0/XI51/XI2/MM0_g N_BL<13>_XI0/XI51/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM1 N_XI0/XI51/XI2/NET33_XI0/XI51/XI2/MM1_d
+ N_XI0/XI51/XI2/NET34_XI0/XI51/XI2/MM1_g N_VSS_XI0/XI51/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM9 N_XI0/XI51/XI2/NET36_XI0/XI51/XI2/MM9_d
+ N_WL<99>_XI0/XI51/XI2/MM9_g N_BL<13>_XI0/XI51/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM6 N_XI0/XI51/XI2/NET35_XI0/XI51/XI2/MM6_d
+ N_XI0/XI51/XI2/NET36_XI0/XI51/XI2/MM6_g N_VSS_XI0/XI51/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM7 N_XI0/XI51/XI2/NET36_XI0/XI51/XI2/MM7_d
+ N_XI0/XI51/XI2/NET35_XI0/XI51/XI2/MM7_g N_VSS_XI0/XI51/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM8 N_XI0/XI51/XI2/NET35_XI0/XI51/XI2/MM8_d
+ N_WL<99>_XI0/XI51/XI2/MM8_g N_BLN<13>_XI0/XI51/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI2/MM5 N_XI0/XI51/XI2/NET34_XI0/XI51/XI2/MM5_d
+ N_XI0/XI51/XI2/NET33_XI0/XI51/XI2/MM5_g N_VDD_XI0/XI51/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI2/MM4 N_XI0/XI51/XI2/NET33_XI0/XI51/XI2/MM4_d
+ N_XI0/XI51/XI2/NET34_XI0/XI51/XI2/MM4_g N_VDD_XI0/XI51/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI2/MM10 N_XI0/XI51/XI2/NET35_XI0/XI51/XI2/MM10_d
+ N_XI0/XI51/XI2/NET36_XI0/XI51/XI2/MM10_g N_VDD_XI0/XI51/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI2/MM11 N_XI0/XI51/XI2/NET36_XI0/XI51/XI2/MM11_d
+ N_XI0/XI51/XI2/NET35_XI0/XI51/XI2/MM11_g N_VDD_XI0/XI51/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI3/MM2 N_XI0/XI51/XI3/NET34_XI0/XI51/XI3/MM2_d
+ N_XI0/XI51/XI3/NET33_XI0/XI51/XI3/MM2_g N_VSS_XI0/XI51/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM3 N_XI0/XI51/XI3/NET33_XI0/XI51/XI3/MM3_d
+ N_WL<98>_XI0/XI51/XI3/MM3_g N_BLN<12>_XI0/XI51/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM0 N_XI0/XI51/XI3/NET34_XI0/XI51/XI3/MM0_d
+ N_WL<98>_XI0/XI51/XI3/MM0_g N_BL<12>_XI0/XI51/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM1 N_XI0/XI51/XI3/NET33_XI0/XI51/XI3/MM1_d
+ N_XI0/XI51/XI3/NET34_XI0/XI51/XI3/MM1_g N_VSS_XI0/XI51/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM9 N_XI0/XI51/XI3/NET36_XI0/XI51/XI3/MM9_d
+ N_WL<99>_XI0/XI51/XI3/MM9_g N_BL<12>_XI0/XI51/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM6 N_XI0/XI51/XI3/NET35_XI0/XI51/XI3/MM6_d
+ N_XI0/XI51/XI3/NET36_XI0/XI51/XI3/MM6_g N_VSS_XI0/XI51/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM7 N_XI0/XI51/XI3/NET36_XI0/XI51/XI3/MM7_d
+ N_XI0/XI51/XI3/NET35_XI0/XI51/XI3/MM7_g N_VSS_XI0/XI51/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM8 N_XI0/XI51/XI3/NET35_XI0/XI51/XI3/MM8_d
+ N_WL<99>_XI0/XI51/XI3/MM8_g N_BLN<12>_XI0/XI51/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI3/MM5 N_XI0/XI51/XI3/NET34_XI0/XI51/XI3/MM5_d
+ N_XI0/XI51/XI3/NET33_XI0/XI51/XI3/MM5_g N_VDD_XI0/XI51/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI3/MM4 N_XI0/XI51/XI3/NET33_XI0/XI51/XI3/MM4_d
+ N_XI0/XI51/XI3/NET34_XI0/XI51/XI3/MM4_g N_VDD_XI0/XI51/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI3/MM10 N_XI0/XI51/XI3/NET35_XI0/XI51/XI3/MM10_d
+ N_XI0/XI51/XI3/NET36_XI0/XI51/XI3/MM10_g N_VDD_XI0/XI51/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI3/MM11 N_XI0/XI51/XI3/NET36_XI0/XI51/XI3/MM11_d
+ N_XI0/XI51/XI3/NET35_XI0/XI51/XI3/MM11_g N_VDD_XI0/XI51/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI4/MM2 N_XI0/XI51/XI4/NET34_XI0/XI51/XI4/MM2_d
+ N_XI0/XI51/XI4/NET33_XI0/XI51/XI4/MM2_g N_VSS_XI0/XI51/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM3 N_XI0/XI51/XI4/NET33_XI0/XI51/XI4/MM3_d
+ N_WL<98>_XI0/XI51/XI4/MM3_g N_BLN<11>_XI0/XI51/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM0 N_XI0/XI51/XI4/NET34_XI0/XI51/XI4/MM0_d
+ N_WL<98>_XI0/XI51/XI4/MM0_g N_BL<11>_XI0/XI51/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM1 N_XI0/XI51/XI4/NET33_XI0/XI51/XI4/MM1_d
+ N_XI0/XI51/XI4/NET34_XI0/XI51/XI4/MM1_g N_VSS_XI0/XI51/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM9 N_XI0/XI51/XI4/NET36_XI0/XI51/XI4/MM9_d
+ N_WL<99>_XI0/XI51/XI4/MM9_g N_BL<11>_XI0/XI51/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM6 N_XI0/XI51/XI4/NET35_XI0/XI51/XI4/MM6_d
+ N_XI0/XI51/XI4/NET36_XI0/XI51/XI4/MM6_g N_VSS_XI0/XI51/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM7 N_XI0/XI51/XI4/NET36_XI0/XI51/XI4/MM7_d
+ N_XI0/XI51/XI4/NET35_XI0/XI51/XI4/MM7_g N_VSS_XI0/XI51/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM8 N_XI0/XI51/XI4/NET35_XI0/XI51/XI4/MM8_d
+ N_WL<99>_XI0/XI51/XI4/MM8_g N_BLN<11>_XI0/XI51/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI4/MM5 N_XI0/XI51/XI4/NET34_XI0/XI51/XI4/MM5_d
+ N_XI0/XI51/XI4/NET33_XI0/XI51/XI4/MM5_g N_VDD_XI0/XI51/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI4/MM4 N_XI0/XI51/XI4/NET33_XI0/XI51/XI4/MM4_d
+ N_XI0/XI51/XI4/NET34_XI0/XI51/XI4/MM4_g N_VDD_XI0/XI51/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI4/MM10 N_XI0/XI51/XI4/NET35_XI0/XI51/XI4/MM10_d
+ N_XI0/XI51/XI4/NET36_XI0/XI51/XI4/MM10_g N_VDD_XI0/XI51/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI4/MM11 N_XI0/XI51/XI4/NET36_XI0/XI51/XI4/MM11_d
+ N_XI0/XI51/XI4/NET35_XI0/XI51/XI4/MM11_g N_VDD_XI0/XI51/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI5/MM2 N_XI0/XI51/XI5/NET34_XI0/XI51/XI5/MM2_d
+ N_XI0/XI51/XI5/NET33_XI0/XI51/XI5/MM2_g N_VSS_XI0/XI51/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM3 N_XI0/XI51/XI5/NET33_XI0/XI51/XI5/MM3_d
+ N_WL<98>_XI0/XI51/XI5/MM3_g N_BLN<10>_XI0/XI51/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM0 N_XI0/XI51/XI5/NET34_XI0/XI51/XI5/MM0_d
+ N_WL<98>_XI0/XI51/XI5/MM0_g N_BL<10>_XI0/XI51/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM1 N_XI0/XI51/XI5/NET33_XI0/XI51/XI5/MM1_d
+ N_XI0/XI51/XI5/NET34_XI0/XI51/XI5/MM1_g N_VSS_XI0/XI51/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM9 N_XI0/XI51/XI5/NET36_XI0/XI51/XI5/MM9_d
+ N_WL<99>_XI0/XI51/XI5/MM9_g N_BL<10>_XI0/XI51/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM6 N_XI0/XI51/XI5/NET35_XI0/XI51/XI5/MM6_d
+ N_XI0/XI51/XI5/NET36_XI0/XI51/XI5/MM6_g N_VSS_XI0/XI51/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM7 N_XI0/XI51/XI5/NET36_XI0/XI51/XI5/MM7_d
+ N_XI0/XI51/XI5/NET35_XI0/XI51/XI5/MM7_g N_VSS_XI0/XI51/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM8 N_XI0/XI51/XI5/NET35_XI0/XI51/XI5/MM8_d
+ N_WL<99>_XI0/XI51/XI5/MM8_g N_BLN<10>_XI0/XI51/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI5/MM5 N_XI0/XI51/XI5/NET34_XI0/XI51/XI5/MM5_d
+ N_XI0/XI51/XI5/NET33_XI0/XI51/XI5/MM5_g N_VDD_XI0/XI51/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI5/MM4 N_XI0/XI51/XI5/NET33_XI0/XI51/XI5/MM4_d
+ N_XI0/XI51/XI5/NET34_XI0/XI51/XI5/MM4_g N_VDD_XI0/XI51/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI5/MM10 N_XI0/XI51/XI5/NET35_XI0/XI51/XI5/MM10_d
+ N_XI0/XI51/XI5/NET36_XI0/XI51/XI5/MM10_g N_VDD_XI0/XI51/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI5/MM11 N_XI0/XI51/XI5/NET36_XI0/XI51/XI5/MM11_d
+ N_XI0/XI51/XI5/NET35_XI0/XI51/XI5/MM11_g N_VDD_XI0/XI51/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI6/MM2 N_XI0/XI51/XI6/NET34_XI0/XI51/XI6/MM2_d
+ N_XI0/XI51/XI6/NET33_XI0/XI51/XI6/MM2_g N_VSS_XI0/XI51/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM3 N_XI0/XI51/XI6/NET33_XI0/XI51/XI6/MM3_d
+ N_WL<98>_XI0/XI51/XI6/MM3_g N_BLN<9>_XI0/XI51/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM0 N_XI0/XI51/XI6/NET34_XI0/XI51/XI6/MM0_d
+ N_WL<98>_XI0/XI51/XI6/MM0_g N_BL<9>_XI0/XI51/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM1 N_XI0/XI51/XI6/NET33_XI0/XI51/XI6/MM1_d
+ N_XI0/XI51/XI6/NET34_XI0/XI51/XI6/MM1_g N_VSS_XI0/XI51/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM9 N_XI0/XI51/XI6/NET36_XI0/XI51/XI6/MM9_d
+ N_WL<99>_XI0/XI51/XI6/MM9_g N_BL<9>_XI0/XI51/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM6 N_XI0/XI51/XI6/NET35_XI0/XI51/XI6/MM6_d
+ N_XI0/XI51/XI6/NET36_XI0/XI51/XI6/MM6_g N_VSS_XI0/XI51/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM7 N_XI0/XI51/XI6/NET36_XI0/XI51/XI6/MM7_d
+ N_XI0/XI51/XI6/NET35_XI0/XI51/XI6/MM7_g N_VSS_XI0/XI51/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM8 N_XI0/XI51/XI6/NET35_XI0/XI51/XI6/MM8_d
+ N_WL<99>_XI0/XI51/XI6/MM8_g N_BLN<9>_XI0/XI51/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI6/MM5 N_XI0/XI51/XI6/NET34_XI0/XI51/XI6/MM5_d
+ N_XI0/XI51/XI6/NET33_XI0/XI51/XI6/MM5_g N_VDD_XI0/XI51/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI6/MM4 N_XI0/XI51/XI6/NET33_XI0/XI51/XI6/MM4_d
+ N_XI0/XI51/XI6/NET34_XI0/XI51/XI6/MM4_g N_VDD_XI0/XI51/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI6/MM10 N_XI0/XI51/XI6/NET35_XI0/XI51/XI6/MM10_d
+ N_XI0/XI51/XI6/NET36_XI0/XI51/XI6/MM10_g N_VDD_XI0/XI51/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI6/MM11 N_XI0/XI51/XI6/NET36_XI0/XI51/XI6/MM11_d
+ N_XI0/XI51/XI6/NET35_XI0/XI51/XI6/MM11_g N_VDD_XI0/XI51/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI7/MM2 N_XI0/XI51/XI7/NET34_XI0/XI51/XI7/MM2_d
+ N_XI0/XI51/XI7/NET33_XI0/XI51/XI7/MM2_g N_VSS_XI0/XI51/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM3 N_XI0/XI51/XI7/NET33_XI0/XI51/XI7/MM3_d
+ N_WL<98>_XI0/XI51/XI7/MM3_g N_BLN<8>_XI0/XI51/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM0 N_XI0/XI51/XI7/NET34_XI0/XI51/XI7/MM0_d
+ N_WL<98>_XI0/XI51/XI7/MM0_g N_BL<8>_XI0/XI51/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM1 N_XI0/XI51/XI7/NET33_XI0/XI51/XI7/MM1_d
+ N_XI0/XI51/XI7/NET34_XI0/XI51/XI7/MM1_g N_VSS_XI0/XI51/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM9 N_XI0/XI51/XI7/NET36_XI0/XI51/XI7/MM9_d
+ N_WL<99>_XI0/XI51/XI7/MM9_g N_BL<8>_XI0/XI51/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM6 N_XI0/XI51/XI7/NET35_XI0/XI51/XI7/MM6_d
+ N_XI0/XI51/XI7/NET36_XI0/XI51/XI7/MM6_g N_VSS_XI0/XI51/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM7 N_XI0/XI51/XI7/NET36_XI0/XI51/XI7/MM7_d
+ N_XI0/XI51/XI7/NET35_XI0/XI51/XI7/MM7_g N_VSS_XI0/XI51/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM8 N_XI0/XI51/XI7/NET35_XI0/XI51/XI7/MM8_d
+ N_WL<99>_XI0/XI51/XI7/MM8_g N_BLN<8>_XI0/XI51/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI7/MM5 N_XI0/XI51/XI7/NET34_XI0/XI51/XI7/MM5_d
+ N_XI0/XI51/XI7/NET33_XI0/XI51/XI7/MM5_g N_VDD_XI0/XI51/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI7/MM4 N_XI0/XI51/XI7/NET33_XI0/XI51/XI7/MM4_d
+ N_XI0/XI51/XI7/NET34_XI0/XI51/XI7/MM4_g N_VDD_XI0/XI51/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI7/MM10 N_XI0/XI51/XI7/NET35_XI0/XI51/XI7/MM10_d
+ N_XI0/XI51/XI7/NET36_XI0/XI51/XI7/MM10_g N_VDD_XI0/XI51/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI7/MM11 N_XI0/XI51/XI7/NET36_XI0/XI51/XI7/MM11_d
+ N_XI0/XI51/XI7/NET35_XI0/XI51/XI7/MM11_g N_VDD_XI0/XI51/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI8/MM2 N_XI0/XI51/XI8/NET34_XI0/XI51/XI8/MM2_d
+ N_XI0/XI51/XI8/NET33_XI0/XI51/XI8/MM2_g N_VSS_XI0/XI51/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM3 N_XI0/XI51/XI8/NET33_XI0/XI51/XI8/MM3_d
+ N_WL<98>_XI0/XI51/XI8/MM3_g N_BLN<7>_XI0/XI51/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM0 N_XI0/XI51/XI8/NET34_XI0/XI51/XI8/MM0_d
+ N_WL<98>_XI0/XI51/XI8/MM0_g N_BL<7>_XI0/XI51/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM1 N_XI0/XI51/XI8/NET33_XI0/XI51/XI8/MM1_d
+ N_XI0/XI51/XI8/NET34_XI0/XI51/XI8/MM1_g N_VSS_XI0/XI51/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM9 N_XI0/XI51/XI8/NET36_XI0/XI51/XI8/MM9_d
+ N_WL<99>_XI0/XI51/XI8/MM9_g N_BL<7>_XI0/XI51/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM6 N_XI0/XI51/XI8/NET35_XI0/XI51/XI8/MM6_d
+ N_XI0/XI51/XI8/NET36_XI0/XI51/XI8/MM6_g N_VSS_XI0/XI51/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM7 N_XI0/XI51/XI8/NET36_XI0/XI51/XI8/MM7_d
+ N_XI0/XI51/XI8/NET35_XI0/XI51/XI8/MM7_g N_VSS_XI0/XI51/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM8 N_XI0/XI51/XI8/NET35_XI0/XI51/XI8/MM8_d
+ N_WL<99>_XI0/XI51/XI8/MM8_g N_BLN<7>_XI0/XI51/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI8/MM5 N_XI0/XI51/XI8/NET34_XI0/XI51/XI8/MM5_d
+ N_XI0/XI51/XI8/NET33_XI0/XI51/XI8/MM5_g N_VDD_XI0/XI51/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI8/MM4 N_XI0/XI51/XI8/NET33_XI0/XI51/XI8/MM4_d
+ N_XI0/XI51/XI8/NET34_XI0/XI51/XI8/MM4_g N_VDD_XI0/XI51/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI8/MM10 N_XI0/XI51/XI8/NET35_XI0/XI51/XI8/MM10_d
+ N_XI0/XI51/XI8/NET36_XI0/XI51/XI8/MM10_g N_VDD_XI0/XI51/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI8/MM11 N_XI0/XI51/XI8/NET36_XI0/XI51/XI8/MM11_d
+ N_XI0/XI51/XI8/NET35_XI0/XI51/XI8/MM11_g N_VDD_XI0/XI51/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI9/MM2 N_XI0/XI51/XI9/NET34_XI0/XI51/XI9/MM2_d
+ N_XI0/XI51/XI9/NET33_XI0/XI51/XI9/MM2_g N_VSS_XI0/XI51/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM3 N_XI0/XI51/XI9/NET33_XI0/XI51/XI9/MM3_d
+ N_WL<98>_XI0/XI51/XI9/MM3_g N_BLN<6>_XI0/XI51/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM0 N_XI0/XI51/XI9/NET34_XI0/XI51/XI9/MM0_d
+ N_WL<98>_XI0/XI51/XI9/MM0_g N_BL<6>_XI0/XI51/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM1 N_XI0/XI51/XI9/NET33_XI0/XI51/XI9/MM1_d
+ N_XI0/XI51/XI9/NET34_XI0/XI51/XI9/MM1_g N_VSS_XI0/XI51/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM9 N_XI0/XI51/XI9/NET36_XI0/XI51/XI9/MM9_d
+ N_WL<99>_XI0/XI51/XI9/MM9_g N_BL<6>_XI0/XI51/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM6 N_XI0/XI51/XI9/NET35_XI0/XI51/XI9/MM6_d
+ N_XI0/XI51/XI9/NET36_XI0/XI51/XI9/MM6_g N_VSS_XI0/XI51/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM7 N_XI0/XI51/XI9/NET36_XI0/XI51/XI9/MM7_d
+ N_XI0/XI51/XI9/NET35_XI0/XI51/XI9/MM7_g N_VSS_XI0/XI51/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM8 N_XI0/XI51/XI9/NET35_XI0/XI51/XI9/MM8_d
+ N_WL<99>_XI0/XI51/XI9/MM8_g N_BLN<6>_XI0/XI51/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI9/MM5 N_XI0/XI51/XI9/NET34_XI0/XI51/XI9/MM5_d
+ N_XI0/XI51/XI9/NET33_XI0/XI51/XI9/MM5_g N_VDD_XI0/XI51/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI9/MM4 N_XI0/XI51/XI9/NET33_XI0/XI51/XI9/MM4_d
+ N_XI0/XI51/XI9/NET34_XI0/XI51/XI9/MM4_g N_VDD_XI0/XI51/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI9/MM10 N_XI0/XI51/XI9/NET35_XI0/XI51/XI9/MM10_d
+ N_XI0/XI51/XI9/NET36_XI0/XI51/XI9/MM10_g N_VDD_XI0/XI51/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI9/MM11 N_XI0/XI51/XI9/NET36_XI0/XI51/XI9/MM11_d
+ N_XI0/XI51/XI9/NET35_XI0/XI51/XI9/MM11_g N_VDD_XI0/XI51/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI10/MM2 N_XI0/XI51/XI10/NET34_XI0/XI51/XI10/MM2_d
+ N_XI0/XI51/XI10/NET33_XI0/XI51/XI10/MM2_g N_VSS_XI0/XI51/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM3 N_XI0/XI51/XI10/NET33_XI0/XI51/XI10/MM3_d
+ N_WL<98>_XI0/XI51/XI10/MM3_g N_BLN<5>_XI0/XI51/XI10/MM3_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM0 N_XI0/XI51/XI10/NET34_XI0/XI51/XI10/MM0_d
+ N_WL<98>_XI0/XI51/XI10/MM0_g N_BL<5>_XI0/XI51/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM1 N_XI0/XI51/XI10/NET33_XI0/XI51/XI10/MM1_d
+ N_XI0/XI51/XI10/NET34_XI0/XI51/XI10/MM1_g N_VSS_XI0/XI51/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM9 N_XI0/XI51/XI10/NET36_XI0/XI51/XI10/MM9_d
+ N_WL<99>_XI0/XI51/XI10/MM9_g N_BL<5>_XI0/XI51/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM6 N_XI0/XI51/XI10/NET35_XI0/XI51/XI10/MM6_d
+ N_XI0/XI51/XI10/NET36_XI0/XI51/XI10/MM6_g N_VSS_XI0/XI51/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM7 N_XI0/XI51/XI10/NET36_XI0/XI51/XI10/MM7_d
+ N_XI0/XI51/XI10/NET35_XI0/XI51/XI10/MM7_g N_VSS_XI0/XI51/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM8 N_XI0/XI51/XI10/NET35_XI0/XI51/XI10/MM8_d
+ N_WL<99>_XI0/XI51/XI10/MM8_g N_BLN<5>_XI0/XI51/XI10/MM8_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI10/MM5 N_XI0/XI51/XI10/NET34_XI0/XI51/XI10/MM5_d
+ N_XI0/XI51/XI10/NET33_XI0/XI51/XI10/MM5_g N_VDD_XI0/XI51/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI10/MM4 N_XI0/XI51/XI10/NET33_XI0/XI51/XI10/MM4_d
+ N_XI0/XI51/XI10/NET34_XI0/XI51/XI10/MM4_g N_VDD_XI0/XI51/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI10/MM10 N_XI0/XI51/XI10/NET35_XI0/XI51/XI10/MM10_d
+ N_XI0/XI51/XI10/NET36_XI0/XI51/XI10/MM10_g N_VDD_XI0/XI51/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI10/MM11 N_XI0/XI51/XI10/NET36_XI0/XI51/XI10/MM11_d
+ N_XI0/XI51/XI10/NET35_XI0/XI51/XI10/MM11_g N_VDD_XI0/XI51/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI11/MM2 N_XI0/XI51/XI11/NET34_XI0/XI51/XI11/MM2_d
+ N_XI0/XI51/XI11/NET33_XI0/XI51/XI11/MM2_g N_VSS_XI0/XI51/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM3 N_XI0/XI51/XI11/NET33_XI0/XI51/XI11/MM3_d
+ N_WL<98>_XI0/XI51/XI11/MM3_g N_BLN<4>_XI0/XI51/XI11/MM3_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM0 N_XI0/XI51/XI11/NET34_XI0/XI51/XI11/MM0_d
+ N_WL<98>_XI0/XI51/XI11/MM0_g N_BL<4>_XI0/XI51/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM1 N_XI0/XI51/XI11/NET33_XI0/XI51/XI11/MM1_d
+ N_XI0/XI51/XI11/NET34_XI0/XI51/XI11/MM1_g N_VSS_XI0/XI51/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM9 N_XI0/XI51/XI11/NET36_XI0/XI51/XI11/MM9_d
+ N_WL<99>_XI0/XI51/XI11/MM9_g N_BL<4>_XI0/XI51/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM6 N_XI0/XI51/XI11/NET35_XI0/XI51/XI11/MM6_d
+ N_XI0/XI51/XI11/NET36_XI0/XI51/XI11/MM6_g N_VSS_XI0/XI51/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM7 N_XI0/XI51/XI11/NET36_XI0/XI51/XI11/MM7_d
+ N_XI0/XI51/XI11/NET35_XI0/XI51/XI11/MM7_g N_VSS_XI0/XI51/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM8 N_XI0/XI51/XI11/NET35_XI0/XI51/XI11/MM8_d
+ N_WL<99>_XI0/XI51/XI11/MM8_g N_BLN<4>_XI0/XI51/XI11/MM8_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI11/MM5 N_XI0/XI51/XI11/NET34_XI0/XI51/XI11/MM5_d
+ N_XI0/XI51/XI11/NET33_XI0/XI51/XI11/MM5_g N_VDD_XI0/XI51/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI11/MM4 N_XI0/XI51/XI11/NET33_XI0/XI51/XI11/MM4_d
+ N_XI0/XI51/XI11/NET34_XI0/XI51/XI11/MM4_g N_VDD_XI0/XI51/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI11/MM10 N_XI0/XI51/XI11/NET35_XI0/XI51/XI11/MM10_d
+ N_XI0/XI51/XI11/NET36_XI0/XI51/XI11/MM10_g N_VDD_XI0/XI51/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI11/MM11 N_XI0/XI51/XI11/NET36_XI0/XI51/XI11/MM11_d
+ N_XI0/XI51/XI11/NET35_XI0/XI51/XI11/MM11_g N_VDD_XI0/XI51/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI12/MM2 N_XI0/XI51/XI12/NET34_XI0/XI51/XI12/MM2_d
+ N_XI0/XI51/XI12/NET33_XI0/XI51/XI12/MM2_g N_VSS_XI0/XI51/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM3 N_XI0/XI51/XI12/NET33_XI0/XI51/XI12/MM3_d
+ N_WL<98>_XI0/XI51/XI12/MM3_g N_BLN<3>_XI0/XI51/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM0 N_XI0/XI51/XI12/NET34_XI0/XI51/XI12/MM0_d
+ N_WL<98>_XI0/XI51/XI12/MM0_g N_BL<3>_XI0/XI51/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM1 N_XI0/XI51/XI12/NET33_XI0/XI51/XI12/MM1_d
+ N_XI0/XI51/XI12/NET34_XI0/XI51/XI12/MM1_g N_VSS_XI0/XI51/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM9 N_XI0/XI51/XI12/NET36_XI0/XI51/XI12/MM9_d
+ N_WL<99>_XI0/XI51/XI12/MM9_g N_BL<3>_XI0/XI51/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM6 N_XI0/XI51/XI12/NET35_XI0/XI51/XI12/MM6_d
+ N_XI0/XI51/XI12/NET36_XI0/XI51/XI12/MM6_g N_VSS_XI0/XI51/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM7 N_XI0/XI51/XI12/NET36_XI0/XI51/XI12/MM7_d
+ N_XI0/XI51/XI12/NET35_XI0/XI51/XI12/MM7_g N_VSS_XI0/XI51/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM8 N_XI0/XI51/XI12/NET35_XI0/XI51/XI12/MM8_d
+ N_WL<99>_XI0/XI51/XI12/MM8_g N_BLN<3>_XI0/XI51/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI12/MM5 N_XI0/XI51/XI12/NET34_XI0/XI51/XI12/MM5_d
+ N_XI0/XI51/XI12/NET33_XI0/XI51/XI12/MM5_g N_VDD_XI0/XI51/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI12/MM4 N_XI0/XI51/XI12/NET33_XI0/XI51/XI12/MM4_d
+ N_XI0/XI51/XI12/NET34_XI0/XI51/XI12/MM4_g N_VDD_XI0/XI51/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI12/MM10 N_XI0/XI51/XI12/NET35_XI0/XI51/XI12/MM10_d
+ N_XI0/XI51/XI12/NET36_XI0/XI51/XI12/MM10_g N_VDD_XI0/XI51/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI12/MM11 N_XI0/XI51/XI12/NET36_XI0/XI51/XI12/MM11_d
+ N_XI0/XI51/XI12/NET35_XI0/XI51/XI12/MM11_g N_VDD_XI0/XI51/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI13/MM2 N_XI0/XI51/XI13/NET34_XI0/XI51/XI13/MM2_d
+ N_XI0/XI51/XI13/NET33_XI0/XI51/XI13/MM2_g N_VSS_XI0/XI51/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM3 N_XI0/XI51/XI13/NET33_XI0/XI51/XI13/MM3_d
+ N_WL<98>_XI0/XI51/XI13/MM3_g N_BLN<2>_XI0/XI51/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM0 N_XI0/XI51/XI13/NET34_XI0/XI51/XI13/MM0_d
+ N_WL<98>_XI0/XI51/XI13/MM0_g N_BL<2>_XI0/XI51/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM1 N_XI0/XI51/XI13/NET33_XI0/XI51/XI13/MM1_d
+ N_XI0/XI51/XI13/NET34_XI0/XI51/XI13/MM1_g N_VSS_XI0/XI51/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM9 N_XI0/XI51/XI13/NET36_XI0/XI51/XI13/MM9_d
+ N_WL<99>_XI0/XI51/XI13/MM9_g N_BL<2>_XI0/XI51/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM6 N_XI0/XI51/XI13/NET35_XI0/XI51/XI13/MM6_d
+ N_XI0/XI51/XI13/NET36_XI0/XI51/XI13/MM6_g N_VSS_XI0/XI51/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM7 N_XI0/XI51/XI13/NET36_XI0/XI51/XI13/MM7_d
+ N_XI0/XI51/XI13/NET35_XI0/XI51/XI13/MM7_g N_VSS_XI0/XI51/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM8 N_XI0/XI51/XI13/NET35_XI0/XI51/XI13/MM8_d
+ N_WL<99>_XI0/XI51/XI13/MM8_g N_BLN<2>_XI0/XI51/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI13/MM5 N_XI0/XI51/XI13/NET34_XI0/XI51/XI13/MM5_d
+ N_XI0/XI51/XI13/NET33_XI0/XI51/XI13/MM5_g N_VDD_XI0/XI51/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI13/MM4 N_XI0/XI51/XI13/NET33_XI0/XI51/XI13/MM4_d
+ N_XI0/XI51/XI13/NET34_XI0/XI51/XI13/MM4_g N_VDD_XI0/XI51/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI13/MM10 N_XI0/XI51/XI13/NET35_XI0/XI51/XI13/MM10_d
+ N_XI0/XI51/XI13/NET36_XI0/XI51/XI13/MM10_g N_VDD_XI0/XI51/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI13/MM11 N_XI0/XI51/XI13/NET36_XI0/XI51/XI13/MM11_d
+ N_XI0/XI51/XI13/NET35_XI0/XI51/XI13/MM11_g N_VDD_XI0/XI51/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI14/MM2 N_XI0/XI51/XI14/NET34_XI0/XI51/XI14/MM2_d
+ N_XI0/XI51/XI14/NET33_XI0/XI51/XI14/MM2_g N_VSS_XI0/XI51/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM3 N_XI0/XI51/XI14/NET33_XI0/XI51/XI14/MM3_d
+ N_WL<98>_XI0/XI51/XI14/MM3_g N_BLN<1>_XI0/XI51/XI14/MM3_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM0 N_XI0/XI51/XI14/NET34_XI0/XI51/XI14/MM0_d
+ N_WL<98>_XI0/XI51/XI14/MM0_g N_BL<1>_XI0/XI51/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM1 N_XI0/XI51/XI14/NET33_XI0/XI51/XI14/MM1_d
+ N_XI0/XI51/XI14/NET34_XI0/XI51/XI14/MM1_g N_VSS_XI0/XI51/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM9 N_XI0/XI51/XI14/NET36_XI0/XI51/XI14/MM9_d
+ N_WL<99>_XI0/XI51/XI14/MM9_g N_BL<1>_XI0/XI51/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM6 N_XI0/XI51/XI14/NET35_XI0/XI51/XI14/MM6_d
+ N_XI0/XI51/XI14/NET36_XI0/XI51/XI14/MM6_g N_VSS_XI0/XI51/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM7 N_XI0/XI51/XI14/NET36_XI0/XI51/XI14/MM7_d
+ N_XI0/XI51/XI14/NET35_XI0/XI51/XI14/MM7_g N_VSS_XI0/XI51/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM8 N_XI0/XI51/XI14/NET35_XI0/XI51/XI14/MM8_d
+ N_WL<99>_XI0/XI51/XI14/MM8_g N_BLN<1>_XI0/XI51/XI14/MM8_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI14/MM5 N_XI0/XI51/XI14/NET34_XI0/XI51/XI14/MM5_d
+ N_XI0/XI51/XI14/NET33_XI0/XI51/XI14/MM5_g N_VDD_XI0/XI51/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI14/MM4 N_XI0/XI51/XI14/NET33_XI0/XI51/XI14/MM4_d
+ N_XI0/XI51/XI14/NET34_XI0/XI51/XI14/MM4_g N_VDD_XI0/XI51/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI14/MM10 N_XI0/XI51/XI14/NET35_XI0/XI51/XI14/MM10_d
+ N_XI0/XI51/XI14/NET36_XI0/XI51/XI14/MM10_g N_VDD_XI0/XI51/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI14/MM11 N_XI0/XI51/XI14/NET36_XI0/XI51/XI14/MM11_d
+ N_XI0/XI51/XI14/NET35_XI0/XI51/XI14/MM11_g N_VDD_XI0/XI51/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI15/MM2 N_XI0/XI51/XI15/NET34_XI0/XI51/XI15/MM2_d
+ N_XI0/XI51/XI15/NET33_XI0/XI51/XI15/MM2_g N_VSS_XI0/XI51/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM3 N_XI0/XI51/XI15/NET33_XI0/XI51/XI15/MM3_d
+ N_WL<98>_XI0/XI51/XI15/MM3_g N_BLN<0>_XI0/XI51/XI15/MM3_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM0 N_XI0/XI51/XI15/NET34_XI0/XI51/XI15/MM0_d
+ N_WL<98>_XI0/XI51/XI15/MM0_g N_BL<0>_XI0/XI51/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM1 N_XI0/XI51/XI15/NET33_XI0/XI51/XI15/MM1_d
+ N_XI0/XI51/XI15/NET34_XI0/XI51/XI15/MM1_g N_VSS_XI0/XI51/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM9 N_XI0/XI51/XI15/NET36_XI0/XI51/XI15/MM9_d
+ N_WL<99>_XI0/XI51/XI15/MM9_g N_BL<0>_XI0/XI51/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM6 N_XI0/XI51/XI15/NET35_XI0/XI51/XI15/MM6_d
+ N_XI0/XI51/XI15/NET36_XI0/XI51/XI15/MM6_g N_VSS_XI0/XI51/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM7 N_XI0/XI51/XI15/NET36_XI0/XI51/XI15/MM7_d
+ N_XI0/XI51/XI15/NET35_XI0/XI51/XI15/MM7_g N_VSS_XI0/XI51/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM8 N_XI0/XI51/XI15/NET35_XI0/XI51/XI15/MM8_d
+ N_WL<99>_XI0/XI51/XI15/MM8_g N_BLN<0>_XI0/XI51/XI15/MM8_s N_VSS_XI1/XI15/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI51/XI15/MM5 N_XI0/XI51/XI15/NET34_XI0/XI51/XI15/MM5_d
+ N_XI0/XI51/XI15/NET33_XI0/XI51/XI15/MM5_g N_VDD_XI0/XI51/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI15/MM4 N_XI0/XI51/XI15/NET33_XI0/XI51/XI15/MM4_d
+ N_XI0/XI51/XI15/NET34_XI0/XI51/XI15/MM4_g N_VDD_XI0/XI51/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI15/MM10 N_XI0/XI51/XI15/NET35_XI0/XI51/XI15/MM10_d
+ N_XI0/XI51/XI15/NET36_XI0/XI51/XI15/MM10_g N_VDD_XI0/XI51/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI51/XI15/MM11 N_XI0/XI51/XI15/NET36_XI0/XI51/XI15/MM11_d
+ N_XI0/XI51/XI15/NET35_XI0/XI51/XI15/MM11_g N_VDD_XI0/XI51/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI0/MM2 N_XI0/XI52/XI0/NET34_XI0/XI52/XI0/MM2_d
+ N_XI0/XI52/XI0/NET33_XI0/XI52/XI0/MM2_g N_VSS_XI0/XI52/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM3 N_XI0/XI52/XI0/NET33_XI0/XI52/XI0/MM3_d
+ N_WL<100>_XI0/XI52/XI0/MM3_g N_BLN<15>_XI0/XI52/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM0 N_XI0/XI52/XI0/NET34_XI0/XI52/XI0/MM0_d
+ N_WL<100>_XI0/XI52/XI0/MM0_g N_BL<15>_XI0/XI52/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM1 N_XI0/XI52/XI0/NET33_XI0/XI52/XI0/MM1_d
+ N_XI0/XI52/XI0/NET34_XI0/XI52/XI0/MM1_g N_VSS_XI0/XI52/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM9 N_XI0/XI52/XI0/NET36_XI0/XI52/XI0/MM9_d
+ N_WL<101>_XI0/XI52/XI0/MM9_g N_BL<15>_XI0/XI52/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM6 N_XI0/XI52/XI0/NET35_XI0/XI52/XI0/MM6_d
+ N_XI0/XI52/XI0/NET36_XI0/XI52/XI0/MM6_g N_VSS_XI0/XI52/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM7 N_XI0/XI52/XI0/NET36_XI0/XI52/XI0/MM7_d
+ N_XI0/XI52/XI0/NET35_XI0/XI52/XI0/MM7_g N_VSS_XI0/XI52/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM8 N_XI0/XI52/XI0/NET35_XI0/XI52/XI0/MM8_d
+ N_WL<101>_XI0/XI52/XI0/MM8_g N_BLN<15>_XI0/XI52/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI0/MM5 N_XI0/XI52/XI0/NET34_XI0/XI52/XI0/MM5_d
+ N_XI0/XI52/XI0/NET33_XI0/XI52/XI0/MM5_g N_VDD_XI0/XI52/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI0/MM4 N_XI0/XI52/XI0/NET33_XI0/XI52/XI0/MM4_d
+ N_XI0/XI52/XI0/NET34_XI0/XI52/XI0/MM4_g N_VDD_XI0/XI52/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI0/MM10 N_XI0/XI52/XI0/NET35_XI0/XI52/XI0/MM10_d
+ N_XI0/XI52/XI0/NET36_XI0/XI52/XI0/MM10_g N_VDD_XI0/XI52/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI0/MM11 N_XI0/XI52/XI0/NET36_XI0/XI52/XI0/MM11_d
+ N_XI0/XI52/XI0/NET35_XI0/XI52/XI0/MM11_g N_VDD_XI0/XI52/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI1/MM2 N_XI0/XI52/XI1/NET34_XI0/XI52/XI1/MM2_d
+ N_XI0/XI52/XI1/NET33_XI0/XI52/XI1/MM2_g N_VSS_XI0/XI52/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM3 N_XI0/XI52/XI1/NET33_XI0/XI52/XI1/MM3_d
+ N_WL<100>_XI0/XI52/XI1/MM3_g N_BLN<14>_XI0/XI52/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM0 N_XI0/XI52/XI1/NET34_XI0/XI52/XI1/MM0_d
+ N_WL<100>_XI0/XI52/XI1/MM0_g N_BL<14>_XI0/XI52/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM1 N_XI0/XI52/XI1/NET33_XI0/XI52/XI1/MM1_d
+ N_XI0/XI52/XI1/NET34_XI0/XI52/XI1/MM1_g N_VSS_XI0/XI52/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM9 N_XI0/XI52/XI1/NET36_XI0/XI52/XI1/MM9_d
+ N_WL<101>_XI0/XI52/XI1/MM9_g N_BL<14>_XI0/XI52/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM6 N_XI0/XI52/XI1/NET35_XI0/XI52/XI1/MM6_d
+ N_XI0/XI52/XI1/NET36_XI0/XI52/XI1/MM6_g N_VSS_XI0/XI52/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM7 N_XI0/XI52/XI1/NET36_XI0/XI52/XI1/MM7_d
+ N_XI0/XI52/XI1/NET35_XI0/XI52/XI1/MM7_g N_VSS_XI0/XI52/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM8 N_XI0/XI52/XI1/NET35_XI0/XI52/XI1/MM8_d
+ N_WL<101>_XI0/XI52/XI1/MM8_g N_BLN<14>_XI0/XI52/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI1/MM5 N_XI0/XI52/XI1/NET34_XI0/XI52/XI1/MM5_d
+ N_XI0/XI52/XI1/NET33_XI0/XI52/XI1/MM5_g N_VDD_XI0/XI52/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI1/MM4 N_XI0/XI52/XI1/NET33_XI0/XI52/XI1/MM4_d
+ N_XI0/XI52/XI1/NET34_XI0/XI52/XI1/MM4_g N_VDD_XI0/XI52/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI1/MM10 N_XI0/XI52/XI1/NET35_XI0/XI52/XI1/MM10_d
+ N_XI0/XI52/XI1/NET36_XI0/XI52/XI1/MM10_g N_VDD_XI0/XI52/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI1/MM11 N_XI0/XI52/XI1/NET36_XI0/XI52/XI1/MM11_d
+ N_XI0/XI52/XI1/NET35_XI0/XI52/XI1/MM11_g N_VDD_XI0/XI52/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI2/MM2 N_XI0/XI52/XI2/NET34_XI0/XI52/XI2/MM2_d
+ N_XI0/XI52/XI2/NET33_XI0/XI52/XI2/MM2_g N_VSS_XI0/XI52/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM3 N_XI0/XI52/XI2/NET33_XI0/XI52/XI2/MM3_d
+ N_WL<100>_XI0/XI52/XI2/MM3_g N_BLN<13>_XI0/XI52/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM0 N_XI0/XI52/XI2/NET34_XI0/XI52/XI2/MM0_d
+ N_WL<100>_XI0/XI52/XI2/MM0_g N_BL<13>_XI0/XI52/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM1 N_XI0/XI52/XI2/NET33_XI0/XI52/XI2/MM1_d
+ N_XI0/XI52/XI2/NET34_XI0/XI52/XI2/MM1_g N_VSS_XI0/XI52/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM9 N_XI0/XI52/XI2/NET36_XI0/XI52/XI2/MM9_d
+ N_WL<101>_XI0/XI52/XI2/MM9_g N_BL<13>_XI0/XI52/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM6 N_XI0/XI52/XI2/NET35_XI0/XI52/XI2/MM6_d
+ N_XI0/XI52/XI2/NET36_XI0/XI52/XI2/MM6_g N_VSS_XI0/XI52/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM7 N_XI0/XI52/XI2/NET36_XI0/XI52/XI2/MM7_d
+ N_XI0/XI52/XI2/NET35_XI0/XI52/XI2/MM7_g N_VSS_XI0/XI52/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM8 N_XI0/XI52/XI2/NET35_XI0/XI52/XI2/MM8_d
+ N_WL<101>_XI0/XI52/XI2/MM8_g N_BLN<13>_XI0/XI52/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI2/MM5 N_XI0/XI52/XI2/NET34_XI0/XI52/XI2/MM5_d
+ N_XI0/XI52/XI2/NET33_XI0/XI52/XI2/MM5_g N_VDD_XI0/XI52/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI2/MM4 N_XI0/XI52/XI2/NET33_XI0/XI52/XI2/MM4_d
+ N_XI0/XI52/XI2/NET34_XI0/XI52/XI2/MM4_g N_VDD_XI0/XI52/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI2/MM10 N_XI0/XI52/XI2/NET35_XI0/XI52/XI2/MM10_d
+ N_XI0/XI52/XI2/NET36_XI0/XI52/XI2/MM10_g N_VDD_XI0/XI52/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI2/MM11 N_XI0/XI52/XI2/NET36_XI0/XI52/XI2/MM11_d
+ N_XI0/XI52/XI2/NET35_XI0/XI52/XI2/MM11_g N_VDD_XI0/XI52/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI3/MM2 N_XI0/XI52/XI3/NET34_XI0/XI52/XI3/MM2_d
+ N_XI0/XI52/XI3/NET33_XI0/XI52/XI3/MM2_g N_VSS_XI0/XI52/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM3 N_XI0/XI52/XI3/NET33_XI0/XI52/XI3/MM3_d
+ N_WL<100>_XI0/XI52/XI3/MM3_g N_BLN<12>_XI0/XI52/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM0 N_XI0/XI52/XI3/NET34_XI0/XI52/XI3/MM0_d
+ N_WL<100>_XI0/XI52/XI3/MM0_g N_BL<12>_XI0/XI52/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM1 N_XI0/XI52/XI3/NET33_XI0/XI52/XI3/MM1_d
+ N_XI0/XI52/XI3/NET34_XI0/XI52/XI3/MM1_g N_VSS_XI0/XI52/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM9 N_XI0/XI52/XI3/NET36_XI0/XI52/XI3/MM9_d
+ N_WL<101>_XI0/XI52/XI3/MM9_g N_BL<12>_XI0/XI52/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM6 N_XI0/XI52/XI3/NET35_XI0/XI52/XI3/MM6_d
+ N_XI0/XI52/XI3/NET36_XI0/XI52/XI3/MM6_g N_VSS_XI0/XI52/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM7 N_XI0/XI52/XI3/NET36_XI0/XI52/XI3/MM7_d
+ N_XI0/XI52/XI3/NET35_XI0/XI52/XI3/MM7_g N_VSS_XI0/XI52/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM8 N_XI0/XI52/XI3/NET35_XI0/XI52/XI3/MM8_d
+ N_WL<101>_XI0/XI52/XI3/MM8_g N_BLN<12>_XI0/XI52/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI3/MM5 N_XI0/XI52/XI3/NET34_XI0/XI52/XI3/MM5_d
+ N_XI0/XI52/XI3/NET33_XI0/XI52/XI3/MM5_g N_VDD_XI0/XI52/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI3/MM4 N_XI0/XI52/XI3/NET33_XI0/XI52/XI3/MM4_d
+ N_XI0/XI52/XI3/NET34_XI0/XI52/XI3/MM4_g N_VDD_XI0/XI52/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI3/MM10 N_XI0/XI52/XI3/NET35_XI0/XI52/XI3/MM10_d
+ N_XI0/XI52/XI3/NET36_XI0/XI52/XI3/MM10_g N_VDD_XI0/XI52/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI3/MM11 N_XI0/XI52/XI3/NET36_XI0/XI52/XI3/MM11_d
+ N_XI0/XI52/XI3/NET35_XI0/XI52/XI3/MM11_g N_VDD_XI0/XI52/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI4/MM2 N_XI0/XI52/XI4/NET34_XI0/XI52/XI4/MM2_d
+ N_XI0/XI52/XI4/NET33_XI0/XI52/XI4/MM2_g N_VSS_XI0/XI52/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM3 N_XI0/XI52/XI4/NET33_XI0/XI52/XI4/MM3_d
+ N_WL<100>_XI0/XI52/XI4/MM3_g N_BLN<11>_XI0/XI52/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM0 N_XI0/XI52/XI4/NET34_XI0/XI52/XI4/MM0_d
+ N_WL<100>_XI0/XI52/XI4/MM0_g N_BL<11>_XI0/XI52/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM1 N_XI0/XI52/XI4/NET33_XI0/XI52/XI4/MM1_d
+ N_XI0/XI52/XI4/NET34_XI0/XI52/XI4/MM1_g N_VSS_XI0/XI52/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM9 N_XI0/XI52/XI4/NET36_XI0/XI52/XI4/MM9_d
+ N_WL<101>_XI0/XI52/XI4/MM9_g N_BL<11>_XI0/XI52/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM6 N_XI0/XI52/XI4/NET35_XI0/XI52/XI4/MM6_d
+ N_XI0/XI52/XI4/NET36_XI0/XI52/XI4/MM6_g N_VSS_XI0/XI52/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM7 N_XI0/XI52/XI4/NET36_XI0/XI52/XI4/MM7_d
+ N_XI0/XI52/XI4/NET35_XI0/XI52/XI4/MM7_g N_VSS_XI0/XI52/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM8 N_XI0/XI52/XI4/NET35_XI0/XI52/XI4/MM8_d
+ N_WL<101>_XI0/XI52/XI4/MM8_g N_BLN<11>_XI0/XI52/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI4/MM5 N_XI0/XI52/XI4/NET34_XI0/XI52/XI4/MM5_d
+ N_XI0/XI52/XI4/NET33_XI0/XI52/XI4/MM5_g N_VDD_XI0/XI52/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI4/MM4 N_XI0/XI52/XI4/NET33_XI0/XI52/XI4/MM4_d
+ N_XI0/XI52/XI4/NET34_XI0/XI52/XI4/MM4_g N_VDD_XI0/XI52/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI4/MM10 N_XI0/XI52/XI4/NET35_XI0/XI52/XI4/MM10_d
+ N_XI0/XI52/XI4/NET36_XI0/XI52/XI4/MM10_g N_VDD_XI0/XI52/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI4/MM11 N_XI0/XI52/XI4/NET36_XI0/XI52/XI4/MM11_d
+ N_XI0/XI52/XI4/NET35_XI0/XI52/XI4/MM11_g N_VDD_XI0/XI52/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI5/MM2 N_XI0/XI52/XI5/NET34_XI0/XI52/XI5/MM2_d
+ N_XI0/XI52/XI5/NET33_XI0/XI52/XI5/MM2_g N_VSS_XI0/XI52/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM3 N_XI0/XI52/XI5/NET33_XI0/XI52/XI5/MM3_d
+ N_WL<100>_XI0/XI52/XI5/MM3_g N_BLN<10>_XI0/XI52/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM0 N_XI0/XI52/XI5/NET34_XI0/XI52/XI5/MM0_d
+ N_WL<100>_XI0/XI52/XI5/MM0_g N_BL<10>_XI0/XI52/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM1 N_XI0/XI52/XI5/NET33_XI0/XI52/XI5/MM1_d
+ N_XI0/XI52/XI5/NET34_XI0/XI52/XI5/MM1_g N_VSS_XI0/XI52/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM9 N_XI0/XI52/XI5/NET36_XI0/XI52/XI5/MM9_d
+ N_WL<101>_XI0/XI52/XI5/MM9_g N_BL<10>_XI0/XI52/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM6 N_XI0/XI52/XI5/NET35_XI0/XI52/XI5/MM6_d
+ N_XI0/XI52/XI5/NET36_XI0/XI52/XI5/MM6_g N_VSS_XI0/XI52/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM7 N_XI0/XI52/XI5/NET36_XI0/XI52/XI5/MM7_d
+ N_XI0/XI52/XI5/NET35_XI0/XI52/XI5/MM7_g N_VSS_XI0/XI52/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM8 N_XI0/XI52/XI5/NET35_XI0/XI52/XI5/MM8_d
+ N_WL<101>_XI0/XI52/XI5/MM8_g N_BLN<10>_XI0/XI52/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI5/MM5 N_XI0/XI52/XI5/NET34_XI0/XI52/XI5/MM5_d
+ N_XI0/XI52/XI5/NET33_XI0/XI52/XI5/MM5_g N_VDD_XI0/XI52/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI5/MM4 N_XI0/XI52/XI5/NET33_XI0/XI52/XI5/MM4_d
+ N_XI0/XI52/XI5/NET34_XI0/XI52/XI5/MM4_g N_VDD_XI0/XI52/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI5/MM10 N_XI0/XI52/XI5/NET35_XI0/XI52/XI5/MM10_d
+ N_XI0/XI52/XI5/NET36_XI0/XI52/XI5/MM10_g N_VDD_XI0/XI52/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI5/MM11 N_XI0/XI52/XI5/NET36_XI0/XI52/XI5/MM11_d
+ N_XI0/XI52/XI5/NET35_XI0/XI52/XI5/MM11_g N_VDD_XI0/XI52/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI6/MM2 N_XI0/XI52/XI6/NET34_XI0/XI52/XI6/MM2_d
+ N_XI0/XI52/XI6/NET33_XI0/XI52/XI6/MM2_g N_VSS_XI0/XI52/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM3 N_XI0/XI52/XI6/NET33_XI0/XI52/XI6/MM3_d
+ N_WL<100>_XI0/XI52/XI6/MM3_g N_BLN<9>_XI0/XI52/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM0 N_XI0/XI52/XI6/NET34_XI0/XI52/XI6/MM0_d
+ N_WL<100>_XI0/XI52/XI6/MM0_g N_BL<9>_XI0/XI52/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM1 N_XI0/XI52/XI6/NET33_XI0/XI52/XI6/MM1_d
+ N_XI0/XI52/XI6/NET34_XI0/XI52/XI6/MM1_g N_VSS_XI0/XI52/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM9 N_XI0/XI52/XI6/NET36_XI0/XI52/XI6/MM9_d
+ N_WL<101>_XI0/XI52/XI6/MM9_g N_BL<9>_XI0/XI52/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM6 N_XI0/XI52/XI6/NET35_XI0/XI52/XI6/MM6_d
+ N_XI0/XI52/XI6/NET36_XI0/XI52/XI6/MM6_g N_VSS_XI0/XI52/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM7 N_XI0/XI52/XI6/NET36_XI0/XI52/XI6/MM7_d
+ N_XI0/XI52/XI6/NET35_XI0/XI52/XI6/MM7_g N_VSS_XI0/XI52/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM8 N_XI0/XI52/XI6/NET35_XI0/XI52/XI6/MM8_d
+ N_WL<101>_XI0/XI52/XI6/MM8_g N_BLN<9>_XI0/XI52/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI6/MM5 N_XI0/XI52/XI6/NET34_XI0/XI52/XI6/MM5_d
+ N_XI0/XI52/XI6/NET33_XI0/XI52/XI6/MM5_g N_VDD_XI0/XI52/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI6/MM4 N_XI0/XI52/XI6/NET33_XI0/XI52/XI6/MM4_d
+ N_XI0/XI52/XI6/NET34_XI0/XI52/XI6/MM4_g N_VDD_XI0/XI52/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI6/MM10 N_XI0/XI52/XI6/NET35_XI0/XI52/XI6/MM10_d
+ N_XI0/XI52/XI6/NET36_XI0/XI52/XI6/MM10_g N_VDD_XI0/XI52/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI6/MM11 N_XI0/XI52/XI6/NET36_XI0/XI52/XI6/MM11_d
+ N_XI0/XI52/XI6/NET35_XI0/XI52/XI6/MM11_g N_VDD_XI0/XI52/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI7/MM2 N_XI0/XI52/XI7/NET34_XI0/XI52/XI7/MM2_d
+ N_XI0/XI52/XI7/NET33_XI0/XI52/XI7/MM2_g N_VSS_XI0/XI52/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM3 N_XI0/XI52/XI7/NET33_XI0/XI52/XI7/MM3_d
+ N_WL<100>_XI0/XI52/XI7/MM3_g N_BLN<8>_XI0/XI52/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM0 N_XI0/XI52/XI7/NET34_XI0/XI52/XI7/MM0_d
+ N_WL<100>_XI0/XI52/XI7/MM0_g N_BL<8>_XI0/XI52/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM1 N_XI0/XI52/XI7/NET33_XI0/XI52/XI7/MM1_d
+ N_XI0/XI52/XI7/NET34_XI0/XI52/XI7/MM1_g N_VSS_XI0/XI52/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM9 N_XI0/XI52/XI7/NET36_XI0/XI52/XI7/MM9_d
+ N_WL<101>_XI0/XI52/XI7/MM9_g N_BL<8>_XI0/XI52/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM6 N_XI0/XI52/XI7/NET35_XI0/XI52/XI7/MM6_d
+ N_XI0/XI52/XI7/NET36_XI0/XI52/XI7/MM6_g N_VSS_XI0/XI52/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM7 N_XI0/XI52/XI7/NET36_XI0/XI52/XI7/MM7_d
+ N_XI0/XI52/XI7/NET35_XI0/XI52/XI7/MM7_g N_VSS_XI0/XI52/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM8 N_XI0/XI52/XI7/NET35_XI0/XI52/XI7/MM8_d
+ N_WL<101>_XI0/XI52/XI7/MM8_g N_BLN<8>_XI0/XI52/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI7/MM5 N_XI0/XI52/XI7/NET34_XI0/XI52/XI7/MM5_d
+ N_XI0/XI52/XI7/NET33_XI0/XI52/XI7/MM5_g N_VDD_XI0/XI52/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI7/MM4 N_XI0/XI52/XI7/NET33_XI0/XI52/XI7/MM4_d
+ N_XI0/XI52/XI7/NET34_XI0/XI52/XI7/MM4_g N_VDD_XI0/XI52/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI7/MM10 N_XI0/XI52/XI7/NET35_XI0/XI52/XI7/MM10_d
+ N_XI0/XI52/XI7/NET36_XI0/XI52/XI7/MM10_g N_VDD_XI0/XI52/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI7/MM11 N_XI0/XI52/XI7/NET36_XI0/XI52/XI7/MM11_d
+ N_XI0/XI52/XI7/NET35_XI0/XI52/XI7/MM11_g N_VDD_XI0/XI52/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI8/MM2 N_XI0/XI52/XI8/NET34_XI0/XI52/XI8/MM2_d
+ N_XI0/XI52/XI8/NET33_XI0/XI52/XI8/MM2_g N_VSS_XI0/XI52/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM3 N_XI0/XI52/XI8/NET33_XI0/XI52/XI8/MM3_d
+ N_WL<100>_XI0/XI52/XI8/MM3_g N_BLN<7>_XI0/XI52/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM0 N_XI0/XI52/XI8/NET34_XI0/XI52/XI8/MM0_d
+ N_WL<100>_XI0/XI52/XI8/MM0_g N_BL<7>_XI0/XI52/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM1 N_XI0/XI52/XI8/NET33_XI0/XI52/XI8/MM1_d
+ N_XI0/XI52/XI8/NET34_XI0/XI52/XI8/MM1_g N_VSS_XI0/XI52/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM9 N_XI0/XI52/XI8/NET36_XI0/XI52/XI8/MM9_d
+ N_WL<101>_XI0/XI52/XI8/MM9_g N_BL<7>_XI0/XI52/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM6 N_XI0/XI52/XI8/NET35_XI0/XI52/XI8/MM6_d
+ N_XI0/XI52/XI8/NET36_XI0/XI52/XI8/MM6_g N_VSS_XI0/XI52/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM7 N_XI0/XI52/XI8/NET36_XI0/XI52/XI8/MM7_d
+ N_XI0/XI52/XI8/NET35_XI0/XI52/XI8/MM7_g N_VSS_XI0/XI52/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM8 N_XI0/XI52/XI8/NET35_XI0/XI52/XI8/MM8_d
+ N_WL<101>_XI0/XI52/XI8/MM8_g N_BLN<7>_XI0/XI52/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI8/MM5 N_XI0/XI52/XI8/NET34_XI0/XI52/XI8/MM5_d
+ N_XI0/XI52/XI8/NET33_XI0/XI52/XI8/MM5_g N_VDD_XI0/XI52/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI8/MM4 N_XI0/XI52/XI8/NET33_XI0/XI52/XI8/MM4_d
+ N_XI0/XI52/XI8/NET34_XI0/XI52/XI8/MM4_g N_VDD_XI0/XI52/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI8/MM10 N_XI0/XI52/XI8/NET35_XI0/XI52/XI8/MM10_d
+ N_XI0/XI52/XI8/NET36_XI0/XI52/XI8/MM10_g N_VDD_XI0/XI52/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI8/MM11 N_XI0/XI52/XI8/NET36_XI0/XI52/XI8/MM11_d
+ N_XI0/XI52/XI8/NET35_XI0/XI52/XI8/MM11_g N_VDD_XI0/XI52/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI9/MM2 N_XI0/XI52/XI9/NET34_XI0/XI52/XI9/MM2_d
+ N_XI0/XI52/XI9/NET33_XI0/XI52/XI9/MM2_g N_VSS_XI0/XI52/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM3 N_XI0/XI52/XI9/NET33_XI0/XI52/XI9/MM3_d
+ N_WL<100>_XI0/XI52/XI9/MM3_g N_BLN<6>_XI0/XI52/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM0 N_XI0/XI52/XI9/NET34_XI0/XI52/XI9/MM0_d
+ N_WL<100>_XI0/XI52/XI9/MM0_g N_BL<6>_XI0/XI52/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM1 N_XI0/XI52/XI9/NET33_XI0/XI52/XI9/MM1_d
+ N_XI0/XI52/XI9/NET34_XI0/XI52/XI9/MM1_g N_VSS_XI0/XI52/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM9 N_XI0/XI52/XI9/NET36_XI0/XI52/XI9/MM9_d
+ N_WL<101>_XI0/XI52/XI9/MM9_g N_BL<6>_XI0/XI52/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM6 N_XI0/XI52/XI9/NET35_XI0/XI52/XI9/MM6_d
+ N_XI0/XI52/XI9/NET36_XI0/XI52/XI9/MM6_g N_VSS_XI0/XI52/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM7 N_XI0/XI52/XI9/NET36_XI0/XI52/XI9/MM7_d
+ N_XI0/XI52/XI9/NET35_XI0/XI52/XI9/MM7_g N_VSS_XI0/XI52/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM8 N_XI0/XI52/XI9/NET35_XI0/XI52/XI9/MM8_d
+ N_WL<101>_XI0/XI52/XI9/MM8_g N_BLN<6>_XI0/XI52/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI9/MM5 N_XI0/XI52/XI9/NET34_XI0/XI52/XI9/MM5_d
+ N_XI0/XI52/XI9/NET33_XI0/XI52/XI9/MM5_g N_VDD_XI0/XI52/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI9/MM4 N_XI0/XI52/XI9/NET33_XI0/XI52/XI9/MM4_d
+ N_XI0/XI52/XI9/NET34_XI0/XI52/XI9/MM4_g N_VDD_XI0/XI52/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI9/MM10 N_XI0/XI52/XI9/NET35_XI0/XI52/XI9/MM10_d
+ N_XI0/XI52/XI9/NET36_XI0/XI52/XI9/MM10_g N_VDD_XI0/XI52/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI9/MM11 N_XI0/XI52/XI9/NET36_XI0/XI52/XI9/MM11_d
+ N_XI0/XI52/XI9/NET35_XI0/XI52/XI9/MM11_g N_VDD_XI0/XI52/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI10/MM2 N_XI0/XI52/XI10/NET34_XI0/XI52/XI10/MM2_d
+ N_XI0/XI52/XI10/NET33_XI0/XI52/XI10/MM2_g N_VSS_XI0/XI52/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM3 N_XI0/XI52/XI10/NET33_XI0/XI52/XI10/MM3_d
+ N_WL<100>_XI0/XI52/XI10/MM3_g N_BLN<5>_XI0/XI52/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM0 N_XI0/XI52/XI10/NET34_XI0/XI52/XI10/MM0_d
+ N_WL<100>_XI0/XI52/XI10/MM0_g N_BL<5>_XI0/XI52/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM1 N_XI0/XI52/XI10/NET33_XI0/XI52/XI10/MM1_d
+ N_XI0/XI52/XI10/NET34_XI0/XI52/XI10/MM1_g N_VSS_XI0/XI52/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM9 N_XI0/XI52/XI10/NET36_XI0/XI52/XI10/MM9_d
+ N_WL<101>_XI0/XI52/XI10/MM9_g N_BL<5>_XI0/XI52/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM6 N_XI0/XI52/XI10/NET35_XI0/XI52/XI10/MM6_d
+ N_XI0/XI52/XI10/NET36_XI0/XI52/XI10/MM6_g N_VSS_XI0/XI52/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM7 N_XI0/XI52/XI10/NET36_XI0/XI52/XI10/MM7_d
+ N_XI0/XI52/XI10/NET35_XI0/XI52/XI10/MM7_g N_VSS_XI0/XI52/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM8 N_XI0/XI52/XI10/NET35_XI0/XI52/XI10/MM8_d
+ N_WL<101>_XI0/XI52/XI10/MM8_g N_BLN<5>_XI0/XI52/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI10/MM5 N_XI0/XI52/XI10/NET34_XI0/XI52/XI10/MM5_d
+ N_XI0/XI52/XI10/NET33_XI0/XI52/XI10/MM5_g N_VDD_XI0/XI52/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI10/MM4 N_XI0/XI52/XI10/NET33_XI0/XI52/XI10/MM4_d
+ N_XI0/XI52/XI10/NET34_XI0/XI52/XI10/MM4_g N_VDD_XI0/XI52/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI10/MM10 N_XI0/XI52/XI10/NET35_XI0/XI52/XI10/MM10_d
+ N_XI0/XI52/XI10/NET36_XI0/XI52/XI10/MM10_g N_VDD_XI0/XI52/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI10/MM11 N_XI0/XI52/XI10/NET36_XI0/XI52/XI10/MM11_d
+ N_XI0/XI52/XI10/NET35_XI0/XI52/XI10/MM11_g N_VDD_XI0/XI52/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI11/MM2 N_XI0/XI52/XI11/NET34_XI0/XI52/XI11/MM2_d
+ N_XI0/XI52/XI11/NET33_XI0/XI52/XI11/MM2_g N_VSS_XI0/XI52/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM3 N_XI0/XI52/XI11/NET33_XI0/XI52/XI11/MM3_d
+ N_WL<100>_XI0/XI52/XI11/MM3_g N_BLN<4>_XI0/XI52/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM0 N_XI0/XI52/XI11/NET34_XI0/XI52/XI11/MM0_d
+ N_WL<100>_XI0/XI52/XI11/MM0_g N_BL<4>_XI0/XI52/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM1 N_XI0/XI52/XI11/NET33_XI0/XI52/XI11/MM1_d
+ N_XI0/XI52/XI11/NET34_XI0/XI52/XI11/MM1_g N_VSS_XI0/XI52/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM9 N_XI0/XI52/XI11/NET36_XI0/XI52/XI11/MM9_d
+ N_WL<101>_XI0/XI52/XI11/MM9_g N_BL<4>_XI0/XI52/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM6 N_XI0/XI52/XI11/NET35_XI0/XI52/XI11/MM6_d
+ N_XI0/XI52/XI11/NET36_XI0/XI52/XI11/MM6_g N_VSS_XI0/XI52/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM7 N_XI0/XI52/XI11/NET36_XI0/XI52/XI11/MM7_d
+ N_XI0/XI52/XI11/NET35_XI0/XI52/XI11/MM7_g N_VSS_XI0/XI52/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM8 N_XI0/XI52/XI11/NET35_XI0/XI52/XI11/MM8_d
+ N_WL<101>_XI0/XI52/XI11/MM8_g N_BLN<4>_XI0/XI52/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI11/MM5 N_XI0/XI52/XI11/NET34_XI0/XI52/XI11/MM5_d
+ N_XI0/XI52/XI11/NET33_XI0/XI52/XI11/MM5_g N_VDD_XI0/XI52/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI11/MM4 N_XI0/XI52/XI11/NET33_XI0/XI52/XI11/MM4_d
+ N_XI0/XI52/XI11/NET34_XI0/XI52/XI11/MM4_g N_VDD_XI0/XI52/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI11/MM10 N_XI0/XI52/XI11/NET35_XI0/XI52/XI11/MM10_d
+ N_XI0/XI52/XI11/NET36_XI0/XI52/XI11/MM10_g N_VDD_XI0/XI52/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI11/MM11 N_XI0/XI52/XI11/NET36_XI0/XI52/XI11/MM11_d
+ N_XI0/XI52/XI11/NET35_XI0/XI52/XI11/MM11_g N_VDD_XI0/XI52/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI12/MM2 N_XI0/XI52/XI12/NET34_XI0/XI52/XI12/MM2_d
+ N_XI0/XI52/XI12/NET33_XI0/XI52/XI12/MM2_g N_VSS_XI0/XI52/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM3 N_XI0/XI52/XI12/NET33_XI0/XI52/XI12/MM3_d
+ N_WL<100>_XI0/XI52/XI12/MM3_g N_BLN<3>_XI0/XI52/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM0 N_XI0/XI52/XI12/NET34_XI0/XI52/XI12/MM0_d
+ N_WL<100>_XI0/XI52/XI12/MM0_g N_BL<3>_XI0/XI52/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM1 N_XI0/XI52/XI12/NET33_XI0/XI52/XI12/MM1_d
+ N_XI0/XI52/XI12/NET34_XI0/XI52/XI12/MM1_g N_VSS_XI0/XI52/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM9 N_XI0/XI52/XI12/NET36_XI0/XI52/XI12/MM9_d
+ N_WL<101>_XI0/XI52/XI12/MM9_g N_BL<3>_XI0/XI52/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM6 N_XI0/XI52/XI12/NET35_XI0/XI52/XI12/MM6_d
+ N_XI0/XI52/XI12/NET36_XI0/XI52/XI12/MM6_g N_VSS_XI0/XI52/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM7 N_XI0/XI52/XI12/NET36_XI0/XI52/XI12/MM7_d
+ N_XI0/XI52/XI12/NET35_XI0/XI52/XI12/MM7_g N_VSS_XI0/XI52/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM8 N_XI0/XI52/XI12/NET35_XI0/XI52/XI12/MM8_d
+ N_WL<101>_XI0/XI52/XI12/MM8_g N_BLN<3>_XI0/XI52/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI12/MM5 N_XI0/XI52/XI12/NET34_XI0/XI52/XI12/MM5_d
+ N_XI0/XI52/XI12/NET33_XI0/XI52/XI12/MM5_g N_VDD_XI0/XI52/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI12/MM4 N_XI0/XI52/XI12/NET33_XI0/XI52/XI12/MM4_d
+ N_XI0/XI52/XI12/NET34_XI0/XI52/XI12/MM4_g N_VDD_XI0/XI52/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI12/MM10 N_XI0/XI52/XI12/NET35_XI0/XI52/XI12/MM10_d
+ N_XI0/XI52/XI12/NET36_XI0/XI52/XI12/MM10_g N_VDD_XI0/XI52/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI12/MM11 N_XI0/XI52/XI12/NET36_XI0/XI52/XI12/MM11_d
+ N_XI0/XI52/XI12/NET35_XI0/XI52/XI12/MM11_g N_VDD_XI0/XI52/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI13/MM2 N_XI0/XI52/XI13/NET34_XI0/XI52/XI13/MM2_d
+ N_XI0/XI52/XI13/NET33_XI0/XI52/XI13/MM2_g N_VSS_XI0/XI52/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM3 N_XI0/XI52/XI13/NET33_XI0/XI52/XI13/MM3_d
+ N_WL<100>_XI0/XI52/XI13/MM3_g N_BLN<2>_XI0/XI52/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM0 N_XI0/XI52/XI13/NET34_XI0/XI52/XI13/MM0_d
+ N_WL<100>_XI0/XI52/XI13/MM0_g N_BL<2>_XI0/XI52/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM1 N_XI0/XI52/XI13/NET33_XI0/XI52/XI13/MM1_d
+ N_XI0/XI52/XI13/NET34_XI0/XI52/XI13/MM1_g N_VSS_XI0/XI52/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM9 N_XI0/XI52/XI13/NET36_XI0/XI52/XI13/MM9_d
+ N_WL<101>_XI0/XI52/XI13/MM9_g N_BL<2>_XI0/XI52/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM6 N_XI0/XI52/XI13/NET35_XI0/XI52/XI13/MM6_d
+ N_XI0/XI52/XI13/NET36_XI0/XI52/XI13/MM6_g N_VSS_XI0/XI52/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM7 N_XI0/XI52/XI13/NET36_XI0/XI52/XI13/MM7_d
+ N_XI0/XI52/XI13/NET35_XI0/XI52/XI13/MM7_g N_VSS_XI0/XI52/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM8 N_XI0/XI52/XI13/NET35_XI0/XI52/XI13/MM8_d
+ N_WL<101>_XI0/XI52/XI13/MM8_g N_BLN<2>_XI0/XI52/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI13/MM5 N_XI0/XI52/XI13/NET34_XI0/XI52/XI13/MM5_d
+ N_XI0/XI52/XI13/NET33_XI0/XI52/XI13/MM5_g N_VDD_XI0/XI52/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI13/MM4 N_XI0/XI52/XI13/NET33_XI0/XI52/XI13/MM4_d
+ N_XI0/XI52/XI13/NET34_XI0/XI52/XI13/MM4_g N_VDD_XI0/XI52/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI13/MM10 N_XI0/XI52/XI13/NET35_XI0/XI52/XI13/MM10_d
+ N_XI0/XI52/XI13/NET36_XI0/XI52/XI13/MM10_g N_VDD_XI0/XI52/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI13/MM11 N_XI0/XI52/XI13/NET36_XI0/XI52/XI13/MM11_d
+ N_XI0/XI52/XI13/NET35_XI0/XI52/XI13/MM11_g N_VDD_XI0/XI52/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI14/MM2 N_XI0/XI52/XI14/NET34_XI0/XI52/XI14/MM2_d
+ N_XI0/XI52/XI14/NET33_XI0/XI52/XI14/MM2_g N_VSS_XI0/XI52/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM3 N_XI0/XI52/XI14/NET33_XI0/XI52/XI14/MM3_d
+ N_WL<100>_XI0/XI52/XI14/MM3_g N_BLN<1>_XI0/XI52/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM0 N_XI0/XI52/XI14/NET34_XI0/XI52/XI14/MM0_d
+ N_WL<100>_XI0/XI52/XI14/MM0_g N_BL<1>_XI0/XI52/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM1 N_XI0/XI52/XI14/NET33_XI0/XI52/XI14/MM1_d
+ N_XI0/XI52/XI14/NET34_XI0/XI52/XI14/MM1_g N_VSS_XI0/XI52/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM9 N_XI0/XI52/XI14/NET36_XI0/XI52/XI14/MM9_d
+ N_WL<101>_XI0/XI52/XI14/MM9_g N_BL<1>_XI0/XI52/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM6 N_XI0/XI52/XI14/NET35_XI0/XI52/XI14/MM6_d
+ N_XI0/XI52/XI14/NET36_XI0/XI52/XI14/MM6_g N_VSS_XI0/XI52/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM7 N_XI0/XI52/XI14/NET36_XI0/XI52/XI14/MM7_d
+ N_XI0/XI52/XI14/NET35_XI0/XI52/XI14/MM7_g N_VSS_XI0/XI52/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM8 N_XI0/XI52/XI14/NET35_XI0/XI52/XI14/MM8_d
+ N_WL<101>_XI0/XI52/XI14/MM8_g N_BLN<1>_XI0/XI52/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI14/MM5 N_XI0/XI52/XI14/NET34_XI0/XI52/XI14/MM5_d
+ N_XI0/XI52/XI14/NET33_XI0/XI52/XI14/MM5_g N_VDD_XI0/XI52/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI14/MM4 N_XI0/XI52/XI14/NET33_XI0/XI52/XI14/MM4_d
+ N_XI0/XI52/XI14/NET34_XI0/XI52/XI14/MM4_g N_VDD_XI0/XI52/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI14/MM10 N_XI0/XI52/XI14/NET35_XI0/XI52/XI14/MM10_d
+ N_XI0/XI52/XI14/NET36_XI0/XI52/XI14/MM10_g N_VDD_XI0/XI52/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI14/MM11 N_XI0/XI52/XI14/NET36_XI0/XI52/XI14/MM11_d
+ N_XI0/XI52/XI14/NET35_XI0/XI52/XI14/MM11_g N_VDD_XI0/XI52/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI15/MM2 N_XI0/XI52/XI15/NET34_XI0/XI52/XI15/MM2_d
+ N_XI0/XI52/XI15/NET33_XI0/XI52/XI15/MM2_g N_VSS_XI0/XI52/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM3 N_XI0/XI52/XI15/NET33_XI0/XI52/XI15/MM3_d
+ N_WL<100>_XI0/XI52/XI15/MM3_g N_BLN<0>_XI0/XI52/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM0 N_XI0/XI52/XI15/NET34_XI0/XI52/XI15/MM0_d
+ N_WL<100>_XI0/XI52/XI15/MM0_g N_BL<0>_XI0/XI52/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM1 N_XI0/XI52/XI15/NET33_XI0/XI52/XI15/MM1_d
+ N_XI0/XI52/XI15/NET34_XI0/XI52/XI15/MM1_g N_VSS_XI0/XI52/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM9 N_XI0/XI52/XI15/NET36_XI0/XI52/XI15/MM9_d
+ N_WL<101>_XI0/XI52/XI15/MM9_g N_BL<0>_XI0/XI52/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM6 N_XI0/XI52/XI15/NET35_XI0/XI52/XI15/MM6_d
+ N_XI0/XI52/XI15/NET36_XI0/XI52/XI15/MM6_g N_VSS_XI0/XI52/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM7 N_XI0/XI52/XI15/NET36_XI0/XI52/XI15/MM7_d
+ N_XI0/XI52/XI15/NET35_XI0/XI52/XI15/MM7_g N_VSS_XI0/XI52/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM8 N_XI0/XI52/XI15/NET35_XI0/XI52/XI15/MM8_d
+ N_WL<101>_XI0/XI52/XI15/MM8_g N_BLN<0>_XI0/XI52/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI52/XI15/MM5 N_XI0/XI52/XI15/NET34_XI0/XI52/XI15/MM5_d
+ N_XI0/XI52/XI15/NET33_XI0/XI52/XI15/MM5_g N_VDD_XI0/XI52/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI15/MM4 N_XI0/XI52/XI15/NET33_XI0/XI52/XI15/MM4_d
+ N_XI0/XI52/XI15/NET34_XI0/XI52/XI15/MM4_g N_VDD_XI0/XI52/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI15/MM10 N_XI0/XI52/XI15/NET35_XI0/XI52/XI15/MM10_d
+ N_XI0/XI52/XI15/NET36_XI0/XI52/XI15/MM10_g N_VDD_XI0/XI52/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI52/XI15/MM11 N_XI0/XI52/XI15/NET36_XI0/XI52/XI15/MM11_d
+ N_XI0/XI52/XI15/NET35_XI0/XI52/XI15/MM11_g N_VDD_XI0/XI52/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI0/MM2 N_XI0/XI53/XI0/NET34_XI0/XI53/XI0/MM2_d
+ N_XI0/XI53/XI0/NET33_XI0/XI53/XI0/MM2_g N_VSS_XI0/XI53/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM3 N_XI0/XI53/XI0/NET33_XI0/XI53/XI0/MM3_d
+ N_WL<102>_XI0/XI53/XI0/MM3_g N_BLN<15>_XI0/XI53/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM0 N_XI0/XI53/XI0/NET34_XI0/XI53/XI0/MM0_d
+ N_WL<102>_XI0/XI53/XI0/MM0_g N_BL<15>_XI0/XI53/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM1 N_XI0/XI53/XI0/NET33_XI0/XI53/XI0/MM1_d
+ N_XI0/XI53/XI0/NET34_XI0/XI53/XI0/MM1_g N_VSS_XI0/XI53/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM9 N_XI0/XI53/XI0/NET36_XI0/XI53/XI0/MM9_d
+ N_WL<103>_XI0/XI53/XI0/MM9_g N_BL<15>_XI0/XI53/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM6 N_XI0/XI53/XI0/NET35_XI0/XI53/XI0/MM6_d
+ N_XI0/XI53/XI0/NET36_XI0/XI53/XI0/MM6_g N_VSS_XI0/XI53/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM7 N_XI0/XI53/XI0/NET36_XI0/XI53/XI0/MM7_d
+ N_XI0/XI53/XI0/NET35_XI0/XI53/XI0/MM7_g N_VSS_XI0/XI53/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM8 N_XI0/XI53/XI0/NET35_XI0/XI53/XI0/MM8_d
+ N_WL<103>_XI0/XI53/XI0/MM8_g N_BLN<15>_XI0/XI53/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI0/MM5 N_XI0/XI53/XI0/NET34_XI0/XI53/XI0/MM5_d
+ N_XI0/XI53/XI0/NET33_XI0/XI53/XI0/MM5_g N_VDD_XI0/XI53/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI0/MM4 N_XI0/XI53/XI0/NET33_XI0/XI53/XI0/MM4_d
+ N_XI0/XI53/XI0/NET34_XI0/XI53/XI0/MM4_g N_VDD_XI0/XI53/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI0/MM10 N_XI0/XI53/XI0/NET35_XI0/XI53/XI0/MM10_d
+ N_XI0/XI53/XI0/NET36_XI0/XI53/XI0/MM10_g N_VDD_XI0/XI53/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI0/MM11 N_XI0/XI53/XI0/NET36_XI0/XI53/XI0/MM11_d
+ N_XI0/XI53/XI0/NET35_XI0/XI53/XI0/MM11_g N_VDD_XI0/XI53/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI1/MM2 N_XI0/XI53/XI1/NET34_XI0/XI53/XI1/MM2_d
+ N_XI0/XI53/XI1/NET33_XI0/XI53/XI1/MM2_g N_VSS_XI0/XI53/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM3 N_XI0/XI53/XI1/NET33_XI0/XI53/XI1/MM3_d
+ N_WL<102>_XI0/XI53/XI1/MM3_g N_BLN<14>_XI0/XI53/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM0 N_XI0/XI53/XI1/NET34_XI0/XI53/XI1/MM0_d
+ N_WL<102>_XI0/XI53/XI1/MM0_g N_BL<14>_XI0/XI53/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM1 N_XI0/XI53/XI1/NET33_XI0/XI53/XI1/MM1_d
+ N_XI0/XI53/XI1/NET34_XI0/XI53/XI1/MM1_g N_VSS_XI0/XI53/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM9 N_XI0/XI53/XI1/NET36_XI0/XI53/XI1/MM9_d
+ N_WL<103>_XI0/XI53/XI1/MM9_g N_BL<14>_XI0/XI53/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM6 N_XI0/XI53/XI1/NET35_XI0/XI53/XI1/MM6_d
+ N_XI0/XI53/XI1/NET36_XI0/XI53/XI1/MM6_g N_VSS_XI0/XI53/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM7 N_XI0/XI53/XI1/NET36_XI0/XI53/XI1/MM7_d
+ N_XI0/XI53/XI1/NET35_XI0/XI53/XI1/MM7_g N_VSS_XI0/XI53/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM8 N_XI0/XI53/XI1/NET35_XI0/XI53/XI1/MM8_d
+ N_WL<103>_XI0/XI53/XI1/MM8_g N_BLN<14>_XI0/XI53/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI1/MM5 N_XI0/XI53/XI1/NET34_XI0/XI53/XI1/MM5_d
+ N_XI0/XI53/XI1/NET33_XI0/XI53/XI1/MM5_g N_VDD_XI0/XI53/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI1/MM4 N_XI0/XI53/XI1/NET33_XI0/XI53/XI1/MM4_d
+ N_XI0/XI53/XI1/NET34_XI0/XI53/XI1/MM4_g N_VDD_XI0/XI53/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI1/MM10 N_XI0/XI53/XI1/NET35_XI0/XI53/XI1/MM10_d
+ N_XI0/XI53/XI1/NET36_XI0/XI53/XI1/MM10_g N_VDD_XI0/XI53/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI1/MM11 N_XI0/XI53/XI1/NET36_XI0/XI53/XI1/MM11_d
+ N_XI0/XI53/XI1/NET35_XI0/XI53/XI1/MM11_g N_VDD_XI0/XI53/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI2/MM2 N_XI0/XI53/XI2/NET34_XI0/XI53/XI2/MM2_d
+ N_XI0/XI53/XI2/NET33_XI0/XI53/XI2/MM2_g N_VSS_XI0/XI53/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM3 N_XI0/XI53/XI2/NET33_XI0/XI53/XI2/MM3_d
+ N_WL<102>_XI0/XI53/XI2/MM3_g N_BLN<13>_XI0/XI53/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM0 N_XI0/XI53/XI2/NET34_XI0/XI53/XI2/MM0_d
+ N_WL<102>_XI0/XI53/XI2/MM0_g N_BL<13>_XI0/XI53/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM1 N_XI0/XI53/XI2/NET33_XI0/XI53/XI2/MM1_d
+ N_XI0/XI53/XI2/NET34_XI0/XI53/XI2/MM1_g N_VSS_XI0/XI53/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM9 N_XI0/XI53/XI2/NET36_XI0/XI53/XI2/MM9_d
+ N_WL<103>_XI0/XI53/XI2/MM9_g N_BL<13>_XI0/XI53/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM6 N_XI0/XI53/XI2/NET35_XI0/XI53/XI2/MM6_d
+ N_XI0/XI53/XI2/NET36_XI0/XI53/XI2/MM6_g N_VSS_XI0/XI53/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM7 N_XI0/XI53/XI2/NET36_XI0/XI53/XI2/MM7_d
+ N_XI0/XI53/XI2/NET35_XI0/XI53/XI2/MM7_g N_VSS_XI0/XI53/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM8 N_XI0/XI53/XI2/NET35_XI0/XI53/XI2/MM8_d
+ N_WL<103>_XI0/XI53/XI2/MM8_g N_BLN<13>_XI0/XI53/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI2/MM5 N_XI0/XI53/XI2/NET34_XI0/XI53/XI2/MM5_d
+ N_XI0/XI53/XI2/NET33_XI0/XI53/XI2/MM5_g N_VDD_XI0/XI53/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI2/MM4 N_XI0/XI53/XI2/NET33_XI0/XI53/XI2/MM4_d
+ N_XI0/XI53/XI2/NET34_XI0/XI53/XI2/MM4_g N_VDD_XI0/XI53/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI2/MM10 N_XI0/XI53/XI2/NET35_XI0/XI53/XI2/MM10_d
+ N_XI0/XI53/XI2/NET36_XI0/XI53/XI2/MM10_g N_VDD_XI0/XI53/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI2/MM11 N_XI0/XI53/XI2/NET36_XI0/XI53/XI2/MM11_d
+ N_XI0/XI53/XI2/NET35_XI0/XI53/XI2/MM11_g N_VDD_XI0/XI53/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI3/MM2 N_XI0/XI53/XI3/NET34_XI0/XI53/XI3/MM2_d
+ N_XI0/XI53/XI3/NET33_XI0/XI53/XI3/MM2_g N_VSS_XI0/XI53/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM3 N_XI0/XI53/XI3/NET33_XI0/XI53/XI3/MM3_d
+ N_WL<102>_XI0/XI53/XI3/MM3_g N_BLN<12>_XI0/XI53/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM0 N_XI0/XI53/XI3/NET34_XI0/XI53/XI3/MM0_d
+ N_WL<102>_XI0/XI53/XI3/MM0_g N_BL<12>_XI0/XI53/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM1 N_XI0/XI53/XI3/NET33_XI0/XI53/XI3/MM1_d
+ N_XI0/XI53/XI3/NET34_XI0/XI53/XI3/MM1_g N_VSS_XI0/XI53/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM9 N_XI0/XI53/XI3/NET36_XI0/XI53/XI3/MM9_d
+ N_WL<103>_XI0/XI53/XI3/MM9_g N_BL<12>_XI0/XI53/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM6 N_XI0/XI53/XI3/NET35_XI0/XI53/XI3/MM6_d
+ N_XI0/XI53/XI3/NET36_XI0/XI53/XI3/MM6_g N_VSS_XI0/XI53/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM7 N_XI0/XI53/XI3/NET36_XI0/XI53/XI3/MM7_d
+ N_XI0/XI53/XI3/NET35_XI0/XI53/XI3/MM7_g N_VSS_XI0/XI53/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM8 N_XI0/XI53/XI3/NET35_XI0/XI53/XI3/MM8_d
+ N_WL<103>_XI0/XI53/XI3/MM8_g N_BLN<12>_XI0/XI53/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI3/MM5 N_XI0/XI53/XI3/NET34_XI0/XI53/XI3/MM5_d
+ N_XI0/XI53/XI3/NET33_XI0/XI53/XI3/MM5_g N_VDD_XI0/XI53/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI3/MM4 N_XI0/XI53/XI3/NET33_XI0/XI53/XI3/MM4_d
+ N_XI0/XI53/XI3/NET34_XI0/XI53/XI3/MM4_g N_VDD_XI0/XI53/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI3/MM10 N_XI0/XI53/XI3/NET35_XI0/XI53/XI3/MM10_d
+ N_XI0/XI53/XI3/NET36_XI0/XI53/XI3/MM10_g N_VDD_XI0/XI53/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI3/MM11 N_XI0/XI53/XI3/NET36_XI0/XI53/XI3/MM11_d
+ N_XI0/XI53/XI3/NET35_XI0/XI53/XI3/MM11_g N_VDD_XI0/XI53/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI4/MM2 N_XI0/XI53/XI4/NET34_XI0/XI53/XI4/MM2_d
+ N_XI0/XI53/XI4/NET33_XI0/XI53/XI4/MM2_g N_VSS_XI0/XI53/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM3 N_XI0/XI53/XI4/NET33_XI0/XI53/XI4/MM3_d
+ N_WL<102>_XI0/XI53/XI4/MM3_g N_BLN<11>_XI0/XI53/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM0 N_XI0/XI53/XI4/NET34_XI0/XI53/XI4/MM0_d
+ N_WL<102>_XI0/XI53/XI4/MM0_g N_BL<11>_XI0/XI53/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM1 N_XI0/XI53/XI4/NET33_XI0/XI53/XI4/MM1_d
+ N_XI0/XI53/XI4/NET34_XI0/XI53/XI4/MM1_g N_VSS_XI0/XI53/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM9 N_XI0/XI53/XI4/NET36_XI0/XI53/XI4/MM9_d
+ N_WL<103>_XI0/XI53/XI4/MM9_g N_BL<11>_XI0/XI53/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM6 N_XI0/XI53/XI4/NET35_XI0/XI53/XI4/MM6_d
+ N_XI0/XI53/XI4/NET36_XI0/XI53/XI4/MM6_g N_VSS_XI0/XI53/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM7 N_XI0/XI53/XI4/NET36_XI0/XI53/XI4/MM7_d
+ N_XI0/XI53/XI4/NET35_XI0/XI53/XI4/MM7_g N_VSS_XI0/XI53/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM8 N_XI0/XI53/XI4/NET35_XI0/XI53/XI4/MM8_d
+ N_WL<103>_XI0/XI53/XI4/MM8_g N_BLN<11>_XI0/XI53/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI4/MM5 N_XI0/XI53/XI4/NET34_XI0/XI53/XI4/MM5_d
+ N_XI0/XI53/XI4/NET33_XI0/XI53/XI4/MM5_g N_VDD_XI0/XI53/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI4/MM4 N_XI0/XI53/XI4/NET33_XI0/XI53/XI4/MM4_d
+ N_XI0/XI53/XI4/NET34_XI0/XI53/XI4/MM4_g N_VDD_XI0/XI53/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI4/MM10 N_XI0/XI53/XI4/NET35_XI0/XI53/XI4/MM10_d
+ N_XI0/XI53/XI4/NET36_XI0/XI53/XI4/MM10_g N_VDD_XI0/XI53/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI4/MM11 N_XI0/XI53/XI4/NET36_XI0/XI53/XI4/MM11_d
+ N_XI0/XI53/XI4/NET35_XI0/XI53/XI4/MM11_g N_VDD_XI0/XI53/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI5/MM2 N_XI0/XI53/XI5/NET34_XI0/XI53/XI5/MM2_d
+ N_XI0/XI53/XI5/NET33_XI0/XI53/XI5/MM2_g N_VSS_XI0/XI53/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM3 N_XI0/XI53/XI5/NET33_XI0/XI53/XI5/MM3_d
+ N_WL<102>_XI0/XI53/XI5/MM3_g N_BLN<10>_XI0/XI53/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM0 N_XI0/XI53/XI5/NET34_XI0/XI53/XI5/MM0_d
+ N_WL<102>_XI0/XI53/XI5/MM0_g N_BL<10>_XI0/XI53/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM1 N_XI0/XI53/XI5/NET33_XI0/XI53/XI5/MM1_d
+ N_XI0/XI53/XI5/NET34_XI0/XI53/XI5/MM1_g N_VSS_XI0/XI53/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM9 N_XI0/XI53/XI5/NET36_XI0/XI53/XI5/MM9_d
+ N_WL<103>_XI0/XI53/XI5/MM9_g N_BL<10>_XI0/XI53/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM6 N_XI0/XI53/XI5/NET35_XI0/XI53/XI5/MM6_d
+ N_XI0/XI53/XI5/NET36_XI0/XI53/XI5/MM6_g N_VSS_XI0/XI53/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM7 N_XI0/XI53/XI5/NET36_XI0/XI53/XI5/MM7_d
+ N_XI0/XI53/XI5/NET35_XI0/XI53/XI5/MM7_g N_VSS_XI0/XI53/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM8 N_XI0/XI53/XI5/NET35_XI0/XI53/XI5/MM8_d
+ N_WL<103>_XI0/XI53/XI5/MM8_g N_BLN<10>_XI0/XI53/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI5/MM5 N_XI0/XI53/XI5/NET34_XI0/XI53/XI5/MM5_d
+ N_XI0/XI53/XI5/NET33_XI0/XI53/XI5/MM5_g N_VDD_XI0/XI53/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI5/MM4 N_XI0/XI53/XI5/NET33_XI0/XI53/XI5/MM4_d
+ N_XI0/XI53/XI5/NET34_XI0/XI53/XI5/MM4_g N_VDD_XI0/XI53/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI5/MM10 N_XI0/XI53/XI5/NET35_XI0/XI53/XI5/MM10_d
+ N_XI0/XI53/XI5/NET36_XI0/XI53/XI5/MM10_g N_VDD_XI0/XI53/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI5/MM11 N_XI0/XI53/XI5/NET36_XI0/XI53/XI5/MM11_d
+ N_XI0/XI53/XI5/NET35_XI0/XI53/XI5/MM11_g N_VDD_XI0/XI53/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI6/MM2 N_XI0/XI53/XI6/NET34_XI0/XI53/XI6/MM2_d
+ N_XI0/XI53/XI6/NET33_XI0/XI53/XI6/MM2_g N_VSS_XI0/XI53/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM3 N_XI0/XI53/XI6/NET33_XI0/XI53/XI6/MM3_d
+ N_WL<102>_XI0/XI53/XI6/MM3_g N_BLN<9>_XI0/XI53/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM0 N_XI0/XI53/XI6/NET34_XI0/XI53/XI6/MM0_d
+ N_WL<102>_XI0/XI53/XI6/MM0_g N_BL<9>_XI0/XI53/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM1 N_XI0/XI53/XI6/NET33_XI0/XI53/XI6/MM1_d
+ N_XI0/XI53/XI6/NET34_XI0/XI53/XI6/MM1_g N_VSS_XI0/XI53/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM9 N_XI0/XI53/XI6/NET36_XI0/XI53/XI6/MM9_d
+ N_WL<103>_XI0/XI53/XI6/MM9_g N_BL<9>_XI0/XI53/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM6 N_XI0/XI53/XI6/NET35_XI0/XI53/XI6/MM6_d
+ N_XI0/XI53/XI6/NET36_XI0/XI53/XI6/MM6_g N_VSS_XI0/XI53/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM7 N_XI0/XI53/XI6/NET36_XI0/XI53/XI6/MM7_d
+ N_XI0/XI53/XI6/NET35_XI0/XI53/XI6/MM7_g N_VSS_XI0/XI53/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM8 N_XI0/XI53/XI6/NET35_XI0/XI53/XI6/MM8_d
+ N_WL<103>_XI0/XI53/XI6/MM8_g N_BLN<9>_XI0/XI53/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI6/MM5 N_XI0/XI53/XI6/NET34_XI0/XI53/XI6/MM5_d
+ N_XI0/XI53/XI6/NET33_XI0/XI53/XI6/MM5_g N_VDD_XI0/XI53/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI6/MM4 N_XI0/XI53/XI6/NET33_XI0/XI53/XI6/MM4_d
+ N_XI0/XI53/XI6/NET34_XI0/XI53/XI6/MM4_g N_VDD_XI0/XI53/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI6/MM10 N_XI0/XI53/XI6/NET35_XI0/XI53/XI6/MM10_d
+ N_XI0/XI53/XI6/NET36_XI0/XI53/XI6/MM10_g N_VDD_XI0/XI53/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI6/MM11 N_XI0/XI53/XI6/NET36_XI0/XI53/XI6/MM11_d
+ N_XI0/XI53/XI6/NET35_XI0/XI53/XI6/MM11_g N_VDD_XI0/XI53/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI7/MM2 N_XI0/XI53/XI7/NET34_XI0/XI53/XI7/MM2_d
+ N_XI0/XI53/XI7/NET33_XI0/XI53/XI7/MM2_g N_VSS_XI0/XI53/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM3 N_XI0/XI53/XI7/NET33_XI0/XI53/XI7/MM3_d
+ N_WL<102>_XI0/XI53/XI7/MM3_g N_BLN<8>_XI0/XI53/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM0 N_XI0/XI53/XI7/NET34_XI0/XI53/XI7/MM0_d
+ N_WL<102>_XI0/XI53/XI7/MM0_g N_BL<8>_XI0/XI53/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM1 N_XI0/XI53/XI7/NET33_XI0/XI53/XI7/MM1_d
+ N_XI0/XI53/XI7/NET34_XI0/XI53/XI7/MM1_g N_VSS_XI0/XI53/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM9 N_XI0/XI53/XI7/NET36_XI0/XI53/XI7/MM9_d
+ N_WL<103>_XI0/XI53/XI7/MM9_g N_BL<8>_XI0/XI53/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM6 N_XI0/XI53/XI7/NET35_XI0/XI53/XI7/MM6_d
+ N_XI0/XI53/XI7/NET36_XI0/XI53/XI7/MM6_g N_VSS_XI0/XI53/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM7 N_XI0/XI53/XI7/NET36_XI0/XI53/XI7/MM7_d
+ N_XI0/XI53/XI7/NET35_XI0/XI53/XI7/MM7_g N_VSS_XI0/XI53/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM8 N_XI0/XI53/XI7/NET35_XI0/XI53/XI7/MM8_d
+ N_WL<103>_XI0/XI53/XI7/MM8_g N_BLN<8>_XI0/XI53/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI7/MM5 N_XI0/XI53/XI7/NET34_XI0/XI53/XI7/MM5_d
+ N_XI0/XI53/XI7/NET33_XI0/XI53/XI7/MM5_g N_VDD_XI0/XI53/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI7/MM4 N_XI0/XI53/XI7/NET33_XI0/XI53/XI7/MM4_d
+ N_XI0/XI53/XI7/NET34_XI0/XI53/XI7/MM4_g N_VDD_XI0/XI53/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI7/MM10 N_XI0/XI53/XI7/NET35_XI0/XI53/XI7/MM10_d
+ N_XI0/XI53/XI7/NET36_XI0/XI53/XI7/MM10_g N_VDD_XI0/XI53/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI7/MM11 N_XI0/XI53/XI7/NET36_XI0/XI53/XI7/MM11_d
+ N_XI0/XI53/XI7/NET35_XI0/XI53/XI7/MM11_g N_VDD_XI0/XI53/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI8/MM2 N_XI0/XI53/XI8/NET34_XI0/XI53/XI8/MM2_d
+ N_XI0/XI53/XI8/NET33_XI0/XI53/XI8/MM2_g N_VSS_XI0/XI53/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM3 N_XI0/XI53/XI8/NET33_XI0/XI53/XI8/MM3_d
+ N_WL<102>_XI0/XI53/XI8/MM3_g N_BLN<7>_XI0/XI53/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM0 N_XI0/XI53/XI8/NET34_XI0/XI53/XI8/MM0_d
+ N_WL<102>_XI0/XI53/XI8/MM0_g N_BL<7>_XI0/XI53/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM1 N_XI0/XI53/XI8/NET33_XI0/XI53/XI8/MM1_d
+ N_XI0/XI53/XI8/NET34_XI0/XI53/XI8/MM1_g N_VSS_XI0/XI53/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM9 N_XI0/XI53/XI8/NET36_XI0/XI53/XI8/MM9_d
+ N_WL<103>_XI0/XI53/XI8/MM9_g N_BL<7>_XI0/XI53/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM6 N_XI0/XI53/XI8/NET35_XI0/XI53/XI8/MM6_d
+ N_XI0/XI53/XI8/NET36_XI0/XI53/XI8/MM6_g N_VSS_XI0/XI53/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM7 N_XI0/XI53/XI8/NET36_XI0/XI53/XI8/MM7_d
+ N_XI0/XI53/XI8/NET35_XI0/XI53/XI8/MM7_g N_VSS_XI0/XI53/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM8 N_XI0/XI53/XI8/NET35_XI0/XI53/XI8/MM8_d
+ N_WL<103>_XI0/XI53/XI8/MM8_g N_BLN<7>_XI0/XI53/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI8/MM5 N_XI0/XI53/XI8/NET34_XI0/XI53/XI8/MM5_d
+ N_XI0/XI53/XI8/NET33_XI0/XI53/XI8/MM5_g N_VDD_XI0/XI53/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI8/MM4 N_XI0/XI53/XI8/NET33_XI0/XI53/XI8/MM4_d
+ N_XI0/XI53/XI8/NET34_XI0/XI53/XI8/MM4_g N_VDD_XI0/XI53/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI8/MM10 N_XI0/XI53/XI8/NET35_XI0/XI53/XI8/MM10_d
+ N_XI0/XI53/XI8/NET36_XI0/XI53/XI8/MM10_g N_VDD_XI0/XI53/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI8/MM11 N_XI0/XI53/XI8/NET36_XI0/XI53/XI8/MM11_d
+ N_XI0/XI53/XI8/NET35_XI0/XI53/XI8/MM11_g N_VDD_XI0/XI53/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI9/MM2 N_XI0/XI53/XI9/NET34_XI0/XI53/XI9/MM2_d
+ N_XI0/XI53/XI9/NET33_XI0/XI53/XI9/MM2_g N_VSS_XI0/XI53/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM3 N_XI0/XI53/XI9/NET33_XI0/XI53/XI9/MM3_d
+ N_WL<102>_XI0/XI53/XI9/MM3_g N_BLN<6>_XI0/XI53/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM0 N_XI0/XI53/XI9/NET34_XI0/XI53/XI9/MM0_d
+ N_WL<102>_XI0/XI53/XI9/MM0_g N_BL<6>_XI0/XI53/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM1 N_XI0/XI53/XI9/NET33_XI0/XI53/XI9/MM1_d
+ N_XI0/XI53/XI9/NET34_XI0/XI53/XI9/MM1_g N_VSS_XI0/XI53/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM9 N_XI0/XI53/XI9/NET36_XI0/XI53/XI9/MM9_d
+ N_WL<103>_XI0/XI53/XI9/MM9_g N_BL<6>_XI0/XI53/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM6 N_XI0/XI53/XI9/NET35_XI0/XI53/XI9/MM6_d
+ N_XI0/XI53/XI9/NET36_XI0/XI53/XI9/MM6_g N_VSS_XI0/XI53/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM7 N_XI0/XI53/XI9/NET36_XI0/XI53/XI9/MM7_d
+ N_XI0/XI53/XI9/NET35_XI0/XI53/XI9/MM7_g N_VSS_XI0/XI53/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM8 N_XI0/XI53/XI9/NET35_XI0/XI53/XI9/MM8_d
+ N_WL<103>_XI0/XI53/XI9/MM8_g N_BLN<6>_XI0/XI53/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI9/MM5 N_XI0/XI53/XI9/NET34_XI0/XI53/XI9/MM5_d
+ N_XI0/XI53/XI9/NET33_XI0/XI53/XI9/MM5_g N_VDD_XI0/XI53/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI9/MM4 N_XI0/XI53/XI9/NET33_XI0/XI53/XI9/MM4_d
+ N_XI0/XI53/XI9/NET34_XI0/XI53/XI9/MM4_g N_VDD_XI0/XI53/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI9/MM10 N_XI0/XI53/XI9/NET35_XI0/XI53/XI9/MM10_d
+ N_XI0/XI53/XI9/NET36_XI0/XI53/XI9/MM10_g N_VDD_XI0/XI53/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI9/MM11 N_XI0/XI53/XI9/NET36_XI0/XI53/XI9/MM11_d
+ N_XI0/XI53/XI9/NET35_XI0/XI53/XI9/MM11_g N_VDD_XI0/XI53/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI10/MM2 N_XI0/XI53/XI10/NET34_XI0/XI53/XI10/MM2_d
+ N_XI0/XI53/XI10/NET33_XI0/XI53/XI10/MM2_g N_VSS_XI0/XI53/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM3 N_XI0/XI53/XI10/NET33_XI0/XI53/XI10/MM3_d
+ N_WL<102>_XI0/XI53/XI10/MM3_g N_BLN<5>_XI0/XI53/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM0 N_XI0/XI53/XI10/NET34_XI0/XI53/XI10/MM0_d
+ N_WL<102>_XI0/XI53/XI10/MM0_g N_BL<5>_XI0/XI53/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM1 N_XI0/XI53/XI10/NET33_XI0/XI53/XI10/MM1_d
+ N_XI0/XI53/XI10/NET34_XI0/XI53/XI10/MM1_g N_VSS_XI0/XI53/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM9 N_XI0/XI53/XI10/NET36_XI0/XI53/XI10/MM9_d
+ N_WL<103>_XI0/XI53/XI10/MM9_g N_BL<5>_XI0/XI53/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM6 N_XI0/XI53/XI10/NET35_XI0/XI53/XI10/MM6_d
+ N_XI0/XI53/XI10/NET36_XI0/XI53/XI10/MM6_g N_VSS_XI0/XI53/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM7 N_XI0/XI53/XI10/NET36_XI0/XI53/XI10/MM7_d
+ N_XI0/XI53/XI10/NET35_XI0/XI53/XI10/MM7_g N_VSS_XI0/XI53/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM8 N_XI0/XI53/XI10/NET35_XI0/XI53/XI10/MM8_d
+ N_WL<103>_XI0/XI53/XI10/MM8_g N_BLN<5>_XI0/XI53/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI10/MM5 N_XI0/XI53/XI10/NET34_XI0/XI53/XI10/MM5_d
+ N_XI0/XI53/XI10/NET33_XI0/XI53/XI10/MM5_g N_VDD_XI0/XI53/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI10/MM4 N_XI0/XI53/XI10/NET33_XI0/XI53/XI10/MM4_d
+ N_XI0/XI53/XI10/NET34_XI0/XI53/XI10/MM4_g N_VDD_XI0/XI53/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI10/MM10 N_XI0/XI53/XI10/NET35_XI0/XI53/XI10/MM10_d
+ N_XI0/XI53/XI10/NET36_XI0/XI53/XI10/MM10_g N_VDD_XI0/XI53/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI10/MM11 N_XI0/XI53/XI10/NET36_XI0/XI53/XI10/MM11_d
+ N_XI0/XI53/XI10/NET35_XI0/XI53/XI10/MM11_g N_VDD_XI0/XI53/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI11/MM2 N_XI0/XI53/XI11/NET34_XI0/XI53/XI11/MM2_d
+ N_XI0/XI53/XI11/NET33_XI0/XI53/XI11/MM2_g N_VSS_XI0/XI53/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM3 N_XI0/XI53/XI11/NET33_XI0/XI53/XI11/MM3_d
+ N_WL<102>_XI0/XI53/XI11/MM3_g N_BLN<4>_XI0/XI53/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM0 N_XI0/XI53/XI11/NET34_XI0/XI53/XI11/MM0_d
+ N_WL<102>_XI0/XI53/XI11/MM0_g N_BL<4>_XI0/XI53/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM1 N_XI0/XI53/XI11/NET33_XI0/XI53/XI11/MM1_d
+ N_XI0/XI53/XI11/NET34_XI0/XI53/XI11/MM1_g N_VSS_XI0/XI53/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM9 N_XI0/XI53/XI11/NET36_XI0/XI53/XI11/MM9_d
+ N_WL<103>_XI0/XI53/XI11/MM9_g N_BL<4>_XI0/XI53/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM6 N_XI0/XI53/XI11/NET35_XI0/XI53/XI11/MM6_d
+ N_XI0/XI53/XI11/NET36_XI0/XI53/XI11/MM6_g N_VSS_XI0/XI53/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM7 N_XI0/XI53/XI11/NET36_XI0/XI53/XI11/MM7_d
+ N_XI0/XI53/XI11/NET35_XI0/XI53/XI11/MM7_g N_VSS_XI0/XI53/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM8 N_XI0/XI53/XI11/NET35_XI0/XI53/XI11/MM8_d
+ N_WL<103>_XI0/XI53/XI11/MM8_g N_BLN<4>_XI0/XI53/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI11/MM5 N_XI0/XI53/XI11/NET34_XI0/XI53/XI11/MM5_d
+ N_XI0/XI53/XI11/NET33_XI0/XI53/XI11/MM5_g N_VDD_XI0/XI53/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI11/MM4 N_XI0/XI53/XI11/NET33_XI0/XI53/XI11/MM4_d
+ N_XI0/XI53/XI11/NET34_XI0/XI53/XI11/MM4_g N_VDD_XI0/XI53/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI11/MM10 N_XI0/XI53/XI11/NET35_XI0/XI53/XI11/MM10_d
+ N_XI0/XI53/XI11/NET36_XI0/XI53/XI11/MM10_g N_VDD_XI0/XI53/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI11/MM11 N_XI0/XI53/XI11/NET36_XI0/XI53/XI11/MM11_d
+ N_XI0/XI53/XI11/NET35_XI0/XI53/XI11/MM11_g N_VDD_XI0/XI53/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI12/MM2 N_XI0/XI53/XI12/NET34_XI0/XI53/XI12/MM2_d
+ N_XI0/XI53/XI12/NET33_XI0/XI53/XI12/MM2_g N_VSS_XI0/XI53/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM3 N_XI0/XI53/XI12/NET33_XI0/XI53/XI12/MM3_d
+ N_WL<102>_XI0/XI53/XI12/MM3_g N_BLN<3>_XI0/XI53/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM0 N_XI0/XI53/XI12/NET34_XI0/XI53/XI12/MM0_d
+ N_WL<102>_XI0/XI53/XI12/MM0_g N_BL<3>_XI0/XI53/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM1 N_XI0/XI53/XI12/NET33_XI0/XI53/XI12/MM1_d
+ N_XI0/XI53/XI12/NET34_XI0/XI53/XI12/MM1_g N_VSS_XI0/XI53/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM9 N_XI0/XI53/XI12/NET36_XI0/XI53/XI12/MM9_d
+ N_WL<103>_XI0/XI53/XI12/MM9_g N_BL<3>_XI0/XI53/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM6 N_XI0/XI53/XI12/NET35_XI0/XI53/XI12/MM6_d
+ N_XI0/XI53/XI12/NET36_XI0/XI53/XI12/MM6_g N_VSS_XI0/XI53/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM7 N_XI0/XI53/XI12/NET36_XI0/XI53/XI12/MM7_d
+ N_XI0/XI53/XI12/NET35_XI0/XI53/XI12/MM7_g N_VSS_XI0/XI53/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM8 N_XI0/XI53/XI12/NET35_XI0/XI53/XI12/MM8_d
+ N_WL<103>_XI0/XI53/XI12/MM8_g N_BLN<3>_XI0/XI53/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI12/MM5 N_XI0/XI53/XI12/NET34_XI0/XI53/XI12/MM5_d
+ N_XI0/XI53/XI12/NET33_XI0/XI53/XI12/MM5_g N_VDD_XI0/XI53/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI12/MM4 N_XI0/XI53/XI12/NET33_XI0/XI53/XI12/MM4_d
+ N_XI0/XI53/XI12/NET34_XI0/XI53/XI12/MM4_g N_VDD_XI0/XI53/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI12/MM10 N_XI0/XI53/XI12/NET35_XI0/XI53/XI12/MM10_d
+ N_XI0/XI53/XI12/NET36_XI0/XI53/XI12/MM10_g N_VDD_XI0/XI53/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI12/MM11 N_XI0/XI53/XI12/NET36_XI0/XI53/XI12/MM11_d
+ N_XI0/XI53/XI12/NET35_XI0/XI53/XI12/MM11_g N_VDD_XI0/XI53/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI13/MM2 N_XI0/XI53/XI13/NET34_XI0/XI53/XI13/MM2_d
+ N_XI0/XI53/XI13/NET33_XI0/XI53/XI13/MM2_g N_VSS_XI0/XI53/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM3 N_XI0/XI53/XI13/NET33_XI0/XI53/XI13/MM3_d
+ N_WL<102>_XI0/XI53/XI13/MM3_g N_BLN<2>_XI0/XI53/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM0 N_XI0/XI53/XI13/NET34_XI0/XI53/XI13/MM0_d
+ N_WL<102>_XI0/XI53/XI13/MM0_g N_BL<2>_XI0/XI53/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM1 N_XI0/XI53/XI13/NET33_XI0/XI53/XI13/MM1_d
+ N_XI0/XI53/XI13/NET34_XI0/XI53/XI13/MM1_g N_VSS_XI0/XI53/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM9 N_XI0/XI53/XI13/NET36_XI0/XI53/XI13/MM9_d
+ N_WL<103>_XI0/XI53/XI13/MM9_g N_BL<2>_XI0/XI53/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM6 N_XI0/XI53/XI13/NET35_XI0/XI53/XI13/MM6_d
+ N_XI0/XI53/XI13/NET36_XI0/XI53/XI13/MM6_g N_VSS_XI0/XI53/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM7 N_XI0/XI53/XI13/NET36_XI0/XI53/XI13/MM7_d
+ N_XI0/XI53/XI13/NET35_XI0/XI53/XI13/MM7_g N_VSS_XI0/XI53/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM8 N_XI0/XI53/XI13/NET35_XI0/XI53/XI13/MM8_d
+ N_WL<103>_XI0/XI53/XI13/MM8_g N_BLN<2>_XI0/XI53/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI13/MM5 N_XI0/XI53/XI13/NET34_XI0/XI53/XI13/MM5_d
+ N_XI0/XI53/XI13/NET33_XI0/XI53/XI13/MM5_g N_VDD_XI0/XI53/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI13/MM4 N_XI0/XI53/XI13/NET33_XI0/XI53/XI13/MM4_d
+ N_XI0/XI53/XI13/NET34_XI0/XI53/XI13/MM4_g N_VDD_XI0/XI53/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI13/MM10 N_XI0/XI53/XI13/NET35_XI0/XI53/XI13/MM10_d
+ N_XI0/XI53/XI13/NET36_XI0/XI53/XI13/MM10_g N_VDD_XI0/XI53/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI13/MM11 N_XI0/XI53/XI13/NET36_XI0/XI53/XI13/MM11_d
+ N_XI0/XI53/XI13/NET35_XI0/XI53/XI13/MM11_g N_VDD_XI0/XI53/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI14/MM2 N_XI0/XI53/XI14/NET34_XI0/XI53/XI14/MM2_d
+ N_XI0/XI53/XI14/NET33_XI0/XI53/XI14/MM2_g N_VSS_XI0/XI53/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM3 N_XI0/XI53/XI14/NET33_XI0/XI53/XI14/MM3_d
+ N_WL<102>_XI0/XI53/XI14/MM3_g N_BLN<1>_XI0/XI53/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM0 N_XI0/XI53/XI14/NET34_XI0/XI53/XI14/MM0_d
+ N_WL<102>_XI0/XI53/XI14/MM0_g N_BL<1>_XI0/XI53/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM1 N_XI0/XI53/XI14/NET33_XI0/XI53/XI14/MM1_d
+ N_XI0/XI53/XI14/NET34_XI0/XI53/XI14/MM1_g N_VSS_XI0/XI53/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM9 N_XI0/XI53/XI14/NET36_XI0/XI53/XI14/MM9_d
+ N_WL<103>_XI0/XI53/XI14/MM9_g N_BL<1>_XI0/XI53/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM6 N_XI0/XI53/XI14/NET35_XI0/XI53/XI14/MM6_d
+ N_XI0/XI53/XI14/NET36_XI0/XI53/XI14/MM6_g N_VSS_XI0/XI53/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM7 N_XI0/XI53/XI14/NET36_XI0/XI53/XI14/MM7_d
+ N_XI0/XI53/XI14/NET35_XI0/XI53/XI14/MM7_g N_VSS_XI0/XI53/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM8 N_XI0/XI53/XI14/NET35_XI0/XI53/XI14/MM8_d
+ N_WL<103>_XI0/XI53/XI14/MM8_g N_BLN<1>_XI0/XI53/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI14/MM5 N_XI0/XI53/XI14/NET34_XI0/XI53/XI14/MM5_d
+ N_XI0/XI53/XI14/NET33_XI0/XI53/XI14/MM5_g N_VDD_XI0/XI53/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI14/MM4 N_XI0/XI53/XI14/NET33_XI0/XI53/XI14/MM4_d
+ N_XI0/XI53/XI14/NET34_XI0/XI53/XI14/MM4_g N_VDD_XI0/XI53/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI14/MM10 N_XI0/XI53/XI14/NET35_XI0/XI53/XI14/MM10_d
+ N_XI0/XI53/XI14/NET36_XI0/XI53/XI14/MM10_g N_VDD_XI0/XI53/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI14/MM11 N_XI0/XI53/XI14/NET36_XI0/XI53/XI14/MM11_d
+ N_XI0/XI53/XI14/NET35_XI0/XI53/XI14/MM11_g N_VDD_XI0/XI53/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI15/MM2 N_XI0/XI53/XI15/NET34_XI0/XI53/XI15/MM2_d
+ N_XI0/XI53/XI15/NET33_XI0/XI53/XI15/MM2_g N_VSS_XI0/XI53/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM3 N_XI0/XI53/XI15/NET33_XI0/XI53/XI15/MM3_d
+ N_WL<102>_XI0/XI53/XI15/MM3_g N_BLN<0>_XI0/XI53/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM0 N_XI0/XI53/XI15/NET34_XI0/XI53/XI15/MM0_d
+ N_WL<102>_XI0/XI53/XI15/MM0_g N_BL<0>_XI0/XI53/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM1 N_XI0/XI53/XI15/NET33_XI0/XI53/XI15/MM1_d
+ N_XI0/XI53/XI15/NET34_XI0/XI53/XI15/MM1_g N_VSS_XI0/XI53/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM9 N_XI0/XI53/XI15/NET36_XI0/XI53/XI15/MM9_d
+ N_WL<103>_XI0/XI53/XI15/MM9_g N_BL<0>_XI0/XI53/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM6 N_XI0/XI53/XI15/NET35_XI0/XI53/XI15/MM6_d
+ N_XI0/XI53/XI15/NET36_XI0/XI53/XI15/MM6_g N_VSS_XI0/XI53/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM7 N_XI0/XI53/XI15/NET36_XI0/XI53/XI15/MM7_d
+ N_XI0/XI53/XI15/NET35_XI0/XI53/XI15/MM7_g N_VSS_XI0/XI53/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM8 N_XI0/XI53/XI15/NET35_XI0/XI53/XI15/MM8_d
+ N_WL<103>_XI0/XI53/XI15/MM8_g N_BLN<0>_XI0/XI53/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI53/XI15/MM5 N_XI0/XI53/XI15/NET34_XI0/XI53/XI15/MM5_d
+ N_XI0/XI53/XI15/NET33_XI0/XI53/XI15/MM5_g N_VDD_XI0/XI53/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI15/MM4 N_XI0/XI53/XI15/NET33_XI0/XI53/XI15/MM4_d
+ N_XI0/XI53/XI15/NET34_XI0/XI53/XI15/MM4_g N_VDD_XI0/XI53/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI15/MM10 N_XI0/XI53/XI15/NET35_XI0/XI53/XI15/MM10_d
+ N_XI0/XI53/XI15/NET36_XI0/XI53/XI15/MM10_g N_VDD_XI0/XI53/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI53/XI15/MM11 N_XI0/XI53/XI15/NET36_XI0/XI53/XI15/MM11_d
+ N_XI0/XI53/XI15/NET35_XI0/XI53/XI15/MM11_g N_VDD_XI0/XI53/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI0/MM2 N_XI0/XI54/XI0/NET34_XI0/XI54/XI0/MM2_d
+ N_XI0/XI54/XI0/NET33_XI0/XI54/XI0/MM2_g N_VSS_XI0/XI54/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM3 N_XI0/XI54/XI0/NET33_XI0/XI54/XI0/MM3_d
+ N_WL<104>_XI0/XI54/XI0/MM3_g N_BLN<15>_XI0/XI54/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM0 N_XI0/XI54/XI0/NET34_XI0/XI54/XI0/MM0_d
+ N_WL<104>_XI0/XI54/XI0/MM0_g N_BL<15>_XI0/XI54/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM1 N_XI0/XI54/XI0/NET33_XI0/XI54/XI0/MM1_d
+ N_XI0/XI54/XI0/NET34_XI0/XI54/XI0/MM1_g N_VSS_XI0/XI54/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM9 N_XI0/XI54/XI0/NET36_XI0/XI54/XI0/MM9_d
+ N_WL<105>_XI0/XI54/XI0/MM9_g N_BL<15>_XI0/XI54/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM6 N_XI0/XI54/XI0/NET35_XI0/XI54/XI0/MM6_d
+ N_XI0/XI54/XI0/NET36_XI0/XI54/XI0/MM6_g N_VSS_XI0/XI54/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM7 N_XI0/XI54/XI0/NET36_XI0/XI54/XI0/MM7_d
+ N_XI0/XI54/XI0/NET35_XI0/XI54/XI0/MM7_g N_VSS_XI0/XI54/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM8 N_XI0/XI54/XI0/NET35_XI0/XI54/XI0/MM8_d
+ N_WL<105>_XI0/XI54/XI0/MM8_g N_BLN<15>_XI0/XI54/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI0/MM5 N_XI0/XI54/XI0/NET34_XI0/XI54/XI0/MM5_d
+ N_XI0/XI54/XI0/NET33_XI0/XI54/XI0/MM5_g N_VDD_XI0/XI54/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI0/MM4 N_XI0/XI54/XI0/NET33_XI0/XI54/XI0/MM4_d
+ N_XI0/XI54/XI0/NET34_XI0/XI54/XI0/MM4_g N_VDD_XI0/XI54/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI0/MM10 N_XI0/XI54/XI0/NET35_XI0/XI54/XI0/MM10_d
+ N_XI0/XI54/XI0/NET36_XI0/XI54/XI0/MM10_g N_VDD_XI0/XI54/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI0/MM11 N_XI0/XI54/XI0/NET36_XI0/XI54/XI0/MM11_d
+ N_XI0/XI54/XI0/NET35_XI0/XI54/XI0/MM11_g N_VDD_XI0/XI54/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI1/MM2 N_XI0/XI54/XI1/NET34_XI0/XI54/XI1/MM2_d
+ N_XI0/XI54/XI1/NET33_XI0/XI54/XI1/MM2_g N_VSS_XI0/XI54/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM3 N_XI0/XI54/XI1/NET33_XI0/XI54/XI1/MM3_d
+ N_WL<104>_XI0/XI54/XI1/MM3_g N_BLN<14>_XI0/XI54/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM0 N_XI0/XI54/XI1/NET34_XI0/XI54/XI1/MM0_d
+ N_WL<104>_XI0/XI54/XI1/MM0_g N_BL<14>_XI0/XI54/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM1 N_XI0/XI54/XI1/NET33_XI0/XI54/XI1/MM1_d
+ N_XI0/XI54/XI1/NET34_XI0/XI54/XI1/MM1_g N_VSS_XI0/XI54/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM9 N_XI0/XI54/XI1/NET36_XI0/XI54/XI1/MM9_d
+ N_WL<105>_XI0/XI54/XI1/MM9_g N_BL<14>_XI0/XI54/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM6 N_XI0/XI54/XI1/NET35_XI0/XI54/XI1/MM6_d
+ N_XI0/XI54/XI1/NET36_XI0/XI54/XI1/MM6_g N_VSS_XI0/XI54/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM7 N_XI0/XI54/XI1/NET36_XI0/XI54/XI1/MM7_d
+ N_XI0/XI54/XI1/NET35_XI0/XI54/XI1/MM7_g N_VSS_XI0/XI54/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM8 N_XI0/XI54/XI1/NET35_XI0/XI54/XI1/MM8_d
+ N_WL<105>_XI0/XI54/XI1/MM8_g N_BLN<14>_XI0/XI54/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI1/MM5 N_XI0/XI54/XI1/NET34_XI0/XI54/XI1/MM5_d
+ N_XI0/XI54/XI1/NET33_XI0/XI54/XI1/MM5_g N_VDD_XI0/XI54/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI1/MM4 N_XI0/XI54/XI1/NET33_XI0/XI54/XI1/MM4_d
+ N_XI0/XI54/XI1/NET34_XI0/XI54/XI1/MM4_g N_VDD_XI0/XI54/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI1/MM10 N_XI0/XI54/XI1/NET35_XI0/XI54/XI1/MM10_d
+ N_XI0/XI54/XI1/NET36_XI0/XI54/XI1/MM10_g N_VDD_XI0/XI54/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI1/MM11 N_XI0/XI54/XI1/NET36_XI0/XI54/XI1/MM11_d
+ N_XI0/XI54/XI1/NET35_XI0/XI54/XI1/MM11_g N_VDD_XI0/XI54/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI2/MM2 N_XI0/XI54/XI2/NET34_XI0/XI54/XI2/MM2_d
+ N_XI0/XI54/XI2/NET33_XI0/XI54/XI2/MM2_g N_VSS_XI0/XI54/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM3 N_XI0/XI54/XI2/NET33_XI0/XI54/XI2/MM3_d
+ N_WL<104>_XI0/XI54/XI2/MM3_g N_BLN<13>_XI0/XI54/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM0 N_XI0/XI54/XI2/NET34_XI0/XI54/XI2/MM0_d
+ N_WL<104>_XI0/XI54/XI2/MM0_g N_BL<13>_XI0/XI54/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM1 N_XI0/XI54/XI2/NET33_XI0/XI54/XI2/MM1_d
+ N_XI0/XI54/XI2/NET34_XI0/XI54/XI2/MM1_g N_VSS_XI0/XI54/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM9 N_XI0/XI54/XI2/NET36_XI0/XI54/XI2/MM9_d
+ N_WL<105>_XI0/XI54/XI2/MM9_g N_BL<13>_XI0/XI54/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM6 N_XI0/XI54/XI2/NET35_XI0/XI54/XI2/MM6_d
+ N_XI0/XI54/XI2/NET36_XI0/XI54/XI2/MM6_g N_VSS_XI0/XI54/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM7 N_XI0/XI54/XI2/NET36_XI0/XI54/XI2/MM7_d
+ N_XI0/XI54/XI2/NET35_XI0/XI54/XI2/MM7_g N_VSS_XI0/XI54/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM8 N_XI0/XI54/XI2/NET35_XI0/XI54/XI2/MM8_d
+ N_WL<105>_XI0/XI54/XI2/MM8_g N_BLN<13>_XI0/XI54/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI2/MM5 N_XI0/XI54/XI2/NET34_XI0/XI54/XI2/MM5_d
+ N_XI0/XI54/XI2/NET33_XI0/XI54/XI2/MM5_g N_VDD_XI0/XI54/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI2/MM4 N_XI0/XI54/XI2/NET33_XI0/XI54/XI2/MM4_d
+ N_XI0/XI54/XI2/NET34_XI0/XI54/XI2/MM4_g N_VDD_XI0/XI54/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI2/MM10 N_XI0/XI54/XI2/NET35_XI0/XI54/XI2/MM10_d
+ N_XI0/XI54/XI2/NET36_XI0/XI54/XI2/MM10_g N_VDD_XI0/XI54/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI2/MM11 N_XI0/XI54/XI2/NET36_XI0/XI54/XI2/MM11_d
+ N_XI0/XI54/XI2/NET35_XI0/XI54/XI2/MM11_g N_VDD_XI0/XI54/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI3/MM2 N_XI0/XI54/XI3/NET34_XI0/XI54/XI3/MM2_d
+ N_XI0/XI54/XI3/NET33_XI0/XI54/XI3/MM2_g N_VSS_XI0/XI54/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM3 N_XI0/XI54/XI3/NET33_XI0/XI54/XI3/MM3_d
+ N_WL<104>_XI0/XI54/XI3/MM3_g N_BLN<12>_XI0/XI54/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM0 N_XI0/XI54/XI3/NET34_XI0/XI54/XI3/MM0_d
+ N_WL<104>_XI0/XI54/XI3/MM0_g N_BL<12>_XI0/XI54/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM1 N_XI0/XI54/XI3/NET33_XI0/XI54/XI3/MM1_d
+ N_XI0/XI54/XI3/NET34_XI0/XI54/XI3/MM1_g N_VSS_XI0/XI54/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM9 N_XI0/XI54/XI3/NET36_XI0/XI54/XI3/MM9_d
+ N_WL<105>_XI0/XI54/XI3/MM9_g N_BL<12>_XI0/XI54/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM6 N_XI0/XI54/XI3/NET35_XI0/XI54/XI3/MM6_d
+ N_XI0/XI54/XI3/NET36_XI0/XI54/XI3/MM6_g N_VSS_XI0/XI54/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM7 N_XI0/XI54/XI3/NET36_XI0/XI54/XI3/MM7_d
+ N_XI0/XI54/XI3/NET35_XI0/XI54/XI3/MM7_g N_VSS_XI0/XI54/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM8 N_XI0/XI54/XI3/NET35_XI0/XI54/XI3/MM8_d
+ N_WL<105>_XI0/XI54/XI3/MM8_g N_BLN<12>_XI0/XI54/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI3/MM5 N_XI0/XI54/XI3/NET34_XI0/XI54/XI3/MM5_d
+ N_XI0/XI54/XI3/NET33_XI0/XI54/XI3/MM5_g N_VDD_XI0/XI54/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI3/MM4 N_XI0/XI54/XI3/NET33_XI0/XI54/XI3/MM4_d
+ N_XI0/XI54/XI3/NET34_XI0/XI54/XI3/MM4_g N_VDD_XI0/XI54/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI3/MM10 N_XI0/XI54/XI3/NET35_XI0/XI54/XI3/MM10_d
+ N_XI0/XI54/XI3/NET36_XI0/XI54/XI3/MM10_g N_VDD_XI0/XI54/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI3/MM11 N_XI0/XI54/XI3/NET36_XI0/XI54/XI3/MM11_d
+ N_XI0/XI54/XI3/NET35_XI0/XI54/XI3/MM11_g N_VDD_XI0/XI54/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI4/MM2 N_XI0/XI54/XI4/NET34_XI0/XI54/XI4/MM2_d
+ N_XI0/XI54/XI4/NET33_XI0/XI54/XI4/MM2_g N_VSS_XI0/XI54/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM3 N_XI0/XI54/XI4/NET33_XI0/XI54/XI4/MM3_d
+ N_WL<104>_XI0/XI54/XI4/MM3_g N_BLN<11>_XI0/XI54/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM0 N_XI0/XI54/XI4/NET34_XI0/XI54/XI4/MM0_d
+ N_WL<104>_XI0/XI54/XI4/MM0_g N_BL<11>_XI0/XI54/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM1 N_XI0/XI54/XI4/NET33_XI0/XI54/XI4/MM1_d
+ N_XI0/XI54/XI4/NET34_XI0/XI54/XI4/MM1_g N_VSS_XI0/XI54/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM9 N_XI0/XI54/XI4/NET36_XI0/XI54/XI4/MM9_d
+ N_WL<105>_XI0/XI54/XI4/MM9_g N_BL<11>_XI0/XI54/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM6 N_XI0/XI54/XI4/NET35_XI0/XI54/XI4/MM6_d
+ N_XI0/XI54/XI4/NET36_XI0/XI54/XI4/MM6_g N_VSS_XI0/XI54/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM7 N_XI0/XI54/XI4/NET36_XI0/XI54/XI4/MM7_d
+ N_XI0/XI54/XI4/NET35_XI0/XI54/XI4/MM7_g N_VSS_XI0/XI54/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM8 N_XI0/XI54/XI4/NET35_XI0/XI54/XI4/MM8_d
+ N_WL<105>_XI0/XI54/XI4/MM8_g N_BLN<11>_XI0/XI54/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI4/MM5 N_XI0/XI54/XI4/NET34_XI0/XI54/XI4/MM5_d
+ N_XI0/XI54/XI4/NET33_XI0/XI54/XI4/MM5_g N_VDD_XI0/XI54/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI4/MM4 N_XI0/XI54/XI4/NET33_XI0/XI54/XI4/MM4_d
+ N_XI0/XI54/XI4/NET34_XI0/XI54/XI4/MM4_g N_VDD_XI0/XI54/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI4/MM10 N_XI0/XI54/XI4/NET35_XI0/XI54/XI4/MM10_d
+ N_XI0/XI54/XI4/NET36_XI0/XI54/XI4/MM10_g N_VDD_XI0/XI54/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI4/MM11 N_XI0/XI54/XI4/NET36_XI0/XI54/XI4/MM11_d
+ N_XI0/XI54/XI4/NET35_XI0/XI54/XI4/MM11_g N_VDD_XI0/XI54/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI5/MM2 N_XI0/XI54/XI5/NET34_XI0/XI54/XI5/MM2_d
+ N_XI0/XI54/XI5/NET33_XI0/XI54/XI5/MM2_g N_VSS_XI0/XI54/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM3 N_XI0/XI54/XI5/NET33_XI0/XI54/XI5/MM3_d
+ N_WL<104>_XI0/XI54/XI5/MM3_g N_BLN<10>_XI0/XI54/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM0 N_XI0/XI54/XI5/NET34_XI0/XI54/XI5/MM0_d
+ N_WL<104>_XI0/XI54/XI5/MM0_g N_BL<10>_XI0/XI54/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM1 N_XI0/XI54/XI5/NET33_XI0/XI54/XI5/MM1_d
+ N_XI0/XI54/XI5/NET34_XI0/XI54/XI5/MM1_g N_VSS_XI0/XI54/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM9 N_XI0/XI54/XI5/NET36_XI0/XI54/XI5/MM9_d
+ N_WL<105>_XI0/XI54/XI5/MM9_g N_BL<10>_XI0/XI54/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM6 N_XI0/XI54/XI5/NET35_XI0/XI54/XI5/MM6_d
+ N_XI0/XI54/XI5/NET36_XI0/XI54/XI5/MM6_g N_VSS_XI0/XI54/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM7 N_XI0/XI54/XI5/NET36_XI0/XI54/XI5/MM7_d
+ N_XI0/XI54/XI5/NET35_XI0/XI54/XI5/MM7_g N_VSS_XI0/XI54/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM8 N_XI0/XI54/XI5/NET35_XI0/XI54/XI5/MM8_d
+ N_WL<105>_XI0/XI54/XI5/MM8_g N_BLN<10>_XI0/XI54/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI5/MM5 N_XI0/XI54/XI5/NET34_XI0/XI54/XI5/MM5_d
+ N_XI0/XI54/XI5/NET33_XI0/XI54/XI5/MM5_g N_VDD_XI0/XI54/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI5/MM4 N_XI0/XI54/XI5/NET33_XI0/XI54/XI5/MM4_d
+ N_XI0/XI54/XI5/NET34_XI0/XI54/XI5/MM4_g N_VDD_XI0/XI54/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI5/MM10 N_XI0/XI54/XI5/NET35_XI0/XI54/XI5/MM10_d
+ N_XI0/XI54/XI5/NET36_XI0/XI54/XI5/MM10_g N_VDD_XI0/XI54/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI5/MM11 N_XI0/XI54/XI5/NET36_XI0/XI54/XI5/MM11_d
+ N_XI0/XI54/XI5/NET35_XI0/XI54/XI5/MM11_g N_VDD_XI0/XI54/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI6/MM2 N_XI0/XI54/XI6/NET34_XI0/XI54/XI6/MM2_d
+ N_XI0/XI54/XI6/NET33_XI0/XI54/XI6/MM2_g N_VSS_XI0/XI54/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM3 N_XI0/XI54/XI6/NET33_XI0/XI54/XI6/MM3_d
+ N_WL<104>_XI0/XI54/XI6/MM3_g N_BLN<9>_XI0/XI54/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM0 N_XI0/XI54/XI6/NET34_XI0/XI54/XI6/MM0_d
+ N_WL<104>_XI0/XI54/XI6/MM0_g N_BL<9>_XI0/XI54/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM1 N_XI0/XI54/XI6/NET33_XI0/XI54/XI6/MM1_d
+ N_XI0/XI54/XI6/NET34_XI0/XI54/XI6/MM1_g N_VSS_XI0/XI54/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM9 N_XI0/XI54/XI6/NET36_XI0/XI54/XI6/MM9_d
+ N_WL<105>_XI0/XI54/XI6/MM9_g N_BL<9>_XI0/XI54/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM6 N_XI0/XI54/XI6/NET35_XI0/XI54/XI6/MM6_d
+ N_XI0/XI54/XI6/NET36_XI0/XI54/XI6/MM6_g N_VSS_XI0/XI54/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM7 N_XI0/XI54/XI6/NET36_XI0/XI54/XI6/MM7_d
+ N_XI0/XI54/XI6/NET35_XI0/XI54/XI6/MM7_g N_VSS_XI0/XI54/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM8 N_XI0/XI54/XI6/NET35_XI0/XI54/XI6/MM8_d
+ N_WL<105>_XI0/XI54/XI6/MM8_g N_BLN<9>_XI0/XI54/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI6/MM5 N_XI0/XI54/XI6/NET34_XI0/XI54/XI6/MM5_d
+ N_XI0/XI54/XI6/NET33_XI0/XI54/XI6/MM5_g N_VDD_XI0/XI54/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI6/MM4 N_XI0/XI54/XI6/NET33_XI0/XI54/XI6/MM4_d
+ N_XI0/XI54/XI6/NET34_XI0/XI54/XI6/MM4_g N_VDD_XI0/XI54/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI6/MM10 N_XI0/XI54/XI6/NET35_XI0/XI54/XI6/MM10_d
+ N_XI0/XI54/XI6/NET36_XI0/XI54/XI6/MM10_g N_VDD_XI0/XI54/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI6/MM11 N_XI0/XI54/XI6/NET36_XI0/XI54/XI6/MM11_d
+ N_XI0/XI54/XI6/NET35_XI0/XI54/XI6/MM11_g N_VDD_XI0/XI54/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI7/MM2 N_XI0/XI54/XI7/NET34_XI0/XI54/XI7/MM2_d
+ N_XI0/XI54/XI7/NET33_XI0/XI54/XI7/MM2_g N_VSS_XI0/XI54/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM3 N_XI0/XI54/XI7/NET33_XI0/XI54/XI7/MM3_d
+ N_WL<104>_XI0/XI54/XI7/MM3_g N_BLN<8>_XI0/XI54/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM0 N_XI0/XI54/XI7/NET34_XI0/XI54/XI7/MM0_d
+ N_WL<104>_XI0/XI54/XI7/MM0_g N_BL<8>_XI0/XI54/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM1 N_XI0/XI54/XI7/NET33_XI0/XI54/XI7/MM1_d
+ N_XI0/XI54/XI7/NET34_XI0/XI54/XI7/MM1_g N_VSS_XI0/XI54/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM9 N_XI0/XI54/XI7/NET36_XI0/XI54/XI7/MM9_d
+ N_WL<105>_XI0/XI54/XI7/MM9_g N_BL<8>_XI0/XI54/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM6 N_XI0/XI54/XI7/NET35_XI0/XI54/XI7/MM6_d
+ N_XI0/XI54/XI7/NET36_XI0/XI54/XI7/MM6_g N_VSS_XI0/XI54/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM7 N_XI0/XI54/XI7/NET36_XI0/XI54/XI7/MM7_d
+ N_XI0/XI54/XI7/NET35_XI0/XI54/XI7/MM7_g N_VSS_XI0/XI54/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM8 N_XI0/XI54/XI7/NET35_XI0/XI54/XI7/MM8_d
+ N_WL<105>_XI0/XI54/XI7/MM8_g N_BLN<8>_XI0/XI54/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI7/MM5 N_XI0/XI54/XI7/NET34_XI0/XI54/XI7/MM5_d
+ N_XI0/XI54/XI7/NET33_XI0/XI54/XI7/MM5_g N_VDD_XI0/XI54/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI7/MM4 N_XI0/XI54/XI7/NET33_XI0/XI54/XI7/MM4_d
+ N_XI0/XI54/XI7/NET34_XI0/XI54/XI7/MM4_g N_VDD_XI0/XI54/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI7/MM10 N_XI0/XI54/XI7/NET35_XI0/XI54/XI7/MM10_d
+ N_XI0/XI54/XI7/NET36_XI0/XI54/XI7/MM10_g N_VDD_XI0/XI54/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI7/MM11 N_XI0/XI54/XI7/NET36_XI0/XI54/XI7/MM11_d
+ N_XI0/XI54/XI7/NET35_XI0/XI54/XI7/MM11_g N_VDD_XI0/XI54/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI8/MM2 N_XI0/XI54/XI8/NET34_XI0/XI54/XI8/MM2_d
+ N_XI0/XI54/XI8/NET33_XI0/XI54/XI8/MM2_g N_VSS_XI0/XI54/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM3 N_XI0/XI54/XI8/NET33_XI0/XI54/XI8/MM3_d
+ N_WL<104>_XI0/XI54/XI8/MM3_g N_BLN<7>_XI0/XI54/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM0 N_XI0/XI54/XI8/NET34_XI0/XI54/XI8/MM0_d
+ N_WL<104>_XI0/XI54/XI8/MM0_g N_BL<7>_XI0/XI54/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM1 N_XI0/XI54/XI8/NET33_XI0/XI54/XI8/MM1_d
+ N_XI0/XI54/XI8/NET34_XI0/XI54/XI8/MM1_g N_VSS_XI0/XI54/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM9 N_XI0/XI54/XI8/NET36_XI0/XI54/XI8/MM9_d
+ N_WL<105>_XI0/XI54/XI8/MM9_g N_BL<7>_XI0/XI54/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM6 N_XI0/XI54/XI8/NET35_XI0/XI54/XI8/MM6_d
+ N_XI0/XI54/XI8/NET36_XI0/XI54/XI8/MM6_g N_VSS_XI0/XI54/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM7 N_XI0/XI54/XI8/NET36_XI0/XI54/XI8/MM7_d
+ N_XI0/XI54/XI8/NET35_XI0/XI54/XI8/MM7_g N_VSS_XI0/XI54/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM8 N_XI0/XI54/XI8/NET35_XI0/XI54/XI8/MM8_d
+ N_WL<105>_XI0/XI54/XI8/MM8_g N_BLN<7>_XI0/XI54/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI8/MM5 N_XI0/XI54/XI8/NET34_XI0/XI54/XI8/MM5_d
+ N_XI0/XI54/XI8/NET33_XI0/XI54/XI8/MM5_g N_VDD_XI0/XI54/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI8/MM4 N_XI0/XI54/XI8/NET33_XI0/XI54/XI8/MM4_d
+ N_XI0/XI54/XI8/NET34_XI0/XI54/XI8/MM4_g N_VDD_XI0/XI54/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI8/MM10 N_XI0/XI54/XI8/NET35_XI0/XI54/XI8/MM10_d
+ N_XI0/XI54/XI8/NET36_XI0/XI54/XI8/MM10_g N_VDD_XI0/XI54/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI8/MM11 N_XI0/XI54/XI8/NET36_XI0/XI54/XI8/MM11_d
+ N_XI0/XI54/XI8/NET35_XI0/XI54/XI8/MM11_g N_VDD_XI0/XI54/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI9/MM2 N_XI0/XI54/XI9/NET34_XI0/XI54/XI9/MM2_d
+ N_XI0/XI54/XI9/NET33_XI0/XI54/XI9/MM2_g N_VSS_XI0/XI54/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM3 N_XI0/XI54/XI9/NET33_XI0/XI54/XI9/MM3_d
+ N_WL<104>_XI0/XI54/XI9/MM3_g N_BLN<6>_XI0/XI54/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM0 N_XI0/XI54/XI9/NET34_XI0/XI54/XI9/MM0_d
+ N_WL<104>_XI0/XI54/XI9/MM0_g N_BL<6>_XI0/XI54/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM1 N_XI0/XI54/XI9/NET33_XI0/XI54/XI9/MM1_d
+ N_XI0/XI54/XI9/NET34_XI0/XI54/XI9/MM1_g N_VSS_XI0/XI54/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM9 N_XI0/XI54/XI9/NET36_XI0/XI54/XI9/MM9_d
+ N_WL<105>_XI0/XI54/XI9/MM9_g N_BL<6>_XI0/XI54/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM6 N_XI0/XI54/XI9/NET35_XI0/XI54/XI9/MM6_d
+ N_XI0/XI54/XI9/NET36_XI0/XI54/XI9/MM6_g N_VSS_XI0/XI54/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM7 N_XI0/XI54/XI9/NET36_XI0/XI54/XI9/MM7_d
+ N_XI0/XI54/XI9/NET35_XI0/XI54/XI9/MM7_g N_VSS_XI0/XI54/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM8 N_XI0/XI54/XI9/NET35_XI0/XI54/XI9/MM8_d
+ N_WL<105>_XI0/XI54/XI9/MM8_g N_BLN<6>_XI0/XI54/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI9/MM5 N_XI0/XI54/XI9/NET34_XI0/XI54/XI9/MM5_d
+ N_XI0/XI54/XI9/NET33_XI0/XI54/XI9/MM5_g N_VDD_XI0/XI54/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI9/MM4 N_XI0/XI54/XI9/NET33_XI0/XI54/XI9/MM4_d
+ N_XI0/XI54/XI9/NET34_XI0/XI54/XI9/MM4_g N_VDD_XI0/XI54/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI9/MM10 N_XI0/XI54/XI9/NET35_XI0/XI54/XI9/MM10_d
+ N_XI0/XI54/XI9/NET36_XI0/XI54/XI9/MM10_g N_VDD_XI0/XI54/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI9/MM11 N_XI0/XI54/XI9/NET36_XI0/XI54/XI9/MM11_d
+ N_XI0/XI54/XI9/NET35_XI0/XI54/XI9/MM11_g N_VDD_XI0/XI54/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI10/MM2 N_XI0/XI54/XI10/NET34_XI0/XI54/XI10/MM2_d
+ N_XI0/XI54/XI10/NET33_XI0/XI54/XI10/MM2_g N_VSS_XI0/XI54/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM3 N_XI0/XI54/XI10/NET33_XI0/XI54/XI10/MM3_d
+ N_WL<104>_XI0/XI54/XI10/MM3_g N_BLN<5>_XI0/XI54/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM0 N_XI0/XI54/XI10/NET34_XI0/XI54/XI10/MM0_d
+ N_WL<104>_XI0/XI54/XI10/MM0_g N_BL<5>_XI0/XI54/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM1 N_XI0/XI54/XI10/NET33_XI0/XI54/XI10/MM1_d
+ N_XI0/XI54/XI10/NET34_XI0/XI54/XI10/MM1_g N_VSS_XI0/XI54/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM9 N_XI0/XI54/XI10/NET36_XI0/XI54/XI10/MM9_d
+ N_WL<105>_XI0/XI54/XI10/MM9_g N_BL<5>_XI0/XI54/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM6 N_XI0/XI54/XI10/NET35_XI0/XI54/XI10/MM6_d
+ N_XI0/XI54/XI10/NET36_XI0/XI54/XI10/MM6_g N_VSS_XI0/XI54/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM7 N_XI0/XI54/XI10/NET36_XI0/XI54/XI10/MM7_d
+ N_XI0/XI54/XI10/NET35_XI0/XI54/XI10/MM7_g N_VSS_XI0/XI54/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM8 N_XI0/XI54/XI10/NET35_XI0/XI54/XI10/MM8_d
+ N_WL<105>_XI0/XI54/XI10/MM8_g N_BLN<5>_XI0/XI54/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI10/MM5 N_XI0/XI54/XI10/NET34_XI0/XI54/XI10/MM5_d
+ N_XI0/XI54/XI10/NET33_XI0/XI54/XI10/MM5_g N_VDD_XI0/XI54/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI10/MM4 N_XI0/XI54/XI10/NET33_XI0/XI54/XI10/MM4_d
+ N_XI0/XI54/XI10/NET34_XI0/XI54/XI10/MM4_g N_VDD_XI0/XI54/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI10/MM10 N_XI0/XI54/XI10/NET35_XI0/XI54/XI10/MM10_d
+ N_XI0/XI54/XI10/NET36_XI0/XI54/XI10/MM10_g N_VDD_XI0/XI54/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI10/MM11 N_XI0/XI54/XI10/NET36_XI0/XI54/XI10/MM11_d
+ N_XI0/XI54/XI10/NET35_XI0/XI54/XI10/MM11_g N_VDD_XI0/XI54/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI11/MM2 N_XI0/XI54/XI11/NET34_XI0/XI54/XI11/MM2_d
+ N_XI0/XI54/XI11/NET33_XI0/XI54/XI11/MM2_g N_VSS_XI0/XI54/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM3 N_XI0/XI54/XI11/NET33_XI0/XI54/XI11/MM3_d
+ N_WL<104>_XI0/XI54/XI11/MM3_g N_BLN<4>_XI0/XI54/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM0 N_XI0/XI54/XI11/NET34_XI0/XI54/XI11/MM0_d
+ N_WL<104>_XI0/XI54/XI11/MM0_g N_BL<4>_XI0/XI54/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM1 N_XI0/XI54/XI11/NET33_XI0/XI54/XI11/MM1_d
+ N_XI0/XI54/XI11/NET34_XI0/XI54/XI11/MM1_g N_VSS_XI0/XI54/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM9 N_XI0/XI54/XI11/NET36_XI0/XI54/XI11/MM9_d
+ N_WL<105>_XI0/XI54/XI11/MM9_g N_BL<4>_XI0/XI54/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM6 N_XI0/XI54/XI11/NET35_XI0/XI54/XI11/MM6_d
+ N_XI0/XI54/XI11/NET36_XI0/XI54/XI11/MM6_g N_VSS_XI0/XI54/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM7 N_XI0/XI54/XI11/NET36_XI0/XI54/XI11/MM7_d
+ N_XI0/XI54/XI11/NET35_XI0/XI54/XI11/MM7_g N_VSS_XI0/XI54/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM8 N_XI0/XI54/XI11/NET35_XI0/XI54/XI11/MM8_d
+ N_WL<105>_XI0/XI54/XI11/MM8_g N_BLN<4>_XI0/XI54/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI11/MM5 N_XI0/XI54/XI11/NET34_XI0/XI54/XI11/MM5_d
+ N_XI0/XI54/XI11/NET33_XI0/XI54/XI11/MM5_g N_VDD_XI0/XI54/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI11/MM4 N_XI0/XI54/XI11/NET33_XI0/XI54/XI11/MM4_d
+ N_XI0/XI54/XI11/NET34_XI0/XI54/XI11/MM4_g N_VDD_XI0/XI54/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI11/MM10 N_XI0/XI54/XI11/NET35_XI0/XI54/XI11/MM10_d
+ N_XI0/XI54/XI11/NET36_XI0/XI54/XI11/MM10_g N_VDD_XI0/XI54/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI11/MM11 N_XI0/XI54/XI11/NET36_XI0/XI54/XI11/MM11_d
+ N_XI0/XI54/XI11/NET35_XI0/XI54/XI11/MM11_g N_VDD_XI0/XI54/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI12/MM2 N_XI0/XI54/XI12/NET34_XI0/XI54/XI12/MM2_d
+ N_XI0/XI54/XI12/NET33_XI0/XI54/XI12/MM2_g N_VSS_XI0/XI54/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM3 N_XI0/XI54/XI12/NET33_XI0/XI54/XI12/MM3_d
+ N_WL<104>_XI0/XI54/XI12/MM3_g N_BLN<3>_XI0/XI54/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM0 N_XI0/XI54/XI12/NET34_XI0/XI54/XI12/MM0_d
+ N_WL<104>_XI0/XI54/XI12/MM0_g N_BL<3>_XI0/XI54/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM1 N_XI0/XI54/XI12/NET33_XI0/XI54/XI12/MM1_d
+ N_XI0/XI54/XI12/NET34_XI0/XI54/XI12/MM1_g N_VSS_XI0/XI54/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM9 N_XI0/XI54/XI12/NET36_XI0/XI54/XI12/MM9_d
+ N_WL<105>_XI0/XI54/XI12/MM9_g N_BL<3>_XI0/XI54/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM6 N_XI0/XI54/XI12/NET35_XI0/XI54/XI12/MM6_d
+ N_XI0/XI54/XI12/NET36_XI0/XI54/XI12/MM6_g N_VSS_XI0/XI54/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM7 N_XI0/XI54/XI12/NET36_XI0/XI54/XI12/MM7_d
+ N_XI0/XI54/XI12/NET35_XI0/XI54/XI12/MM7_g N_VSS_XI0/XI54/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM8 N_XI0/XI54/XI12/NET35_XI0/XI54/XI12/MM8_d
+ N_WL<105>_XI0/XI54/XI12/MM8_g N_BLN<3>_XI0/XI54/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI12/MM5 N_XI0/XI54/XI12/NET34_XI0/XI54/XI12/MM5_d
+ N_XI0/XI54/XI12/NET33_XI0/XI54/XI12/MM5_g N_VDD_XI0/XI54/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI12/MM4 N_XI0/XI54/XI12/NET33_XI0/XI54/XI12/MM4_d
+ N_XI0/XI54/XI12/NET34_XI0/XI54/XI12/MM4_g N_VDD_XI0/XI54/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI12/MM10 N_XI0/XI54/XI12/NET35_XI0/XI54/XI12/MM10_d
+ N_XI0/XI54/XI12/NET36_XI0/XI54/XI12/MM10_g N_VDD_XI0/XI54/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI12/MM11 N_XI0/XI54/XI12/NET36_XI0/XI54/XI12/MM11_d
+ N_XI0/XI54/XI12/NET35_XI0/XI54/XI12/MM11_g N_VDD_XI0/XI54/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI13/MM2 N_XI0/XI54/XI13/NET34_XI0/XI54/XI13/MM2_d
+ N_XI0/XI54/XI13/NET33_XI0/XI54/XI13/MM2_g N_VSS_XI0/XI54/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM3 N_XI0/XI54/XI13/NET33_XI0/XI54/XI13/MM3_d
+ N_WL<104>_XI0/XI54/XI13/MM3_g N_BLN<2>_XI0/XI54/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM0 N_XI0/XI54/XI13/NET34_XI0/XI54/XI13/MM0_d
+ N_WL<104>_XI0/XI54/XI13/MM0_g N_BL<2>_XI0/XI54/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM1 N_XI0/XI54/XI13/NET33_XI0/XI54/XI13/MM1_d
+ N_XI0/XI54/XI13/NET34_XI0/XI54/XI13/MM1_g N_VSS_XI0/XI54/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM9 N_XI0/XI54/XI13/NET36_XI0/XI54/XI13/MM9_d
+ N_WL<105>_XI0/XI54/XI13/MM9_g N_BL<2>_XI0/XI54/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM6 N_XI0/XI54/XI13/NET35_XI0/XI54/XI13/MM6_d
+ N_XI0/XI54/XI13/NET36_XI0/XI54/XI13/MM6_g N_VSS_XI0/XI54/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM7 N_XI0/XI54/XI13/NET36_XI0/XI54/XI13/MM7_d
+ N_XI0/XI54/XI13/NET35_XI0/XI54/XI13/MM7_g N_VSS_XI0/XI54/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM8 N_XI0/XI54/XI13/NET35_XI0/XI54/XI13/MM8_d
+ N_WL<105>_XI0/XI54/XI13/MM8_g N_BLN<2>_XI0/XI54/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI13/MM5 N_XI0/XI54/XI13/NET34_XI0/XI54/XI13/MM5_d
+ N_XI0/XI54/XI13/NET33_XI0/XI54/XI13/MM5_g N_VDD_XI0/XI54/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI13/MM4 N_XI0/XI54/XI13/NET33_XI0/XI54/XI13/MM4_d
+ N_XI0/XI54/XI13/NET34_XI0/XI54/XI13/MM4_g N_VDD_XI0/XI54/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI13/MM10 N_XI0/XI54/XI13/NET35_XI0/XI54/XI13/MM10_d
+ N_XI0/XI54/XI13/NET36_XI0/XI54/XI13/MM10_g N_VDD_XI0/XI54/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI13/MM11 N_XI0/XI54/XI13/NET36_XI0/XI54/XI13/MM11_d
+ N_XI0/XI54/XI13/NET35_XI0/XI54/XI13/MM11_g N_VDD_XI0/XI54/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI14/MM2 N_XI0/XI54/XI14/NET34_XI0/XI54/XI14/MM2_d
+ N_XI0/XI54/XI14/NET33_XI0/XI54/XI14/MM2_g N_VSS_XI0/XI54/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM3 N_XI0/XI54/XI14/NET33_XI0/XI54/XI14/MM3_d
+ N_WL<104>_XI0/XI54/XI14/MM3_g N_BLN<1>_XI0/XI54/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM0 N_XI0/XI54/XI14/NET34_XI0/XI54/XI14/MM0_d
+ N_WL<104>_XI0/XI54/XI14/MM0_g N_BL<1>_XI0/XI54/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM1 N_XI0/XI54/XI14/NET33_XI0/XI54/XI14/MM1_d
+ N_XI0/XI54/XI14/NET34_XI0/XI54/XI14/MM1_g N_VSS_XI0/XI54/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM9 N_XI0/XI54/XI14/NET36_XI0/XI54/XI14/MM9_d
+ N_WL<105>_XI0/XI54/XI14/MM9_g N_BL<1>_XI0/XI54/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM6 N_XI0/XI54/XI14/NET35_XI0/XI54/XI14/MM6_d
+ N_XI0/XI54/XI14/NET36_XI0/XI54/XI14/MM6_g N_VSS_XI0/XI54/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM7 N_XI0/XI54/XI14/NET36_XI0/XI54/XI14/MM7_d
+ N_XI0/XI54/XI14/NET35_XI0/XI54/XI14/MM7_g N_VSS_XI0/XI54/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM8 N_XI0/XI54/XI14/NET35_XI0/XI54/XI14/MM8_d
+ N_WL<105>_XI0/XI54/XI14/MM8_g N_BLN<1>_XI0/XI54/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI14/MM5 N_XI0/XI54/XI14/NET34_XI0/XI54/XI14/MM5_d
+ N_XI0/XI54/XI14/NET33_XI0/XI54/XI14/MM5_g N_VDD_XI0/XI54/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI14/MM4 N_XI0/XI54/XI14/NET33_XI0/XI54/XI14/MM4_d
+ N_XI0/XI54/XI14/NET34_XI0/XI54/XI14/MM4_g N_VDD_XI0/XI54/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI14/MM10 N_XI0/XI54/XI14/NET35_XI0/XI54/XI14/MM10_d
+ N_XI0/XI54/XI14/NET36_XI0/XI54/XI14/MM10_g N_VDD_XI0/XI54/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI14/MM11 N_XI0/XI54/XI14/NET36_XI0/XI54/XI14/MM11_d
+ N_XI0/XI54/XI14/NET35_XI0/XI54/XI14/MM11_g N_VDD_XI0/XI54/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI15/MM2 N_XI0/XI54/XI15/NET34_XI0/XI54/XI15/MM2_d
+ N_XI0/XI54/XI15/NET33_XI0/XI54/XI15/MM2_g N_VSS_XI0/XI54/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM3 N_XI0/XI54/XI15/NET33_XI0/XI54/XI15/MM3_d
+ N_WL<104>_XI0/XI54/XI15/MM3_g N_BLN<0>_XI0/XI54/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM0 N_XI0/XI54/XI15/NET34_XI0/XI54/XI15/MM0_d
+ N_WL<104>_XI0/XI54/XI15/MM0_g N_BL<0>_XI0/XI54/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM1 N_XI0/XI54/XI15/NET33_XI0/XI54/XI15/MM1_d
+ N_XI0/XI54/XI15/NET34_XI0/XI54/XI15/MM1_g N_VSS_XI0/XI54/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM9 N_XI0/XI54/XI15/NET36_XI0/XI54/XI15/MM9_d
+ N_WL<105>_XI0/XI54/XI15/MM9_g N_BL<0>_XI0/XI54/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM6 N_XI0/XI54/XI15/NET35_XI0/XI54/XI15/MM6_d
+ N_XI0/XI54/XI15/NET36_XI0/XI54/XI15/MM6_g N_VSS_XI0/XI54/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM7 N_XI0/XI54/XI15/NET36_XI0/XI54/XI15/MM7_d
+ N_XI0/XI54/XI15/NET35_XI0/XI54/XI15/MM7_g N_VSS_XI0/XI54/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM8 N_XI0/XI54/XI15/NET35_XI0/XI54/XI15/MM8_d
+ N_WL<105>_XI0/XI54/XI15/MM8_g N_BLN<0>_XI0/XI54/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI54/XI15/MM5 N_XI0/XI54/XI15/NET34_XI0/XI54/XI15/MM5_d
+ N_XI0/XI54/XI15/NET33_XI0/XI54/XI15/MM5_g N_VDD_XI0/XI54/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI15/MM4 N_XI0/XI54/XI15/NET33_XI0/XI54/XI15/MM4_d
+ N_XI0/XI54/XI15/NET34_XI0/XI54/XI15/MM4_g N_VDD_XI0/XI54/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI15/MM10 N_XI0/XI54/XI15/NET35_XI0/XI54/XI15/MM10_d
+ N_XI0/XI54/XI15/NET36_XI0/XI54/XI15/MM10_g N_VDD_XI0/XI54/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI54/XI15/MM11 N_XI0/XI54/XI15/NET36_XI0/XI54/XI15/MM11_d
+ N_XI0/XI54/XI15/NET35_XI0/XI54/XI15/MM11_g N_VDD_XI0/XI54/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI0/MM2 N_XI0/XI55/XI0/NET34_XI0/XI55/XI0/MM2_d
+ N_XI0/XI55/XI0/NET33_XI0/XI55/XI0/MM2_g N_VSS_XI0/XI55/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM3 N_XI0/XI55/XI0/NET33_XI0/XI55/XI0/MM3_d
+ N_WL<106>_XI0/XI55/XI0/MM3_g N_BLN<15>_XI0/XI55/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM0 N_XI0/XI55/XI0/NET34_XI0/XI55/XI0/MM0_d
+ N_WL<106>_XI0/XI55/XI0/MM0_g N_BL<15>_XI0/XI55/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM1 N_XI0/XI55/XI0/NET33_XI0/XI55/XI0/MM1_d
+ N_XI0/XI55/XI0/NET34_XI0/XI55/XI0/MM1_g N_VSS_XI0/XI55/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM9 N_XI0/XI55/XI0/NET36_XI0/XI55/XI0/MM9_d
+ N_WL<107>_XI0/XI55/XI0/MM9_g N_BL<15>_XI0/XI55/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM6 N_XI0/XI55/XI0/NET35_XI0/XI55/XI0/MM6_d
+ N_XI0/XI55/XI0/NET36_XI0/XI55/XI0/MM6_g N_VSS_XI0/XI55/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM7 N_XI0/XI55/XI0/NET36_XI0/XI55/XI0/MM7_d
+ N_XI0/XI55/XI0/NET35_XI0/XI55/XI0/MM7_g N_VSS_XI0/XI55/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM8 N_XI0/XI55/XI0/NET35_XI0/XI55/XI0/MM8_d
+ N_WL<107>_XI0/XI55/XI0/MM8_g N_BLN<15>_XI0/XI55/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI0/MM5 N_XI0/XI55/XI0/NET34_XI0/XI55/XI0/MM5_d
+ N_XI0/XI55/XI0/NET33_XI0/XI55/XI0/MM5_g N_VDD_XI0/XI55/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI0/MM4 N_XI0/XI55/XI0/NET33_XI0/XI55/XI0/MM4_d
+ N_XI0/XI55/XI0/NET34_XI0/XI55/XI0/MM4_g N_VDD_XI0/XI55/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI0/MM10 N_XI0/XI55/XI0/NET35_XI0/XI55/XI0/MM10_d
+ N_XI0/XI55/XI0/NET36_XI0/XI55/XI0/MM10_g N_VDD_XI0/XI55/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI0/MM11 N_XI0/XI55/XI0/NET36_XI0/XI55/XI0/MM11_d
+ N_XI0/XI55/XI0/NET35_XI0/XI55/XI0/MM11_g N_VDD_XI0/XI55/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI1/MM2 N_XI0/XI55/XI1/NET34_XI0/XI55/XI1/MM2_d
+ N_XI0/XI55/XI1/NET33_XI0/XI55/XI1/MM2_g N_VSS_XI0/XI55/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM3 N_XI0/XI55/XI1/NET33_XI0/XI55/XI1/MM3_d
+ N_WL<106>_XI0/XI55/XI1/MM3_g N_BLN<14>_XI0/XI55/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM0 N_XI0/XI55/XI1/NET34_XI0/XI55/XI1/MM0_d
+ N_WL<106>_XI0/XI55/XI1/MM0_g N_BL<14>_XI0/XI55/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM1 N_XI0/XI55/XI1/NET33_XI0/XI55/XI1/MM1_d
+ N_XI0/XI55/XI1/NET34_XI0/XI55/XI1/MM1_g N_VSS_XI0/XI55/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM9 N_XI0/XI55/XI1/NET36_XI0/XI55/XI1/MM9_d
+ N_WL<107>_XI0/XI55/XI1/MM9_g N_BL<14>_XI0/XI55/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM6 N_XI0/XI55/XI1/NET35_XI0/XI55/XI1/MM6_d
+ N_XI0/XI55/XI1/NET36_XI0/XI55/XI1/MM6_g N_VSS_XI0/XI55/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM7 N_XI0/XI55/XI1/NET36_XI0/XI55/XI1/MM7_d
+ N_XI0/XI55/XI1/NET35_XI0/XI55/XI1/MM7_g N_VSS_XI0/XI55/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM8 N_XI0/XI55/XI1/NET35_XI0/XI55/XI1/MM8_d
+ N_WL<107>_XI0/XI55/XI1/MM8_g N_BLN<14>_XI0/XI55/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI1/MM5 N_XI0/XI55/XI1/NET34_XI0/XI55/XI1/MM5_d
+ N_XI0/XI55/XI1/NET33_XI0/XI55/XI1/MM5_g N_VDD_XI0/XI55/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI1/MM4 N_XI0/XI55/XI1/NET33_XI0/XI55/XI1/MM4_d
+ N_XI0/XI55/XI1/NET34_XI0/XI55/XI1/MM4_g N_VDD_XI0/XI55/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI1/MM10 N_XI0/XI55/XI1/NET35_XI0/XI55/XI1/MM10_d
+ N_XI0/XI55/XI1/NET36_XI0/XI55/XI1/MM10_g N_VDD_XI0/XI55/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI1/MM11 N_XI0/XI55/XI1/NET36_XI0/XI55/XI1/MM11_d
+ N_XI0/XI55/XI1/NET35_XI0/XI55/XI1/MM11_g N_VDD_XI0/XI55/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI2/MM2 N_XI0/XI55/XI2/NET34_XI0/XI55/XI2/MM2_d
+ N_XI0/XI55/XI2/NET33_XI0/XI55/XI2/MM2_g N_VSS_XI0/XI55/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM3 N_XI0/XI55/XI2/NET33_XI0/XI55/XI2/MM3_d
+ N_WL<106>_XI0/XI55/XI2/MM3_g N_BLN<13>_XI0/XI55/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM0 N_XI0/XI55/XI2/NET34_XI0/XI55/XI2/MM0_d
+ N_WL<106>_XI0/XI55/XI2/MM0_g N_BL<13>_XI0/XI55/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM1 N_XI0/XI55/XI2/NET33_XI0/XI55/XI2/MM1_d
+ N_XI0/XI55/XI2/NET34_XI0/XI55/XI2/MM1_g N_VSS_XI0/XI55/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM9 N_XI0/XI55/XI2/NET36_XI0/XI55/XI2/MM9_d
+ N_WL<107>_XI0/XI55/XI2/MM9_g N_BL<13>_XI0/XI55/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM6 N_XI0/XI55/XI2/NET35_XI0/XI55/XI2/MM6_d
+ N_XI0/XI55/XI2/NET36_XI0/XI55/XI2/MM6_g N_VSS_XI0/XI55/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM7 N_XI0/XI55/XI2/NET36_XI0/XI55/XI2/MM7_d
+ N_XI0/XI55/XI2/NET35_XI0/XI55/XI2/MM7_g N_VSS_XI0/XI55/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM8 N_XI0/XI55/XI2/NET35_XI0/XI55/XI2/MM8_d
+ N_WL<107>_XI0/XI55/XI2/MM8_g N_BLN<13>_XI0/XI55/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI2/MM5 N_XI0/XI55/XI2/NET34_XI0/XI55/XI2/MM5_d
+ N_XI0/XI55/XI2/NET33_XI0/XI55/XI2/MM5_g N_VDD_XI0/XI55/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI2/MM4 N_XI0/XI55/XI2/NET33_XI0/XI55/XI2/MM4_d
+ N_XI0/XI55/XI2/NET34_XI0/XI55/XI2/MM4_g N_VDD_XI0/XI55/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI2/MM10 N_XI0/XI55/XI2/NET35_XI0/XI55/XI2/MM10_d
+ N_XI0/XI55/XI2/NET36_XI0/XI55/XI2/MM10_g N_VDD_XI0/XI55/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI2/MM11 N_XI0/XI55/XI2/NET36_XI0/XI55/XI2/MM11_d
+ N_XI0/XI55/XI2/NET35_XI0/XI55/XI2/MM11_g N_VDD_XI0/XI55/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI3/MM2 N_XI0/XI55/XI3/NET34_XI0/XI55/XI3/MM2_d
+ N_XI0/XI55/XI3/NET33_XI0/XI55/XI3/MM2_g N_VSS_XI0/XI55/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM3 N_XI0/XI55/XI3/NET33_XI0/XI55/XI3/MM3_d
+ N_WL<106>_XI0/XI55/XI3/MM3_g N_BLN<12>_XI0/XI55/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM0 N_XI0/XI55/XI3/NET34_XI0/XI55/XI3/MM0_d
+ N_WL<106>_XI0/XI55/XI3/MM0_g N_BL<12>_XI0/XI55/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM1 N_XI0/XI55/XI3/NET33_XI0/XI55/XI3/MM1_d
+ N_XI0/XI55/XI3/NET34_XI0/XI55/XI3/MM1_g N_VSS_XI0/XI55/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM9 N_XI0/XI55/XI3/NET36_XI0/XI55/XI3/MM9_d
+ N_WL<107>_XI0/XI55/XI3/MM9_g N_BL<12>_XI0/XI55/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM6 N_XI0/XI55/XI3/NET35_XI0/XI55/XI3/MM6_d
+ N_XI0/XI55/XI3/NET36_XI0/XI55/XI3/MM6_g N_VSS_XI0/XI55/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM7 N_XI0/XI55/XI3/NET36_XI0/XI55/XI3/MM7_d
+ N_XI0/XI55/XI3/NET35_XI0/XI55/XI3/MM7_g N_VSS_XI0/XI55/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM8 N_XI0/XI55/XI3/NET35_XI0/XI55/XI3/MM8_d
+ N_WL<107>_XI0/XI55/XI3/MM8_g N_BLN<12>_XI0/XI55/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI3/MM5 N_XI0/XI55/XI3/NET34_XI0/XI55/XI3/MM5_d
+ N_XI0/XI55/XI3/NET33_XI0/XI55/XI3/MM5_g N_VDD_XI0/XI55/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI3/MM4 N_XI0/XI55/XI3/NET33_XI0/XI55/XI3/MM4_d
+ N_XI0/XI55/XI3/NET34_XI0/XI55/XI3/MM4_g N_VDD_XI0/XI55/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI3/MM10 N_XI0/XI55/XI3/NET35_XI0/XI55/XI3/MM10_d
+ N_XI0/XI55/XI3/NET36_XI0/XI55/XI3/MM10_g N_VDD_XI0/XI55/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI3/MM11 N_XI0/XI55/XI3/NET36_XI0/XI55/XI3/MM11_d
+ N_XI0/XI55/XI3/NET35_XI0/XI55/XI3/MM11_g N_VDD_XI0/XI55/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI4/MM2 N_XI0/XI55/XI4/NET34_XI0/XI55/XI4/MM2_d
+ N_XI0/XI55/XI4/NET33_XI0/XI55/XI4/MM2_g N_VSS_XI0/XI55/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM3 N_XI0/XI55/XI4/NET33_XI0/XI55/XI4/MM3_d
+ N_WL<106>_XI0/XI55/XI4/MM3_g N_BLN<11>_XI0/XI55/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM0 N_XI0/XI55/XI4/NET34_XI0/XI55/XI4/MM0_d
+ N_WL<106>_XI0/XI55/XI4/MM0_g N_BL<11>_XI0/XI55/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM1 N_XI0/XI55/XI4/NET33_XI0/XI55/XI4/MM1_d
+ N_XI0/XI55/XI4/NET34_XI0/XI55/XI4/MM1_g N_VSS_XI0/XI55/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM9 N_XI0/XI55/XI4/NET36_XI0/XI55/XI4/MM9_d
+ N_WL<107>_XI0/XI55/XI4/MM9_g N_BL<11>_XI0/XI55/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM6 N_XI0/XI55/XI4/NET35_XI0/XI55/XI4/MM6_d
+ N_XI0/XI55/XI4/NET36_XI0/XI55/XI4/MM6_g N_VSS_XI0/XI55/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM7 N_XI0/XI55/XI4/NET36_XI0/XI55/XI4/MM7_d
+ N_XI0/XI55/XI4/NET35_XI0/XI55/XI4/MM7_g N_VSS_XI0/XI55/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM8 N_XI0/XI55/XI4/NET35_XI0/XI55/XI4/MM8_d
+ N_WL<107>_XI0/XI55/XI4/MM8_g N_BLN<11>_XI0/XI55/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI4/MM5 N_XI0/XI55/XI4/NET34_XI0/XI55/XI4/MM5_d
+ N_XI0/XI55/XI4/NET33_XI0/XI55/XI4/MM5_g N_VDD_XI0/XI55/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI4/MM4 N_XI0/XI55/XI4/NET33_XI0/XI55/XI4/MM4_d
+ N_XI0/XI55/XI4/NET34_XI0/XI55/XI4/MM4_g N_VDD_XI0/XI55/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI4/MM10 N_XI0/XI55/XI4/NET35_XI0/XI55/XI4/MM10_d
+ N_XI0/XI55/XI4/NET36_XI0/XI55/XI4/MM10_g N_VDD_XI0/XI55/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI4/MM11 N_XI0/XI55/XI4/NET36_XI0/XI55/XI4/MM11_d
+ N_XI0/XI55/XI4/NET35_XI0/XI55/XI4/MM11_g N_VDD_XI0/XI55/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI5/MM2 N_XI0/XI55/XI5/NET34_XI0/XI55/XI5/MM2_d
+ N_XI0/XI55/XI5/NET33_XI0/XI55/XI5/MM2_g N_VSS_XI0/XI55/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM3 N_XI0/XI55/XI5/NET33_XI0/XI55/XI5/MM3_d
+ N_WL<106>_XI0/XI55/XI5/MM3_g N_BLN<10>_XI0/XI55/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM0 N_XI0/XI55/XI5/NET34_XI0/XI55/XI5/MM0_d
+ N_WL<106>_XI0/XI55/XI5/MM0_g N_BL<10>_XI0/XI55/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM1 N_XI0/XI55/XI5/NET33_XI0/XI55/XI5/MM1_d
+ N_XI0/XI55/XI5/NET34_XI0/XI55/XI5/MM1_g N_VSS_XI0/XI55/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM9 N_XI0/XI55/XI5/NET36_XI0/XI55/XI5/MM9_d
+ N_WL<107>_XI0/XI55/XI5/MM9_g N_BL<10>_XI0/XI55/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM6 N_XI0/XI55/XI5/NET35_XI0/XI55/XI5/MM6_d
+ N_XI0/XI55/XI5/NET36_XI0/XI55/XI5/MM6_g N_VSS_XI0/XI55/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM7 N_XI0/XI55/XI5/NET36_XI0/XI55/XI5/MM7_d
+ N_XI0/XI55/XI5/NET35_XI0/XI55/XI5/MM7_g N_VSS_XI0/XI55/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM8 N_XI0/XI55/XI5/NET35_XI0/XI55/XI5/MM8_d
+ N_WL<107>_XI0/XI55/XI5/MM8_g N_BLN<10>_XI0/XI55/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI5/MM5 N_XI0/XI55/XI5/NET34_XI0/XI55/XI5/MM5_d
+ N_XI0/XI55/XI5/NET33_XI0/XI55/XI5/MM5_g N_VDD_XI0/XI55/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI5/MM4 N_XI0/XI55/XI5/NET33_XI0/XI55/XI5/MM4_d
+ N_XI0/XI55/XI5/NET34_XI0/XI55/XI5/MM4_g N_VDD_XI0/XI55/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI5/MM10 N_XI0/XI55/XI5/NET35_XI0/XI55/XI5/MM10_d
+ N_XI0/XI55/XI5/NET36_XI0/XI55/XI5/MM10_g N_VDD_XI0/XI55/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI5/MM11 N_XI0/XI55/XI5/NET36_XI0/XI55/XI5/MM11_d
+ N_XI0/XI55/XI5/NET35_XI0/XI55/XI5/MM11_g N_VDD_XI0/XI55/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI6/MM2 N_XI0/XI55/XI6/NET34_XI0/XI55/XI6/MM2_d
+ N_XI0/XI55/XI6/NET33_XI0/XI55/XI6/MM2_g N_VSS_XI0/XI55/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM3 N_XI0/XI55/XI6/NET33_XI0/XI55/XI6/MM3_d
+ N_WL<106>_XI0/XI55/XI6/MM3_g N_BLN<9>_XI0/XI55/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM0 N_XI0/XI55/XI6/NET34_XI0/XI55/XI6/MM0_d
+ N_WL<106>_XI0/XI55/XI6/MM0_g N_BL<9>_XI0/XI55/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM1 N_XI0/XI55/XI6/NET33_XI0/XI55/XI6/MM1_d
+ N_XI0/XI55/XI6/NET34_XI0/XI55/XI6/MM1_g N_VSS_XI0/XI55/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM9 N_XI0/XI55/XI6/NET36_XI0/XI55/XI6/MM9_d
+ N_WL<107>_XI0/XI55/XI6/MM9_g N_BL<9>_XI0/XI55/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM6 N_XI0/XI55/XI6/NET35_XI0/XI55/XI6/MM6_d
+ N_XI0/XI55/XI6/NET36_XI0/XI55/XI6/MM6_g N_VSS_XI0/XI55/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM7 N_XI0/XI55/XI6/NET36_XI0/XI55/XI6/MM7_d
+ N_XI0/XI55/XI6/NET35_XI0/XI55/XI6/MM7_g N_VSS_XI0/XI55/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM8 N_XI0/XI55/XI6/NET35_XI0/XI55/XI6/MM8_d
+ N_WL<107>_XI0/XI55/XI6/MM8_g N_BLN<9>_XI0/XI55/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI6/MM5 N_XI0/XI55/XI6/NET34_XI0/XI55/XI6/MM5_d
+ N_XI0/XI55/XI6/NET33_XI0/XI55/XI6/MM5_g N_VDD_XI0/XI55/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI6/MM4 N_XI0/XI55/XI6/NET33_XI0/XI55/XI6/MM4_d
+ N_XI0/XI55/XI6/NET34_XI0/XI55/XI6/MM4_g N_VDD_XI0/XI55/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI6/MM10 N_XI0/XI55/XI6/NET35_XI0/XI55/XI6/MM10_d
+ N_XI0/XI55/XI6/NET36_XI0/XI55/XI6/MM10_g N_VDD_XI0/XI55/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI6/MM11 N_XI0/XI55/XI6/NET36_XI0/XI55/XI6/MM11_d
+ N_XI0/XI55/XI6/NET35_XI0/XI55/XI6/MM11_g N_VDD_XI0/XI55/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI7/MM2 N_XI0/XI55/XI7/NET34_XI0/XI55/XI7/MM2_d
+ N_XI0/XI55/XI7/NET33_XI0/XI55/XI7/MM2_g N_VSS_XI0/XI55/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM3 N_XI0/XI55/XI7/NET33_XI0/XI55/XI7/MM3_d
+ N_WL<106>_XI0/XI55/XI7/MM3_g N_BLN<8>_XI0/XI55/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM0 N_XI0/XI55/XI7/NET34_XI0/XI55/XI7/MM0_d
+ N_WL<106>_XI0/XI55/XI7/MM0_g N_BL<8>_XI0/XI55/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM1 N_XI0/XI55/XI7/NET33_XI0/XI55/XI7/MM1_d
+ N_XI0/XI55/XI7/NET34_XI0/XI55/XI7/MM1_g N_VSS_XI0/XI55/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM9 N_XI0/XI55/XI7/NET36_XI0/XI55/XI7/MM9_d
+ N_WL<107>_XI0/XI55/XI7/MM9_g N_BL<8>_XI0/XI55/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM6 N_XI0/XI55/XI7/NET35_XI0/XI55/XI7/MM6_d
+ N_XI0/XI55/XI7/NET36_XI0/XI55/XI7/MM6_g N_VSS_XI0/XI55/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM7 N_XI0/XI55/XI7/NET36_XI0/XI55/XI7/MM7_d
+ N_XI0/XI55/XI7/NET35_XI0/XI55/XI7/MM7_g N_VSS_XI0/XI55/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM8 N_XI0/XI55/XI7/NET35_XI0/XI55/XI7/MM8_d
+ N_WL<107>_XI0/XI55/XI7/MM8_g N_BLN<8>_XI0/XI55/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI7/MM5 N_XI0/XI55/XI7/NET34_XI0/XI55/XI7/MM5_d
+ N_XI0/XI55/XI7/NET33_XI0/XI55/XI7/MM5_g N_VDD_XI0/XI55/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI7/MM4 N_XI0/XI55/XI7/NET33_XI0/XI55/XI7/MM4_d
+ N_XI0/XI55/XI7/NET34_XI0/XI55/XI7/MM4_g N_VDD_XI0/XI55/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI7/MM10 N_XI0/XI55/XI7/NET35_XI0/XI55/XI7/MM10_d
+ N_XI0/XI55/XI7/NET36_XI0/XI55/XI7/MM10_g N_VDD_XI0/XI55/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI7/MM11 N_XI0/XI55/XI7/NET36_XI0/XI55/XI7/MM11_d
+ N_XI0/XI55/XI7/NET35_XI0/XI55/XI7/MM11_g N_VDD_XI0/XI55/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI8/MM2 N_XI0/XI55/XI8/NET34_XI0/XI55/XI8/MM2_d
+ N_XI0/XI55/XI8/NET33_XI0/XI55/XI8/MM2_g N_VSS_XI0/XI55/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM3 N_XI0/XI55/XI8/NET33_XI0/XI55/XI8/MM3_d
+ N_WL<106>_XI0/XI55/XI8/MM3_g N_BLN<7>_XI0/XI55/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM0 N_XI0/XI55/XI8/NET34_XI0/XI55/XI8/MM0_d
+ N_WL<106>_XI0/XI55/XI8/MM0_g N_BL<7>_XI0/XI55/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM1 N_XI0/XI55/XI8/NET33_XI0/XI55/XI8/MM1_d
+ N_XI0/XI55/XI8/NET34_XI0/XI55/XI8/MM1_g N_VSS_XI0/XI55/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM9 N_XI0/XI55/XI8/NET36_XI0/XI55/XI8/MM9_d
+ N_WL<107>_XI0/XI55/XI8/MM9_g N_BL<7>_XI0/XI55/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM6 N_XI0/XI55/XI8/NET35_XI0/XI55/XI8/MM6_d
+ N_XI0/XI55/XI8/NET36_XI0/XI55/XI8/MM6_g N_VSS_XI0/XI55/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM7 N_XI0/XI55/XI8/NET36_XI0/XI55/XI8/MM7_d
+ N_XI0/XI55/XI8/NET35_XI0/XI55/XI8/MM7_g N_VSS_XI0/XI55/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM8 N_XI0/XI55/XI8/NET35_XI0/XI55/XI8/MM8_d
+ N_WL<107>_XI0/XI55/XI8/MM8_g N_BLN<7>_XI0/XI55/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI8/MM5 N_XI0/XI55/XI8/NET34_XI0/XI55/XI8/MM5_d
+ N_XI0/XI55/XI8/NET33_XI0/XI55/XI8/MM5_g N_VDD_XI0/XI55/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI8/MM4 N_XI0/XI55/XI8/NET33_XI0/XI55/XI8/MM4_d
+ N_XI0/XI55/XI8/NET34_XI0/XI55/XI8/MM4_g N_VDD_XI0/XI55/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI8/MM10 N_XI0/XI55/XI8/NET35_XI0/XI55/XI8/MM10_d
+ N_XI0/XI55/XI8/NET36_XI0/XI55/XI8/MM10_g N_VDD_XI0/XI55/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI8/MM11 N_XI0/XI55/XI8/NET36_XI0/XI55/XI8/MM11_d
+ N_XI0/XI55/XI8/NET35_XI0/XI55/XI8/MM11_g N_VDD_XI0/XI55/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI9/MM2 N_XI0/XI55/XI9/NET34_XI0/XI55/XI9/MM2_d
+ N_XI0/XI55/XI9/NET33_XI0/XI55/XI9/MM2_g N_VSS_XI0/XI55/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM3 N_XI0/XI55/XI9/NET33_XI0/XI55/XI9/MM3_d
+ N_WL<106>_XI0/XI55/XI9/MM3_g N_BLN<6>_XI0/XI55/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM0 N_XI0/XI55/XI9/NET34_XI0/XI55/XI9/MM0_d
+ N_WL<106>_XI0/XI55/XI9/MM0_g N_BL<6>_XI0/XI55/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM1 N_XI0/XI55/XI9/NET33_XI0/XI55/XI9/MM1_d
+ N_XI0/XI55/XI9/NET34_XI0/XI55/XI9/MM1_g N_VSS_XI0/XI55/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM9 N_XI0/XI55/XI9/NET36_XI0/XI55/XI9/MM9_d
+ N_WL<107>_XI0/XI55/XI9/MM9_g N_BL<6>_XI0/XI55/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM6 N_XI0/XI55/XI9/NET35_XI0/XI55/XI9/MM6_d
+ N_XI0/XI55/XI9/NET36_XI0/XI55/XI9/MM6_g N_VSS_XI0/XI55/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM7 N_XI0/XI55/XI9/NET36_XI0/XI55/XI9/MM7_d
+ N_XI0/XI55/XI9/NET35_XI0/XI55/XI9/MM7_g N_VSS_XI0/XI55/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM8 N_XI0/XI55/XI9/NET35_XI0/XI55/XI9/MM8_d
+ N_WL<107>_XI0/XI55/XI9/MM8_g N_BLN<6>_XI0/XI55/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI9/MM5 N_XI0/XI55/XI9/NET34_XI0/XI55/XI9/MM5_d
+ N_XI0/XI55/XI9/NET33_XI0/XI55/XI9/MM5_g N_VDD_XI0/XI55/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI9/MM4 N_XI0/XI55/XI9/NET33_XI0/XI55/XI9/MM4_d
+ N_XI0/XI55/XI9/NET34_XI0/XI55/XI9/MM4_g N_VDD_XI0/XI55/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI9/MM10 N_XI0/XI55/XI9/NET35_XI0/XI55/XI9/MM10_d
+ N_XI0/XI55/XI9/NET36_XI0/XI55/XI9/MM10_g N_VDD_XI0/XI55/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI9/MM11 N_XI0/XI55/XI9/NET36_XI0/XI55/XI9/MM11_d
+ N_XI0/XI55/XI9/NET35_XI0/XI55/XI9/MM11_g N_VDD_XI0/XI55/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI10/MM2 N_XI0/XI55/XI10/NET34_XI0/XI55/XI10/MM2_d
+ N_XI0/XI55/XI10/NET33_XI0/XI55/XI10/MM2_g N_VSS_XI0/XI55/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM3 N_XI0/XI55/XI10/NET33_XI0/XI55/XI10/MM3_d
+ N_WL<106>_XI0/XI55/XI10/MM3_g N_BLN<5>_XI0/XI55/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM0 N_XI0/XI55/XI10/NET34_XI0/XI55/XI10/MM0_d
+ N_WL<106>_XI0/XI55/XI10/MM0_g N_BL<5>_XI0/XI55/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM1 N_XI0/XI55/XI10/NET33_XI0/XI55/XI10/MM1_d
+ N_XI0/XI55/XI10/NET34_XI0/XI55/XI10/MM1_g N_VSS_XI0/XI55/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM9 N_XI0/XI55/XI10/NET36_XI0/XI55/XI10/MM9_d
+ N_WL<107>_XI0/XI55/XI10/MM9_g N_BL<5>_XI0/XI55/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM6 N_XI0/XI55/XI10/NET35_XI0/XI55/XI10/MM6_d
+ N_XI0/XI55/XI10/NET36_XI0/XI55/XI10/MM6_g N_VSS_XI0/XI55/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM7 N_XI0/XI55/XI10/NET36_XI0/XI55/XI10/MM7_d
+ N_XI0/XI55/XI10/NET35_XI0/XI55/XI10/MM7_g N_VSS_XI0/XI55/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM8 N_XI0/XI55/XI10/NET35_XI0/XI55/XI10/MM8_d
+ N_WL<107>_XI0/XI55/XI10/MM8_g N_BLN<5>_XI0/XI55/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI10/MM5 N_XI0/XI55/XI10/NET34_XI0/XI55/XI10/MM5_d
+ N_XI0/XI55/XI10/NET33_XI0/XI55/XI10/MM5_g N_VDD_XI0/XI55/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI10/MM4 N_XI0/XI55/XI10/NET33_XI0/XI55/XI10/MM4_d
+ N_XI0/XI55/XI10/NET34_XI0/XI55/XI10/MM4_g N_VDD_XI0/XI55/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI10/MM10 N_XI0/XI55/XI10/NET35_XI0/XI55/XI10/MM10_d
+ N_XI0/XI55/XI10/NET36_XI0/XI55/XI10/MM10_g N_VDD_XI0/XI55/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI10/MM11 N_XI0/XI55/XI10/NET36_XI0/XI55/XI10/MM11_d
+ N_XI0/XI55/XI10/NET35_XI0/XI55/XI10/MM11_g N_VDD_XI0/XI55/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI11/MM2 N_XI0/XI55/XI11/NET34_XI0/XI55/XI11/MM2_d
+ N_XI0/XI55/XI11/NET33_XI0/XI55/XI11/MM2_g N_VSS_XI0/XI55/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM3 N_XI0/XI55/XI11/NET33_XI0/XI55/XI11/MM3_d
+ N_WL<106>_XI0/XI55/XI11/MM3_g N_BLN<4>_XI0/XI55/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM0 N_XI0/XI55/XI11/NET34_XI0/XI55/XI11/MM0_d
+ N_WL<106>_XI0/XI55/XI11/MM0_g N_BL<4>_XI0/XI55/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM1 N_XI0/XI55/XI11/NET33_XI0/XI55/XI11/MM1_d
+ N_XI0/XI55/XI11/NET34_XI0/XI55/XI11/MM1_g N_VSS_XI0/XI55/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM9 N_XI0/XI55/XI11/NET36_XI0/XI55/XI11/MM9_d
+ N_WL<107>_XI0/XI55/XI11/MM9_g N_BL<4>_XI0/XI55/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM6 N_XI0/XI55/XI11/NET35_XI0/XI55/XI11/MM6_d
+ N_XI0/XI55/XI11/NET36_XI0/XI55/XI11/MM6_g N_VSS_XI0/XI55/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM7 N_XI0/XI55/XI11/NET36_XI0/XI55/XI11/MM7_d
+ N_XI0/XI55/XI11/NET35_XI0/XI55/XI11/MM7_g N_VSS_XI0/XI55/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM8 N_XI0/XI55/XI11/NET35_XI0/XI55/XI11/MM8_d
+ N_WL<107>_XI0/XI55/XI11/MM8_g N_BLN<4>_XI0/XI55/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI11/MM5 N_XI0/XI55/XI11/NET34_XI0/XI55/XI11/MM5_d
+ N_XI0/XI55/XI11/NET33_XI0/XI55/XI11/MM5_g N_VDD_XI0/XI55/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI11/MM4 N_XI0/XI55/XI11/NET33_XI0/XI55/XI11/MM4_d
+ N_XI0/XI55/XI11/NET34_XI0/XI55/XI11/MM4_g N_VDD_XI0/XI55/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI11/MM10 N_XI0/XI55/XI11/NET35_XI0/XI55/XI11/MM10_d
+ N_XI0/XI55/XI11/NET36_XI0/XI55/XI11/MM10_g N_VDD_XI0/XI55/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI11/MM11 N_XI0/XI55/XI11/NET36_XI0/XI55/XI11/MM11_d
+ N_XI0/XI55/XI11/NET35_XI0/XI55/XI11/MM11_g N_VDD_XI0/XI55/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI12/MM2 N_XI0/XI55/XI12/NET34_XI0/XI55/XI12/MM2_d
+ N_XI0/XI55/XI12/NET33_XI0/XI55/XI12/MM2_g N_VSS_XI0/XI55/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM3 N_XI0/XI55/XI12/NET33_XI0/XI55/XI12/MM3_d
+ N_WL<106>_XI0/XI55/XI12/MM3_g N_BLN<3>_XI0/XI55/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM0 N_XI0/XI55/XI12/NET34_XI0/XI55/XI12/MM0_d
+ N_WL<106>_XI0/XI55/XI12/MM0_g N_BL<3>_XI0/XI55/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM1 N_XI0/XI55/XI12/NET33_XI0/XI55/XI12/MM1_d
+ N_XI0/XI55/XI12/NET34_XI0/XI55/XI12/MM1_g N_VSS_XI0/XI55/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM9 N_XI0/XI55/XI12/NET36_XI0/XI55/XI12/MM9_d
+ N_WL<107>_XI0/XI55/XI12/MM9_g N_BL<3>_XI0/XI55/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM6 N_XI0/XI55/XI12/NET35_XI0/XI55/XI12/MM6_d
+ N_XI0/XI55/XI12/NET36_XI0/XI55/XI12/MM6_g N_VSS_XI0/XI55/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM7 N_XI0/XI55/XI12/NET36_XI0/XI55/XI12/MM7_d
+ N_XI0/XI55/XI12/NET35_XI0/XI55/XI12/MM7_g N_VSS_XI0/XI55/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM8 N_XI0/XI55/XI12/NET35_XI0/XI55/XI12/MM8_d
+ N_WL<107>_XI0/XI55/XI12/MM8_g N_BLN<3>_XI0/XI55/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI12/MM5 N_XI0/XI55/XI12/NET34_XI0/XI55/XI12/MM5_d
+ N_XI0/XI55/XI12/NET33_XI0/XI55/XI12/MM5_g N_VDD_XI0/XI55/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI12/MM4 N_XI0/XI55/XI12/NET33_XI0/XI55/XI12/MM4_d
+ N_XI0/XI55/XI12/NET34_XI0/XI55/XI12/MM4_g N_VDD_XI0/XI55/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI12/MM10 N_XI0/XI55/XI12/NET35_XI0/XI55/XI12/MM10_d
+ N_XI0/XI55/XI12/NET36_XI0/XI55/XI12/MM10_g N_VDD_XI0/XI55/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI12/MM11 N_XI0/XI55/XI12/NET36_XI0/XI55/XI12/MM11_d
+ N_XI0/XI55/XI12/NET35_XI0/XI55/XI12/MM11_g N_VDD_XI0/XI55/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI13/MM2 N_XI0/XI55/XI13/NET34_XI0/XI55/XI13/MM2_d
+ N_XI0/XI55/XI13/NET33_XI0/XI55/XI13/MM2_g N_VSS_XI0/XI55/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM3 N_XI0/XI55/XI13/NET33_XI0/XI55/XI13/MM3_d
+ N_WL<106>_XI0/XI55/XI13/MM3_g N_BLN<2>_XI0/XI55/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM0 N_XI0/XI55/XI13/NET34_XI0/XI55/XI13/MM0_d
+ N_WL<106>_XI0/XI55/XI13/MM0_g N_BL<2>_XI0/XI55/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM1 N_XI0/XI55/XI13/NET33_XI0/XI55/XI13/MM1_d
+ N_XI0/XI55/XI13/NET34_XI0/XI55/XI13/MM1_g N_VSS_XI0/XI55/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM9 N_XI0/XI55/XI13/NET36_XI0/XI55/XI13/MM9_d
+ N_WL<107>_XI0/XI55/XI13/MM9_g N_BL<2>_XI0/XI55/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM6 N_XI0/XI55/XI13/NET35_XI0/XI55/XI13/MM6_d
+ N_XI0/XI55/XI13/NET36_XI0/XI55/XI13/MM6_g N_VSS_XI0/XI55/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM7 N_XI0/XI55/XI13/NET36_XI0/XI55/XI13/MM7_d
+ N_XI0/XI55/XI13/NET35_XI0/XI55/XI13/MM7_g N_VSS_XI0/XI55/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM8 N_XI0/XI55/XI13/NET35_XI0/XI55/XI13/MM8_d
+ N_WL<107>_XI0/XI55/XI13/MM8_g N_BLN<2>_XI0/XI55/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI13/MM5 N_XI0/XI55/XI13/NET34_XI0/XI55/XI13/MM5_d
+ N_XI0/XI55/XI13/NET33_XI0/XI55/XI13/MM5_g N_VDD_XI0/XI55/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI13/MM4 N_XI0/XI55/XI13/NET33_XI0/XI55/XI13/MM4_d
+ N_XI0/XI55/XI13/NET34_XI0/XI55/XI13/MM4_g N_VDD_XI0/XI55/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI13/MM10 N_XI0/XI55/XI13/NET35_XI0/XI55/XI13/MM10_d
+ N_XI0/XI55/XI13/NET36_XI0/XI55/XI13/MM10_g N_VDD_XI0/XI55/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI13/MM11 N_XI0/XI55/XI13/NET36_XI0/XI55/XI13/MM11_d
+ N_XI0/XI55/XI13/NET35_XI0/XI55/XI13/MM11_g N_VDD_XI0/XI55/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI14/MM2 N_XI0/XI55/XI14/NET34_XI0/XI55/XI14/MM2_d
+ N_XI0/XI55/XI14/NET33_XI0/XI55/XI14/MM2_g N_VSS_XI0/XI55/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM3 N_XI0/XI55/XI14/NET33_XI0/XI55/XI14/MM3_d
+ N_WL<106>_XI0/XI55/XI14/MM3_g N_BLN<1>_XI0/XI55/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM0 N_XI0/XI55/XI14/NET34_XI0/XI55/XI14/MM0_d
+ N_WL<106>_XI0/XI55/XI14/MM0_g N_BL<1>_XI0/XI55/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM1 N_XI0/XI55/XI14/NET33_XI0/XI55/XI14/MM1_d
+ N_XI0/XI55/XI14/NET34_XI0/XI55/XI14/MM1_g N_VSS_XI0/XI55/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM9 N_XI0/XI55/XI14/NET36_XI0/XI55/XI14/MM9_d
+ N_WL<107>_XI0/XI55/XI14/MM9_g N_BL<1>_XI0/XI55/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM6 N_XI0/XI55/XI14/NET35_XI0/XI55/XI14/MM6_d
+ N_XI0/XI55/XI14/NET36_XI0/XI55/XI14/MM6_g N_VSS_XI0/XI55/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM7 N_XI0/XI55/XI14/NET36_XI0/XI55/XI14/MM7_d
+ N_XI0/XI55/XI14/NET35_XI0/XI55/XI14/MM7_g N_VSS_XI0/XI55/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM8 N_XI0/XI55/XI14/NET35_XI0/XI55/XI14/MM8_d
+ N_WL<107>_XI0/XI55/XI14/MM8_g N_BLN<1>_XI0/XI55/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI14/MM5 N_XI0/XI55/XI14/NET34_XI0/XI55/XI14/MM5_d
+ N_XI0/XI55/XI14/NET33_XI0/XI55/XI14/MM5_g N_VDD_XI0/XI55/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI14/MM4 N_XI0/XI55/XI14/NET33_XI0/XI55/XI14/MM4_d
+ N_XI0/XI55/XI14/NET34_XI0/XI55/XI14/MM4_g N_VDD_XI0/XI55/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI14/MM10 N_XI0/XI55/XI14/NET35_XI0/XI55/XI14/MM10_d
+ N_XI0/XI55/XI14/NET36_XI0/XI55/XI14/MM10_g N_VDD_XI0/XI55/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI14/MM11 N_XI0/XI55/XI14/NET36_XI0/XI55/XI14/MM11_d
+ N_XI0/XI55/XI14/NET35_XI0/XI55/XI14/MM11_g N_VDD_XI0/XI55/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI15/MM2 N_XI0/XI55/XI15/NET34_XI0/XI55/XI15/MM2_d
+ N_XI0/XI55/XI15/NET33_XI0/XI55/XI15/MM2_g N_VSS_XI0/XI55/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM3 N_XI0/XI55/XI15/NET33_XI0/XI55/XI15/MM3_d
+ N_WL<106>_XI0/XI55/XI15/MM3_g N_BLN<0>_XI0/XI55/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM0 N_XI0/XI55/XI15/NET34_XI0/XI55/XI15/MM0_d
+ N_WL<106>_XI0/XI55/XI15/MM0_g N_BL<0>_XI0/XI55/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM1 N_XI0/XI55/XI15/NET33_XI0/XI55/XI15/MM1_d
+ N_XI0/XI55/XI15/NET34_XI0/XI55/XI15/MM1_g N_VSS_XI0/XI55/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM9 N_XI0/XI55/XI15/NET36_XI0/XI55/XI15/MM9_d
+ N_WL<107>_XI0/XI55/XI15/MM9_g N_BL<0>_XI0/XI55/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM6 N_XI0/XI55/XI15/NET35_XI0/XI55/XI15/MM6_d
+ N_XI0/XI55/XI15/NET36_XI0/XI55/XI15/MM6_g N_VSS_XI0/XI55/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM7 N_XI0/XI55/XI15/NET36_XI0/XI55/XI15/MM7_d
+ N_XI0/XI55/XI15/NET35_XI0/XI55/XI15/MM7_g N_VSS_XI0/XI55/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM8 N_XI0/XI55/XI15/NET35_XI0/XI55/XI15/MM8_d
+ N_WL<107>_XI0/XI55/XI15/MM8_g N_BLN<0>_XI0/XI55/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI55/XI15/MM5 N_XI0/XI55/XI15/NET34_XI0/XI55/XI15/MM5_d
+ N_XI0/XI55/XI15/NET33_XI0/XI55/XI15/MM5_g N_VDD_XI0/XI55/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI15/MM4 N_XI0/XI55/XI15/NET33_XI0/XI55/XI15/MM4_d
+ N_XI0/XI55/XI15/NET34_XI0/XI55/XI15/MM4_g N_VDD_XI0/XI55/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI15/MM10 N_XI0/XI55/XI15/NET35_XI0/XI55/XI15/MM10_d
+ N_XI0/XI55/XI15/NET36_XI0/XI55/XI15/MM10_g N_VDD_XI0/XI55/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI55/XI15/MM11 N_XI0/XI55/XI15/NET36_XI0/XI55/XI15/MM11_d
+ N_XI0/XI55/XI15/NET35_XI0/XI55/XI15/MM11_g N_VDD_XI0/XI55/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI0/MM2 N_XI0/XI56/XI0/NET34_XI0/XI56/XI0/MM2_d
+ N_XI0/XI56/XI0/NET33_XI0/XI56/XI0/MM2_g N_VSS_XI0/XI56/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM3 N_XI0/XI56/XI0/NET33_XI0/XI56/XI0/MM3_d
+ N_WL<108>_XI0/XI56/XI0/MM3_g N_BLN<15>_XI0/XI56/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM0 N_XI0/XI56/XI0/NET34_XI0/XI56/XI0/MM0_d
+ N_WL<108>_XI0/XI56/XI0/MM0_g N_BL<15>_XI0/XI56/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM1 N_XI0/XI56/XI0/NET33_XI0/XI56/XI0/MM1_d
+ N_XI0/XI56/XI0/NET34_XI0/XI56/XI0/MM1_g N_VSS_XI0/XI56/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM9 N_XI0/XI56/XI0/NET36_XI0/XI56/XI0/MM9_d
+ N_WL<109>_XI0/XI56/XI0/MM9_g N_BL<15>_XI0/XI56/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM6 N_XI0/XI56/XI0/NET35_XI0/XI56/XI0/MM6_d
+ N_XI0/XI56/XI0/NET36_XI0/XI56/XI0/MM6_g N_VSS_XI0/XI56/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM7 N_XI0/XI56/XI0/NET36_XI0/XI56/XI0/MM7_d
+ N_XI0/XI56/XI0/NET35_XI0/XI56/XI0/MM7_g N_VSS_XI0/XI56/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM8 N_XI0/XI56/XI0/NET35_XI0/XI56/XI0/MM8_d
+ N_WL<109>_XI0/XI56/XI0/MM8_g N_BLN<15>_XI0/XI56/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI0/MM5 N_XI0/XI56/XI0/NET34_XI0/XI56/XI0/MM5_d
+ N_XI0/XI56/XI0/NET33_XI0/XI56/XI0/MM5_g N_VDD_XI0/XI56/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI0/MM4 N_XI0/XI56/XI0/NET33_XI0/XI56/XI0/MM4_d
+ N_XI0/XI56/XI0/NET34_XI0/XI56/XI0/MM4_g N_VDD_XI0/XI56/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI0/MM10 N_XI0/XI56/XI0/NET35_XI0/XI56/XI0/MM10_d
+ N_XI0/XI56/XI0/NET36_XI0/XI56/XI0/MM10_g N_VDD_XI0/XI56/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI0/MM11 N_XI0/XI56/XI0/NET36_XI0/XI56/XI0/MM11_d
+ N_XI0/XI56/XI0/NET35_XI0/XI56/XI0/MM11_g N_VDD_XI0/XI56/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI1/MM2 N_XI0/XI56/XI1/NET34_XI0/XI56/XI1/MM2_d
+ N_XI0/XI56/XI1/NET33_XI0/XI56/XI1/MM2_g N_VSS_XI0/XI56/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM3 N_XI0/XI56/XI1/NET33_XI0/XI56/XI1/MM3_d
+ N_WL<108>_XI0/XI56/XI1/MM3_g N_BLN<14>_XI0/XI56/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM0 N_XI0/XI56/XI1/NET34_XI0/XI56/XI1/MM0_d
+ N_WL<108>_XI0/XI56/XI1/MM0_g N_BL<14>_XI0/XI56/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM1 N_XI0/XI56/XI1/NET33_XI0/XI56/XI1/MM1_d
+ N_XI0/XI56/XI1/NET34_XI0/XI56/XI1/MM1_g N_VSS_XI0/XI56/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM9 N_XI0/XI56/XI1/NET36_XI0/XI56/XI1/MM9_d
+ N_WL<109>_XI0/XI56/XI1/MM9_g N_BL<14>_XI0/XI56/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM6 N_XI0/XI56/XI1/NET35_XI0/XI56/XI1/MM6_d
+ N_XI0/XI56/XI1/NET36_XI0/XI56/XI1/MM6_g N_VSS_XI0/XI56/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM7 N_XI0/XI56/XI1/NET36_XI0/XI56/XI1/MM7_d
+ N_XI0/XI56/XI1/NET35_XI0/XI56/XI1/MM7_g N_VSS_XI0/XI56/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM8 N_XI0/XI56/XI1/NET35_XI0/XI56/XI1/MM8_d
+ N_WL<109>_XI0/XI56/XI1/MM8_g N_BLN<14>_XI0/XI56/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI1/MM5 N_XI0/XI56/XI1/NET34_XI0/XI56/XI1/MM5_d
+ N_XI0/XI56/XI1/NET33_XI0/XI56/XI1/MM5_g N_VDD_XI0/XI56/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI1/MM4 N_XI0/XI56/XI1/NET33_XI0/XI56/XI1/MM4_d
+ N_XI0/XI56/XI1/NET34_XI0/XI56/XI1/MM4_g N_VDD_XI0/XI56/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI1/MM10 N_XI0/XI56/XI1/NET35_XI0/XI56/XI1/MM10_d
+ N_XI0/XI56/XI1/NET36_XI0/XI56/XI1/MM10_g N_VDD_XI0/XI56/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI1/MM11 N_XI0/XI56/XI1/NET36_XI0/XI56/XI1/MM11_d
+ N_XI0/XI56/XI1/NET35_XI0/XI56/XI1/MM11_g N_VDD_XI0/XI56/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI2/MM2 N_XI0/XI56/XI2/NET34_XI0/XI56/XI2/MM2_d
+ N_XI0/XI56/XI2/NET33_XI0/XI56/XI2/MM2_g N_VSS_XI0/XI56/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM3 N_XI0/XI56/XI2/NET33_XI0/XI56/XI2/MM3_d
+ N_WL<108>_XI0/XI56/XI2/MM3_g N_BLN<13>_XI0/XI56/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM0 N_XI0/XI56/XI2/NET34_XI0/XI56/XI2/MM0_d
+ N_WL<108>_XI0/XI56/XI2/MM0_g N_BL<13>_XI0/XI56/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM1 N_XI0/XI56/XI2/NET33_XI0/XI56/XI2/MM1_d
+ N_XI0/XI56/XI2/NET34_XI0/XI56/XI2/MM1_g N_VSS_XI0/XI56/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM9 N_XI0/XI56/XI2/NET36_XI0/XI56/XI2/MM9_d
+ N_WL<109>_XI0/XI56/XI2/MM9_g N_BL<13>_XI0/XI56/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM6 N_XI0/XI56/XI2/NET35_XI0/XI56/XI2/MM6_d
+ N_XI0/XI56/XI2/NET36_XI0/XI56/XI2/MM6_g N_VSS_XI0/XI56/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM7 N_XI0/XI56/XI2/NET36_XI0/XI56/XI2/MM7_d
+ N_XI0/XI56/XI2/NET35_XI0/XI56/XI2/MM7_g N_VSS_XI0/XI56/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM8 N_XI0/XI56/XI2/NET35_XI0/XI56/XI2/MM8_d
+ N_WL<109>_XI0/XI56/XI2/MM8_g N_BLN<13>_XI0/XI56/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI2/MM5 N_XI0/XI56/XI2/NET34_XI0/XI56/XI2/MM5_d
+ N_XI0/XI56/XI2/NET33_XI0/XI56/XI2/MM5_g N_VDD_XI0/XI56/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI2/MM4 N_XI0/XI56/XI2/NET33_XI0/XI56/XI2/MM4_d
+ N_XI0/XI56/XI2/NET34_XI0/XI56/XI2/MM4_g N_VDD_XI0/XI56/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI2/MM10 N_XI0/XI56/XI2/NET35_XI0/XI56/XI2/MM10_d
+ N_XI0/XI56/XI2/NET36_XI0/XI56/XI2/MM10_g N_VDD_XI0/XI56/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI2/MM11 N_XI0/XI56/XI2/NET36_XI0/XI56/XI2/MM11_d
+ N_XI0/XI56/XI2/NET35_XI0/XI56/XI2/MM11_g N_VDD_XI0/XI56/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI3/MM2 N_XI0/XI56/XI3/NET34_XI0/XI56/XI3/MM2_d
+ N_XI0/XI56/XI3/NET33_XI0/XI56/XI3/MM2_g N_VSS_XI0/XI56/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM3 N_XI0/XI56/XI3/NET33_XI0/XI56/XI3/MM3_d
+ N_WL<108>_XI0/XI56/XI3/MM3_g N_BLN<12>_XI0/XI56/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM0 N_XI0/XI56/XI3/NET34_XI0/XI56/XI3/MM0_d
+ N_WL<108>_XI0/XI56/XI3/MM0_g N_BL<12>_XI0/XI56/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM1 N_XI0/XI56/XI3/NET33_XI0/XI56/XI3/MM1_d
+ N_XI0/XI56/XI3/NET34_XI0/XI56/XI3/MM1_g N_VSS_XI0/XI56/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM9 N_XI0/XI56/XI3/NET36_XI0/XI56/XI3/MM9_d
+ N_WL<109>_XI0/XI56/XI3/MM9_g N_BL<12>_XI0/XI56/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM6 N_XI0/XI56/XI3/NET35_XI0/XI56/XI3/MM6_d
+ N_XI0/XI56/XI3/NET36_XI0/XI56/XI3/MM6_g N_VSS_XI0/XI56/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM7 N_XI0/XI56/XI3/NET36_XI0/XI56/XI3/MM7_d
+ N_XI0/XI56/XI3/NET35_XI0/XI56/XI3/MM7_g N_VSS_XI0/XI56/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM8 N_XI0/XI56/XI3/NET35_XI0/XI56/XI3/MM8_d
+ N_WL<109>_XI0/XI56/XI3/MM8_g N_BLN<12>_XI0/XI56/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI3/MM5 N_XI0/XI56/XI3/NET34_XI0/XI56/XI3/MM5_d
+ N_XI0/XI56/XI3/NET33_XI0/XI56/XI3/MM5_g N_VDD_XI0/XI56/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI3/MM4 N_XI0/XI56/XI3/NET33_XI0/XI56/XI3/MM4_d
+ N_XI0/XI56/XI3/NET34_XI0/XI56/XI3/MM4_g N_VDD_XI0/XI56/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI3/MM10 N_XI0/XI56/XI3/NET35_XI0/XI56/XI3/MM10_d
+ N_XI0/XI56/XI3/NET36_XI0/XI56/XI3/MM10_g N_VDD_XI0/XI56/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI3/MM11 N_XI0/XI56/XI3/NET36_XI0/XI56/XI3/MM11_d
+ N_XI0/XI56/XI3/NET35_XI0/XI56/XI3/MM11_g N_VDD_XI0/XI56/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI4/MM2 N_XI0/XI56/XI4/NET34_XI0/XI56/XI4/MM2_d
+ N_XI0/XI56/XI4/NET33_XI0/XI56/XI4/MM2_g N_VSS_XI0/XI56/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM3 N_XI0/XI56/XI4/NET33_XI0/XI56/XI4/MM3_d
+ N_WL<108>_XI0/XI56/XI4/MM3_g N_BLN<11>_XI0/XI56/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM0 N_XI0/XI56/XI4/NET34_XI0/XI56/XI4/MM0_d
+ N_WL<108>_XI0/XI56/XI4/MM0_g N_BL<11>_XI0/XI56/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM1 N_XI0/XI56/XI4/NET33_XI0/XI56/XI4/MM1_d
+ N_XI0/XI56/XI4/NET34_XI0/XI56/XI4/MM1_g N_VSS_XI0/XI56/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM9 N_XI0/XI56/XI4/NET36_XI0/XI56/XI4/MM9_d
+ N_WL<109>_XI0/XI56/XI4/MM9_g N_BL<11>_XI0/XI56/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM6 N_XI0/XI56/XI4/NET35_XI0/XI56/XI4/MM6_d
+ N_XI0/XI56/XI4/NET36_XI0/XI56/XI4/MM6_g N_VSS_XI0/XI56/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM7 N_XI0/XI56/XI4/NET36_XI0/XI56/XI4/MM7_d
+ N_XI0/XI56/XI4/NET35_XI0/XI56/XI4/MM7_g N_VSS_XI0/XI56/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM8 N_XI0/XI56/XI4/NET35_XI0/XI56/XI4/MM8_d
+ N_WL<109>_XI0/XI56/XI4/MM8_g N_BLN<11>_XI0/XI56/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI4/MM5 N_XI0/XI56/XI4/NET34_XI0/XI56/XI4/MM5_d
+ N_XI0/XI56/XI4/NET33_XI0/XI56/XI4/MM5_g N_VDD_XI0/XI56/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI4/MM4 N_XI0/XI56/XI4/NET33_XI0/XI56/XI4/MM4_d
+ N_XI0/XI56/XI4/NET34_XI0/XI56/XI4/MM4_g N_VDD_XI0/XI56/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI4/MM10 N_XI0/XI56/XI4/NET35_XI0/XI56/XI4/MM10_d
+ N_XI0/XI56/XI4/NET36_XI0/XI56/XI4/MM10_g N_VDD_XI0/XI56/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI4/MM11 N_XI0/XI56/XI4/NET36_XI0/XI56/XI4/MM11_d
+ N_XI0/XI56/XI4/NET35_XI0/XI56/XI4/MM11_g N_VDD_XI0/XI56/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI5/MM2 N_XI0/XI56/XI5/NET34_XI0/XI56/XI5/MM2_d
+ N_XI0/XI56/XI5/NET33_XI0/XI56/XI5/MM2_g N_VSS_XI0/XI56/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM3 N_XI0/XI56/XI5/NET33_XI0/XI56/XI5/MM3_d
+ N_WL<108>_XI0/XI56/XI5/MM3_g N_BLN<10>_XI0/XI56/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM0 N_XI0/XI56/XI5/NET34_XI0/XI56/XI5/MM0_d
+ N_WL<108>_XI0/XI56/XI5/MM0_g N_BL<10>_XI0/XI56/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM1 N_XI0/XI56/XI5/NET33_XI0/XI56/XI5/MM1_d
+ N_XI0/XI56/XI5/NET34_XI0/XI56/XI5/MM1_g N_VSS_XI0/XI56/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM9 N_XI0/XI56/XI5/NET36_XI0/XI56/XI5/MM9_d
+ N_WL<109>_XI0/XI56/XI5/MM9_g N_BL<10>_XI0/XI56/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM6 N_XI0/XI56/XI5/NET35_XI0/XI56/XI5/MM6_d
+ N_XI0/XI56/XI5/NET36_XI0/XI56/XI5/MM6_g N_VSS_XI0/XI56/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM7 N_XI0/XI56/XI5/NET36_XI0/XI56/XI5/MM7_d
+ N_XI0/XI56/XI5/NET35_XI0/XI56/XI5/MM7_g N_VSS_XI0/XI56/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM8 N_XI0/XI56/XI5/NET35_XI0/XI56/XI5/MM8_d
+ N_WL<109>_XI0/XI56/XI5/MM8_g N_BLN<10>_XI0/XI56/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI5/MM5 N_XI0/XI56/XI5/NET34_XI0/XI56/XI5/MM5_d
+ N_XI0/XI56/XI5/NET33_XI0/XI56/XI5/MM5_g N_VDD_XI0/XI56/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI5/MM4 N_XI0/XI56/XI5/NET33_XI0/XI56/XI5/MM4_d
+ N_XI0/XI56/XI5/NET34_XI0/XI56/XI5/MM4_g N_VDD_XI0/XI56/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI5/MM10 N_XI0/XI56/XI5/NET35_XI0/XI56/XI5/MM10_d
+ N_XI0/XI56/XI5/NET36_XI0/XI56/XI5/MM10_g N_VDD_XI0/XI56/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI5/MM11 N_XI0/XI56/XI5/NET36_XI0/XI56/XI5/MM11_d
+ N_XI0/XI56/XI5/NET35_XI0/XI56/XI5/MM11_g N_VDD_XI0/XI56/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI6/MM2 N_XI0/XI56/XI6/NET34_XI0/XI56/XI6/MM2_d
+ N_XI0/XI56/XI6/NET33_XI0/XI56/XI6/MM2_g N_VSS_XI0/XI56/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM3 N_XI0/XI56/XI6/NET33_XI0/XI56/XI6/MM3_d
+ N_WL<108>_XI0/XI56/XI6/MM3_g N_BLN<9>_XI0/XI56/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM0 N_XI0/XI56/XI6/NET34_XI0/XI56/XI6/MM0_d
+ N_WL<108>_XI0/XI56/XI6/MM0_g N_BL<9>_XI0/XI56/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM1 N_XI0/XI56/XI6/NET33_XI0/XI56/XI6/MM1_d
+ N_XI0/XI56/XI6/NET34_XI0/XI56/XI6/MM1_g N_VSS_XI0/XI56/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM9 N_XI0/XI56/XI6/NET36_XI0/XI56/XI6/MM9_d
+ N_WL<109>_XI0/XI56/XI6/MM9_g N_BL<9>_XI0/XI56/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM6 N_XI0/XI56/XI6/NET35_XI0/XI56/XI6/MM6_d
+ N_XI0/XI56/XI6/NET36_XI0/XI56/XI6/MM6_g N_VSS_XI0/XI56/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM7 N_XI0/XI56/XI6/NET36_XI0/XI56/XI6/MM7_d
+ N_XI0/XI56/XI6/NET35_XI0/XI56/XI6/MM7_g N_VSS_XI0/XI56/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM8 N_XI0/XI56/XI6/NET35_XI0/XI56/XI6/MM8_d
+ N_WL<109>_XI0/XI56/XI6/MM8_g N_BLN<9>_XI0/XI56/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI6/MM5 N_XI0/XI56/XI6/NET34_XI0/XI56/XI6/MM5_d
+ N_XI0/XI56/XI6/NET33_XI0/XI56/XI6/MM5_g N_VDD_XI0/XI56/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI6/MM4 N_XI0/XI56/XI6/NET33_XI0/XI56/XI6/MM4_d
+ N_XI0/XI56/XI6/NET34_XI0/XI56/XI6/MM4_g N_VDD_XI0/XI56/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI6/MM10 N_XI0/XI56/XI6/NET35_XI0/XI56/XI6/MM10_d
+ N_XI0/XI56/XI6/NET36_XI0/XI56/XI6/MM10_g N_VDD_XI0/XI56/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI6/MM11 N_XI0/XI56/XI6/NET36_XI0/XI56/XI6/MM11_d
+ N_XI0/XI56/XI6/NET35_XI0/XI56/XI6/MM11_g N_VDD_XI0/XI56/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI7/MM2 N_XI0/XI56/XI7/NET34_XI0/XI56/XI7/MM2_d
+ N_XI0/XI56/XI7/NET33_XI0/XI56/XI7/MM2_g N_VSS_XI0/XI56/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM3 N_XI0/XI56/XI7/NET33_XI0/XI56/XI7/MM3_d
+ N_WL<108>_XI0/XI56/XI7/MM3_g N_BLN<8>_XI0/XI56/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM0 N_XI0/XI56/XI7/NET34_XI0/XI56/XI7/MM0_d
+ N_WL<108>_XI0/XI56/XI7/MM0_g N_BL<8>_XI0/XI56/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM1 N_XI0/XI56/XI7/NET33_XI0/XI56/XI7/MM1_d
+ N_XI0/XI56/XI7/NET34_XI0/XI56/XI7/MM1_g N_VSS_XI0/XI56/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM9 N_XI0/XI56/XI7/NET36_XI0/XI56/XI7/MM9_d
+ N_WL<109>_XI0/XI56/XI7/MM9_g N_BL<8>_XI0/XI56/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM6 N_XI0/XI56/XI7/NET35_XI0/XI56/XI7/MM6_d
+ N_XI0/XI56/XI7/NET36_XI0/XI56/XI7/MM6_g N_VSS_XI0/XI56/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM7 N_XI0/XI56/XI7/NET36_XI0/XI56/XI7/MM7_d
+ N_XI0/XI56/XI7/NET35_XI0/XI56/XI7/MM7_g N_VSS_XI0/XI56/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM8 N_XI0/XI56/XI7/NET35_XI0/XI56/XI7/MM8_d
+ N_WL<109>_XI0/XI56/XI7/MM8_g N_BLN<8>_XI0/XI56/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI7/MM5 N_XI0/XI56/XI7/NET34_XI0/XI56/XI7/MM5_d
+ N_XI0/XI56/XI7/NET33_XI0/XI56/XI7/MM5_g N_VDD_XI0/XI56/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI7/MM4 N_XI0/XI56/XI7/NET33_XI0/XI56/XI7/MM4_d
+ N_XI0/XI56/XI7/NET34_XI0/XI56/XI7/MM4_g N_VDD_XI0/XI56/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI7/MM10 N_XI0/XI56/XI7/NET35_XI0/XI56/XI7/MM10_d
+ N_XI0/XI56/XI7/NET36_XI0/XI56/XI7/MM10_g N_VDD_XI0/XI56/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI7/MM11 N_XI0/XI56/XI7/NET36_XI0/XI56/XI7/MM11_d
+ N_XI0/XI56/XI7/NET35_XI0/XI56/XI7/MM11_g N_VDD_XI0/XI56/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI8/MM2 N_XI0/XI56/XI8/NET34_XI0/XI56/XI8/MM2_d
+ N_XI0/XI56/XI8/NET33_XI0/XI56/XI8/MM2_g N_VSS_XI0/XI56/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM3 N_XI0/XI56/XI8/NET33_XI0/XI56/XI8/MM3_d
+ N_WL<108>_XI0/XI56/XI8/MM3_g N_BLN<7>_XI0/XI56/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM0 N_XI0/XI56/XI8/NET34_XI0/XI56/XI8/MM0_d
+ N_WL<108>_XI0/XI56/XI8/MM0_g N_BL<7>_XI0/XI56/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM1 N_XI0/XI56/XI8/NET33_XI0/XI56/XI8/MM1_d
+ N_XI0/XI56/XI8/NET34_XI0/XI56/XI8/MM1_g N_VSS_XI0/XI56/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM9 N_XI0/XI56/XI8/NET36_XI0/XI56/XI8/MM9_d
+ N_WL<109>_XI0/XI56/XI8/MM9_g N_BL<7>_XI0/XI56/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM6 N_XI0/XI56/XI8/NET35_XI0/XI56/XI8/MM6_d
+ N_XI0/XI56/XI8/NET36_XI0/XI56/XI8/MM6_g N_VSS_XI0/XI56/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM7 N_XI0/XI56/XI8/NET36_XI0/XI56/XI8/MM7_d
+ N_XI0/XI56/XI8/NET35_XI0/XI56/XI8/MM7_g N_VSS_XI0/XI56/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM8 N_XI0/XI56/XI8/NET35_XI0/XI56/XI8/MM8_d
+ N_WL<109>_XI0/XI56/XI8/MM8_g N_BLN<7>_XI0/XI56/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI8/MM5 N_XI0/XI56/XI8/NET34_XI0/XI56/XI8/MM5_d
+ N_XI0/XI56/XI8/NET33_XI0/XI56/XI8/MM5_g N_VDD_XI0/XI56/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI8/MM4 N_XI0/XI56/XI8/NET33_XI0/XI56/XI8/MM4_d
+ N_XI0/XI56/XI8/NET34_XI0/XI56/XI8/MM4_g N_VDD_XI0/XI56/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI8/MM10 N_XI0/XI56/XI8/NET35_XI0/XI56/XI8/MM10_d
+ N_XI0/XI56/XI8/NET36_XI0/XI56/XI8/MM10_g N_VDD_XI0/XI56/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI8/MM11 N_XI0/XI56/XI8/NET36_XI0/XI56/XI8/MM11_d
+ N_XI0/XI56/XI8/NET35_XI0/XI56/XI8/MM11_g N_VDD_XI0/XI56/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI9/MM2 N_XI0/XI56/XI9/NET34_XI0/XI56/XI9/MM2_d
+ N_XI0/XI56/XI9/NET33_XI0/XI56/XI9/MM2_g N_VSS_XI0/XI56/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM3 N_XI0/XI56/XI9/NET33_XI0/XI56/XI9/MM3_d
+ N_WL<108>_XI0/XI56/XI9/MM3_g N_BLN<6>_XI0/XI56/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM0 N_XI0/XI56/XI9/NET34_XI0/XI56/XI9/MM0_d
+ N_WL<108>_XI0/XI56/XI9/MM0_g N_BL<6>_XI0/XI56/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM1 N_XI0/XI56/XI9/NET33_XI0/XI56/XI9/MM1_d
+ N_XI0/XI56/XI9/NET34_XI0/XI56/XI9/MM1_g N_VSS_XI0/XI56/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM9 N_XI0/XI56/XI9/NET36_XI0/XI56/XI9/MM9_d
+ N_WL<109>_XI0/XI56/XI9/MM9_g N_BL<6>_XI0/XI56/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM6 N_XI0/XI56/XI9/NET35_XI0/XI56/XI9/MM6_d
+ N_XI0/XI56/XI9/NET36_XI0/XI56/XI9/MM6_g N_VSS_XI0/XI56/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM7 N_XI0/XI56/XI9/NET36_XI0/XI56/XI9/MM7_d
+ N_XI0/XI56/XI9/NET35_XI0/XI56/XI9/MM7_g N_VSS_XI0/XI56/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM8 N_XI0/XI56/XI9/NET35_XI0/XI56/XI9/MM8_d
+ N_WL<109>_XI0/XI56/XI9/MM8_g N_BLN<6>_XI0/XI56/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI9/MM5 N_XI0/XI56/XI9/NET34_XI0/XI56/XI9/MM5_d
+ N_XI0/XI56/XI9/NET33_XI0/XI56/XI9/MM5_g N_VDD_XI0/XI56/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI9/MM4 N_XI0/XI56/XI9/NET33_XI0/XI56/XI9/MM4_d
+ N_XI0/XI56/XI9/NET34_XI0/XI56/XI9/MM4_g N_VDD_XI0/XI56/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI9/MM10 N_XI0/XI56/XI9/NET35_XI0/XI56/XI9/MM10_d
+ N_XI0/XI56/XI9/NET36_XI0/XI56/XI9/MM10_g N_VDD_XI0/XI56/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI9/MM11 N_XI0/XI56/XI9/NET36_XI0/XI56/XI9/MM11_d
+ N_XI0/XI56/XI9/NET35_XI0/XI56/XI9/MM11_g N_VDD_XI0/XI56/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI10/MM2 N_XI0/XI56/XI10/NET34_XI0/XI56/XI10/MM2_d
+ N_XI0/XI56/XI10/NET33_XI0/XI56/XI10/MM2_g N_VSS_XI0/XI56/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM3 N_XI0/XI56/XI10/NET33_XI0/XI56/XI10/MM3_d
+ N_WL<108>_XI0/XI56/XI10/MM3_g N_BLN<5>_XI0/XI56/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM0 N_XI0/XI56/XI10/NET34_XI0/XI56/XI10/MM0_d
+ N_WL<108>_XI0/XI56/XI10/MM0_g N_BL<5>_XI0/XI56/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM1 N_XI0/XI56/XI10/NET33_XI0/XI56/XI10/MM1_d
+ N_XI0/XI56/XI10/NET34_XI0/XI56/XI10/MM1_g N_VSS_XI0/XI56/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM9 N_XI0/XI56/XI10/NET36_XI0/XI56/XI10/MM9_d
+ N_WL<109>_XI0/XI56/XI10/MM9_g N_BL<5>_XI0/XI56/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM6 N_XI0/XI56/XI10/NET35_XI0/XI56/XI10/MM6_d
+ N_XI0/XI56/XI10/NET36_XI0/XI56/XI10/MM6_g N_VSS_XI0/XI56/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM7 N_XI0/XI56/XI10/NET36_XI0/XI56/XI10/MM7_d
+ N_XI0/XI56/XI10/NET35_XI0/XI56/XI10/MM7_g N_VSS_XI0/XI56/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM8 N_XI0/XI56/XI10/NET35_XI0/XI56/XI10/MM8_d
+ N_WL<109>_XI0/XI56/XI10/MM8_g N_BLN<5>_XI0/XI56/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI10/MM5 N_XI0/XI56/XI10/NET34_XI0/XI56/XI10/MM5_d
+ N_XI0/XI56/XI10/NET33_XI0/XI56/XI10/MM5_g N_VDD_XI0/XI56/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI10/MM4 N_XI0/XI56/XI10/NET33_XI0/XI56/XI10/MM4_d
+ N_XI0/XI56/XI10/NET34_XI0/XI56/XI10/MM4_g N_VDD_XI0/XI56/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI10/MM10 N_XI0/XI56/XI10/NET35_XI0/XI56/XI10/MM10_d
+ N_XI0/XI56/XI10/NET36_XI0/XI56/XI10/MM10_g N_VDD_XI0/XI56/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI10/MM11 N_XI0/XI56/XI10/NET36_XI0/XI56/XI10/MM11_d
+ N_XI0/XI56/XI10/NET35_XI0/XI56/XI10/MM11_g N_VDD_XI0/XI56/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI11/MM2 N_XI0/XI56/XI11/NET34_XI0/XI56/XI11/MM2_d
+ N_XI0/XI56/XI11/NET33_XI0/XI56/XI11/MM2_g N_VSS_XI0/XI56/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM3 N_XI0/XI56/XI11/NET33_XI0/XI56/XI11/MM3_d
+ N_WL<108>_XI0/XI56/XI11/MM3_g N_BLN<4>_XI0/XI56/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM0 N_XI0/XI56/XI11/NET34_XI0/XI56/XI11/MM0_d
+ N_WL<108>_XI0/XI56/XI11/MM0_g N_BL<4>_XI0/XI56/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM1 N_XI0/XI56/XI11/NET33_XI0/XI56/XI11/MM1_d
+ N_XI0/XI56/XI11/NET34_XI0/XI56/XI11/MM1_g N_VSS_XI0/XI56/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM9 N_XI0/XI56/XI11/NET36_XI0/XI56/XI11/MM9_d
+ N_WL<109>_XI0/XI56/XI11/MM9_g N_BL<4>_XI0/XI56/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM6 N_XI0/XI56/XI11/NET35_XI0/XI56/XI11/MM6_d
+ N_XI0/XI56/XI11/NET36_XI0/XI56/XI11/MM6_g N_VSS_XI0/XI56/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM7 N_XI0/XI56/XI11/NET36_XI0/XI56/XI11/MM7_d
+ N_XI0/XI56/XI11/NET35_XI0/XI56/XI11/MM7_g N_VSS_XI0/XI56/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM8 N_XI0/XI56/XI11/NET35_XI0/XI56/XI11/MM8_d
+ N_WL<109>_XI0/XI56/XI11/MM8_g N_BLN<4>_XI0/XI56/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI11/MM5 N_XI0/XI56/XI11/NET34_XI0/XI56/XI11/MM5_d
+ N_XI0/XI56/XI11/NET33_XI0/XI56/XI11/MM5_g N_VDD_XI0/XI56/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI11/MM4 N_XI0/XI56/XI11/NET33_XI0/XI56/XI11/MM4_d
+ N_XI0/XI56/XI11/NET34_XI0/XI56/XI11/MM4_g N_VDD_XI0/XI56/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI11/MM10 N_XI0/XI56/XI11/NET35_XI0/XI56/XI11/MM10_d
+ N_XI0/XI56/XI11/NET36_XI0/XI56/XI11/MM10_g N_VDD_XI0/XI56/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI11/MM11 N_XI0/XI56/XI11/NET36_XI0/XI56/XI11/MM11_d
+ N_XI0/XI56/XI11/NET35_XI0/XI56/XI11/MM11_g N_VDD_XI0/XI56/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI12/MM2 N_XI0/XI56/XI12/NET34_XI0/XI56/XI12/MM2_d
+ N_XI0/XI56/XI12/NET33_XI0/XI56/XI12/MM2_g N_VSS_XI0/XI56/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM3 N_XI0/XI56/XI12/NET33_XI0/XI56/XI12/MM3_d
+ N_WL<108>_XI0/XI56/XI12/MM3_g N_BLN<3>_XI0/XI56/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM0 N_XI0/XI56/XI12/NET34_XI0/XI56/XI12/MM0_d
+ N_WL<108>_XI0/XI56/XI12/MM0_g N_BL<3>_XI0/XI56/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM1 N_XI0/XI56/XI12/NET33_XI0/XI56/XI12/MM1_d
+ N_XI0/XI56/XI12/NET34_XI0/XI56/XI12/MM1_g N_VSS_XI0/XI56/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM9 N_XI0/XI56/XI12/NET36_XI0/XI56/XI12/MM9_d
+ N_WL<109>_XI0/XI56/XI12/MM9_g N_BL<3>_XI0/XI56/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM6 N_XI0/XI56/XI12/NET35_XI0/XI56/XI12/MM6_d
+ N_XI0/XI56/XI12/NET36_XI0/XI56/XI12/MM6_g N_VSS_XI0/XI56/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM7 N_XI0/XI56/XI12/NET36_XI0/XI56/XI12/MM7_d
+ N_XI0/XI56/XI12/NET35_XI0/XI56/XI12/MM7_g N_VSS_XI0/XI56/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM8 N_XI0/XI56/XI12/NET35_XI0/XI56/XI12/MM8_d
+ N_WL<109>_XI0/XI56/XI12/MM8_g N_BLN<3>_XI0/XI56/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI12/MM5 N_XI0/XI56/XI12/NET34_XI0/XI56/XI12/MM5_d
+ N_XI0/XI56/XI12/NET33_XI0/XI56/XI12/MM5_g N_VDD_XI0/XI56/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI12/MM4 N_XI0/XI56/XI12/NET33_XI0/XI56/XI12/MM4_d
+ N_XI0/XI56/XI12/NET34_XI0/XI56/XI12/MM4_g N_VDD_XI0/XI56/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI12/MM10 N_XI0/XI56/XI12/NET35_XI0/XI56/XI12/MM10_d
+ N_XI0/XI56/XI12/NET36_XI0/XI56/XI12/MM10_g N_VDD_XI0/XI56/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI12/MM11 N_XI0/XI56/XI12/NET36_XI0/XI56/XI12/MM11_d
+ N_XI0/XI56/XI12/NET35_XI0/XI56/XI12/MM11_g N_VDD_XI0/XI56/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI13/MM2 N_XI0/XI56/XI13/NET34_XI0/XI56/XI13/MM2_d
+ N_XI0/XI56/XI13/NET33_XI0/XI56/XI13/MM2_g N_VSS_XI0/XI56/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM3 N_XI0/XI56/XI13/NET33_XI0/XI56/XI13/MM3_d
+ N_WL<108>_XI0/XI56/XI13/MM3_g N_BLN<2>_XI0/XI56/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM0 N_XI0/XI56/XI13/NET34_XI0/XI56/XI13/MM0_d
+ N_WL<108>_XI0/XI56/XI13/MM0_g N_BL<2>_XI0/XI56/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM1 N_XI0/XI56/XI13/NET33_XI0/XI56/XI13/MM1_d
+ N_XI0/XI56/XI13/NET34_XI0/XI56/XI13/MM1_g N_VSS_XI0/XI56/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM9 N_XI0/XI56/XI13/NET36_XI0/XI56/XI13/MM9_d
+ N_WL<109>_XI0/XI56/XI13/MM9_g N_BL<2>_XI0/XI56/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM6 N_XI0/XI56/XI13/NET35_XI0/XI56/XI13/MM6_d
+ N_XI0/XI56/XI13/NET36_XI0/XI56/XI13/MM6_g N_VSS_XI0/XI56/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM7 N_XI0/XI56/XI13/NET36_XI0/XI56/XI13/MM7_d
+ N_XI0/XI56/XI13/NET35_XI0/XI56/XI13/MM7_g N_VSS_XI0/XI56/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM8 N_XI0/XI56/XI13/NET35_XI0/XI56/XI13/MM8_d
+ N_WL<109>_XI0/XI56/XI13/MM8_g N_BLN<2>_XI0/XI56/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI13/MM5 N_XI0/XI56/XI13/NET34_XI0/XI56/XI13/MM5_d
+ N_XI0/XI56/XI13/NET33_XI0/XI56/XI13/MM5_g N_VDD_XI0/XI56/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI13/MM4 N_XI0/XI56/XI13/NET33_XI0/XI56/XI13/MM4_d
+ N_XI0/XI56/XI13/NET34_XI0/XI56/XI13/MM4_g N_VDD_XI0/XI56/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI13/MM10 N_XI0/XI56/XI13/NET35_XI0/XI56/XI13/MM10_d
+ N_XI0/XI56/XI13/NET36_XI0/XI56/XI13/MM10_g N_VDD_XI0/XI56/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI13/MM11 N_XI0/XI56/XI13/NET36_XI0/XI56/XI13/MM11_d
+ N_XI0/XI56/XI13/NET35_XI0/XI56/XI13/MM11_g N_VDD_XI0/XI56/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI14/MM2 N_XI0/XI56/XI14/NET34_XI0/XI56/XI14/MM2_d
+ N_XI0/XI56/XI14/NET33_XI0/XI56/XI14/MM2_g N_VSS_XI0/XI56/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM3 N_XI0/XI56/XI14/NET33_XI0/XI56/XI14/MM3_d
+ N_WL<108>_XI0/XI56/XI14/MM3_g N_BLN<1>_XI0/XI56/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM0 N_XI0/XI56/XI14/NET34_XI0/XI56/XI14/MM0_d
+ N_WL<108>_XI0/XI56/XI14/MM0_g N_BL<1>_XI0/XI56/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM1 N_XI0/XI56/XI14/NET33_XI0/XI56/XI14/MM1_d
+ N_XI0/XI56/XI14/NET34_XI0/XI56/XI14/MM1_g N_VSS_XI0/XI56/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM9 N_XI0/XI56/XI14/NET36_XI0/XI56/XI14/MM9_d
+ N_WL<109>_XI0/XI56/XI14/MM9_g N_BL<1>_XI0/XI56/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM6 N_XI0/XI56/XI14/NET35_XI0/XI56/XI14/MM6_d
+ N_XI0/XI56/XI14/NET36_XI0/XI56/XI14/MM6_g N_VSS_XI0/XI56/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM7 N_XI0/XI56/XI14/NET36_XI0/XI56/XI14/MM7_d
+ N_XI0/XI56/XI14/NET35_XI0/XI56/XI14/MM7_g N_VSS_XI0/XI56/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM8 N_XI0/XI56/XI14/NET35_XI0/XI56/XI14/MM8_d
+ N_WL<109>_XI0/XI56/XI14/MM8_g N_BLN<1>_XI0/XI56/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI14/MM5 N_XI0/XI56/XI14/NET34_XI0/XI56/XI14/MM5_d
+ N_XI0/XI56/XI14/NET33_XI0/XI56/XI14/MM5_g N_VDD_XI0/XI56/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI14/MM4 N_XI0/XI56/XI14/NET33_XI0/XI56/XI14/MM4_d
+ N_XI0/XI56/XI14/NET34_XI0/XI56/XI14/MM4_g N_VDD_XI0/XI56/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI14/MM10 N_XI0/XI56/XI14/NET35_XI0/XI56/XI14/MM10_d
+ N_XI0/XI56/XI14/NET36_XI0/XI56/XI14/MM10_g N_VDD_XI0/XI56/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI14/MM11 N_XI0/XI56/XI14/NET36_XI0/XI56/XI14/MM11_d
+ N_XI0/XI56/XI14/NET35_XI0/XI56/XI14/MM11_g N_VDD_XI0/XI56/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI15/MM2 N_XI0/XI56/XI15/NET34_XI0/XI56/XI15/MM2_d
+ N_XI0/XI56/XI15/NET33_XI0/XI56/XI15/MM2_g N_VSS_XI0/XI56/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM3 N_XI0/XI56/XI15/NET33_XI0/XI56/XI15/MM3_d
+ N_WL<108>_XI0/XI56/XI15/MM3_g N_BLN<0>_XI0/XI56/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM0 N_XI0/XI56/XI15/NET34_XI0/XI56/XI15/MM0_d
+ N_WL<108>_XI0/XI56/XI15/MM0_g N_BL<0>_XI0/XI56/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM1 N_XI0/XI56/XI15/NET33_XI0/XI56/XI15/MM1_d
+ N_XI0/XI56/XI15/NET34_XI0/XI56/XI15/MM1_g N_VSS_XI0/XI56/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM9 N_XI0/XI56/XI15/NET36_XI0/XI56/XI15/MM9_d
+ N_WL<109>_XI0/XI56/XI15/MM9_g N_BL<0>_XI0/XI56/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM6 N_XI0/XI56/XI15/NET35_XI0/XI56/XI15/MM6_d
+ N_XI0/XI56/XI15/NET36_XI0/XI56/XI15/MM6_g N_VSS_XI0/XI56/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM7 N_XI0/XI56/XI15/NET36_XI0/XI56/XI15/MM7_d
+ N_XI0/XI56/XI15/NET35_XI0/XI56/XI15/MM7_g N_VSS_XI0/XI56/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM8 N_XI0/XI56/XI15/NET35_XI0/XI56/XI15/MM8_d
+ N_WL<109>_XI0/XI56/XI15/MM8_g N_BLN<0>_XI0/XI56/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI56/XI15/MM5 N_XI0/XI56/XI15/NET34_XI0/XI56/XI15/MM5_d
+ N_XI0/XI56/XI15/NET33_XI0/XI56/XI15/MM5_g N_VDD_XI0/XI56/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI15/MM4 N_XI0/XI56/XI15/NET33_XI0/XI56/XI15/MM4_d
+ N_XI0/XI56/XI15/NET34_XI0/XI56/XI15/MM4_g N_VDD_XI0/XI56/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI15/MM10 N_XI0/XI56/XI15/NET35_XI0/XI56/XI15/MM10_d
+ N_XI0/XI56/XI15/NET36_XI0/XI56/XI15/MM10_g N_VDD_XI0/XI56/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI56/XI15/MM11 N_XI0/XI56/XI15/NET36_XI0/XI56/XI15/MM11_d
+ N_XI0/XI56/XI15/NET35_XI0/XI56/XI15/MM11_g N_VDD_XI0/XI56/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI0/MM2 N_XI0/XI57/XI0/NET34_XI0/XI57/XI0/MM2_d
+ N_XI0/XI57/XI0/NET33_XI0/XI57/XI0/MM2_g N_VSS_XI0/XI57/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM3 N_XI0/XI57/XI0/NET33_XI0/XI57/XI0/MM3_d
+ N_WL<110>_XI0/XI57/XI0/MM3_g N_BLN<15>_XI0/XI57/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM0 N_XI0/XI57/XI0/NET34_XI0/XI57/XI0/MM0_d
+ N_WL<110>_XI0/XI57/XI0/MM0_g N_BL<15>_XI0/XI57/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM1 N_XI0/XI57/XI0/NET33_XI0/XI57/XI0/MM1_d
+ N_XI0/XI57/XI0/NET34_XI0/XI57/XI0/MM1_g N_VSS_XI0/XI57/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM9 N_XI0/XI57/XI0/NET36_XI0/XI57/XI0/MM9_d
+ N_WL<111>_XI0/XI57/XI0/MM9_g N_BL<15>_XI0/XI57/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM6 N_XI0/XI57/XI0/NET35_XI0/XI57/XI0/MM6_d
+ N_XI0/XI57/XI0/NET36_XI0/XI57/XI0/MM6_g N_VSS_XI0/XI57/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM7 N_XI0/XI57/XI0/NET36_XI0/XI57/XI0/MM7_d
+ N_XI0/XI57/XI0/NET35_XI0/XI57/XI0/MM7_g N_VSS_XI0/XI57/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM8 N_XI0/XI57/XI0/NET35_XI0/XI57/XI0/MM8_d
+ N_WL<111>_XI0/XI57/XI0/MM8_g N_BLN<15>_XI0/XI57/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI0/MM5 N_XI0/XI57/XI0/NET34_XI0/XI57/XI0/MM5_d
+ N_XI0/XI57/XI0/NET33_XI0/XI57/XI0/MM5_g N_VDD_XI0/XI57/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI0/MM4 N_XI0/XI57/XI0/NET33_XI0/XI57/XI0/MM4_d
+ N_XI0/XI57/XI0/NET34_XI0/XI57/XI0/MM4_g N_VDD_XI0/XI57/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI0/MM10 N_XI0/XI57/XI0/NET35_XI0/XI57/XI0/MM10_d
+ N_XI0/XI57/XI0/NET36_XI0/XI57/XI0/MM10_g N_VDD_XI0/XI57/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI0/MM11 N_XI0/XI57/XI0/NET36_XI0/XI57/XI0/MM11_d
+ N_XI0/XI57/XI0/NET35_XI0/XI57/XI0/MM11_g N_VDD_XI0/XI57/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI1/MM2 N_XI0/XI57/XI1/NET34_XI0/XI57/XI1/MM2_d
+ N_XI0/XI57/XI1/NET33_XI0/XI57/XI1/MM2_g N_VSS_XI0/XI57/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM3 N_XI0/XI57/XI1/NET33_XI0/XI57/XI1/MM3_d
+ N_WL<110>_XI0/XI57/XI1/MM3_g N_BLN<14>_XI0/XI57/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM0 N_XI0/XI57/XI1/NET34_XI0/XI57/XI1/MM0_d
+ N_WL<110>_XI0/XI57/XI1/MM0_g N_BL<14>_XI0/XI57/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM1 N_XI0/XI57/XI1/NET33_XI0/XI57/XI1/MM1_d
+ N_XI0/XI57/XI1/NET34_XI0/XI57/XI1/MM1_g N_VSS_XI0/XI57/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM9 N_XI0/XI57/XI1/NET36_XI0/XI57/XI1/MM9_d
+ N_WL<111>_XI0/XI57/XI1/MM9_g N_BL<14>_XI0/XI57/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM6 N_XI0/XI57/XI1/NET35_XI0/XI57/XI1/MM6_d
+ N_XI0/XI57/XI1/NET36_XI0/XI57/XI1/MM6_g N_VSS_XI0/XI57/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM7 N_XI0/XI57/XI1/NET36_XI0/XI57/XI1/MM7_d
+ N_XI0/XI57/XI1/NET35_XI0/XI57/XI1/MM7_g N_VSS_XI0/XI57/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM8 N_XI0/XI57/XI1/NET35_XI0/XI57/XI1/MM8_d
+ N_WL<111>_XI0/XI57/XI1/MM8_g N_BLN<14>_XI0/XI57/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI1/MM5 N_XI0/XI57/XI1/NET34_XI0/XI57/XI1/MM5_d
+ N_XI0/XI57/XI1/NET33_XI0/XI57/XI1/MM5_g N_VDD_XI0/XI57/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI1/MM4 N_XI0/XI57/XI1/NET33_XI0/XI57/XI1/MM4_d
+ N_XI0/XI57/XI1/NET34_XI0/XI57/XI1/MM4_g N_VDD_XI0/XI57/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI1/MM10 N_XI0/XI57/XI1/NET35_XI0/XI57/XI1/MM10_d
+ N_XI0/XI57/XI1/NET36_XI0/XI57/XI1/MM10_g N_VDD_XI0/XI57/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI1/MM11 N_XI0/XI57/XI1/NET36_XI0/XI57/XI1/MM11_d
+ N_XI0/XI57/XI1/NET35_XI0/XI57/XI1/MM11_g N_VDD_XI0/XI57/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI2/MM2 N_XI0/XI57/XI2/NET34_XI0/XI57/XI2/MM2_d
+ N_XI0/XI57/XI2/NET33_XI0/XI57/XI2/MM2_g N_VSS_XI0/XI57/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM3 N_XI0/XI57/XI2/NET33_XI0/XI57/XI2/MM3_d
+ N_WL<110>_XI0/XI57/XI2/MM3_g N_BLN<13>_XI0/XI57/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM0 N_XI0/XI57/XI2/NET34_XI0/XI57/XI2/MM0_d
+ N_WL<110>_XI0/XI57/XI2/MM0_g N_BL<13>_XI0/XI57/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM1 N_XI0/XI57/XI2/NET33_XI0/XI57/XI2/MM1_d
+ N_XI0/XI57/XI2/NET34_XI0/XI57/XI2/MM1_g N_VSS_XI0/XI57/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM9 N_XI0/XI57/XI2/NET36_XI0/XI57/XI2/MM9_d
+ N_WL<111>_XI0/XI57/XI2/MM9_g N_BL<13>_XI0/XI57/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM6 N_XI0/XI57/XI2/NET35_XI0/XI57/XI2/MM6_d
+ N_XI0/XI57/XI2/NET36_XI0/XI57/XI2/MM6_g N_VSS_XI0/XI57/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM7 N_XI0/XI57/XI2/NET36_XI0/XI57/XI2/MM7_d
+ N_XI0/XI57/XI2/NET35_XI0/XI57/XI2/MM7_g N_VSS_XI0/XI57/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM8 N_XI0/XI57/XI2/NET35_XI0/XI57/XI2/MM8_d
+ N_WL<111>_XI0/XI57/XI2/MM8_g N_BLN<13>_XI0/XI57/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI2/MM5 N_XI0/XI57/XI2/NET34_XI0/XI57/XI2/MM5_d
+ N_XI0/XI57/XI2/NET33_XI0/XI57/XI2/MM5_g N_VDD_XI0/XI57/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI2/MM4 N_XI0/XI57/XI2/NET33_XI0/XI57/XI2/MM4_d
+ N_XI0/XI57/XI2/NET34_XI0/XI57/XI2/MM4_g N_VDD_XI0/XI57/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI2/MM10 N_XI0/XI57/XI2/NET35_XI0/XI57/XI2/MM10_d
+ N_XI0/XI57/XI2/NET36_XI0/XI57/XI2/MM10_g N_VDD_XI0/XI57/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI2/MM11 N_XI0/XI57/XI2/NET36_XI0/XI57/XI2/MM11_d
+ N_XI0/XI57/XI2/NET35_XI0/XI57/XI2/MM11_g N_VDD_XI0/XI57/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI3/MM2 N_XI0/XI57/XI3/NET34_XI0/XI57/XI3/MM2_d
+ N_XI0/XI57/XI3/NET33_XI0/XI57/XI3/MM2_g N_VSS_XI0/XI57/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM3 N_XI0/XI57/XI3/NET33_XI0/XI57/XI3/MM3_d
+ N_WL<110>_XI0/XI57/XI3/MM3_g N_BLN<12>_XI0/XI57/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM0 N_XI0/XI57/XI3/NET34_XI0/XI57/XI3/MM0_d
+ N_WL<110>_XI0/XI57/XI3/MM0_g N_BL<12>_XI0/XI57/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM1 N_XI0/XI57/XI3/NET33_XI0/XI57/XI3/MM1_d
+ N_XI0/XI57/XI3/NET34_XI0/XI57/XI3/MM1_g N_VSS_XI0/XI57/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM9 N_XI0/XI57/XI3/NET36_XI0/XI57/XI3/MM9_d
+ N_WL<111>_XI0/XI57/XI3/MM9_g N_BL<12>_XI0/XI57/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM6 N_XI0/XI57/XI3/NET35_XI0/XI57/XI3/MM6_d
+ N_XI0/XI57/XI3/NET36_XI0/XI57/XI3/MM6_g N_VSS_XI0/XI57/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM7 N_XI0/XI57/XI3/NET36_XI0/XI57/XI3/MM7_d
+ N_XI0/XI57/XI3/NET35_XI0/XI57/XI3/MM7_g N_VSS_XI0/XI57/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM8 N_XI0/XI57/XI3/NET35_XI0/XI57/XI3/MM8_d
+ N_WL<111>_XI0/XI57/XI3/MM8_g N_BLN<12>_XI0/XI57/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI3/MM5 N_XI0/XI57/XI3/NET34_XI0/XI57/XI3/MM5_d
+ N_XI0/XI57/XI3/NET33_XI0/XI57/XI3/MM5_g N_VDD_XI0/XI57/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI3/MM4 N_XI0/XI57/XI3/NET33_XI0/XI57/XI3/MM4_d
+ N_XI0/XI57/XI3/NET34_XI0/XI57/XI3/MM4_g N_VDD_XI0/XI57/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI3/MM10 N_XI0/XI57/XI3/NET35_XI0/XI57/XI3/MM10_d
+ N_XI0/XI57/XI3/NET36_XI0/XI57/XI3/MM10_g N_VDD_XI0/XI57/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI3/MM11 N_XI0/XI57/XI3/NET36_XI0/XI57/XI3/MM11_d
+ N_XI0/XI57/XI3/NET35_XI0/XI57/XI3/MM11_g N_VDD_XI0/XI57/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI4/MM2 N_XI0/XI57/XI4/NET34_XI0/XI57/XI4/MM2_d
+ N_XI0/XI57/XI4/NET33_XI0/XI57/XI4/MM2_g N_VSS_XI0/XI57/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM3 N_XI0/XI57/XI4/NET33_XI0/XI57/XI4/MM3_d
+ N_WL<110>_XI0/XI57/XI4/MM3_g N_BLN<11>_XI0/XI57/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM0 N_XI0/XI57/XI4/NET34_XI0/XI57/XI4/MM0_d
+ N_WL<110>_XI0/XI57/XI4/MM0_g N_BL<11>_XI0/XI57/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM1 N_XI0/XI57/XI4/NET33_XI0/XI57/XI4/MM1_d
+ N_XI0/XI57/XI4/NET34_XI0/XI57/XI4/MM1_g N_VSS_XI0/XI57/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM9 N_XI0/XI57/XI4/NET36_XI0/XI57/XI4/MM9_d
+ N_WL<111>_XI0/XI57/XI4/MM9_g N_BL<11>_XI0/XI57/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM6 N_XI0/XI57/XI4/NET35_XI0/XI57/XI4/MM6_d
+ N_XI0/XI57/XI4/NET36_XI0/XI57/XI4/MM6_g N_VSS_XI0/XI57/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM7 N_XI0/XI57/XI4/NET36_XI0/XI57/XI4/MM7_d
+ N_XI0/XI57/XI4/NET35_XI0/XI57/XI4/MM7_g N_VSS_XI0/XI57/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM8 N_XI0/XI57/XI4/NET35_XI0/XI57/XI4/MM8_d
+ N_WL<111>_XI0/XI57/XI4/MM8_g N_BLN<11>_XI0/XI57/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI4/MM5 N_XI0/XI57/XI4/NET34_XI0/XI57/XI4/MM5_d
+ N_XI0/XI57/XI4/NET33_XI0/XI57/XI4/MM5_g N_VDD_XI0/XI57/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI4/MM4 N_XI0/XI57/XI4/NET33_XI0/XI57/XI4/MM4_d
+ N_XI0/XI57/XI4/NET34_XI0/XI57/XI4/MM4_g N_VDD_XI0/XI57/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI4/MM10 N_XI0/XI57/XI4/NET35_XI0/XI57/XI4/MM10_d
+ N_XI0/XI57/XI4/NET36_XI0/XI57/XI4/MM10_g N_VDD_XI0/XI57/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI4/MM11 N_XI0/XI57/XI4/NET36_XI0/XI57/XI4/MM11_d
+ N_XI0/XI57/XI4/NET35_XI0/XI57/XI4/MM11_g N_VDD_XI0/XI57/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI5/MM2 N_XI0/XI57/XI5/NET34_XI0/XI57/XI5/MM2_d
+ N_XI0/XI57/XI5/NET33_XI0/XI57/XI5/MM2_g N_VSS_XI0/XI57/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM3 N_XI0/XI57/XI5/NET33_XI0/XI57/XI5/MM3_d
+ N_WL<110>_XI0/XI57/XI5/MM3_g N_BLN<10>_XI0/XI57/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM0 N_XI0/XI57/XI5/NET34_XI0/XI57/XI5/MM0_d
+ N_WL<110>_XI0/XI57/XI5/MM0_g N_BL<10>_XI0/XI57/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM1 N_XI0/XI57/XI5/NET33_XI0/XI57/XI5/MM1_d
+ N_XI0/XI57/XI5/NET34_XI0/XI57/XI5/MM1_g N_VSS_XI0/XI57/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM9 N_XI0/XI57/XI5/NET36_XI0/XI57/XI5/MM9_d
+ N_WL<111>_XI0/XI57/XI5/MM9_g N_BL<10>_XI0/XI57/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM6 N_XI0/XI57/XI5/NET35_XI0/XI57/XI5/MM6_d
+ N_XI0/XI57/XI5/NET36_XI0/XI57/XI5/MM6_g N_VSS_XI0/XI57/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM7 N_XI0/XI57/XI5/NET36_XI0/XI57/XI5/MM7_d
+ N_XI0/XI57/XI5/NET35_XI0/XI57/XI5/MM7_g N_VSS_XI0/XI57/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM8 N_XI0/XI57/XI5/NET35_XI0/XI57/XI5/MM8_d
+ N_WL<111>_XI0/XI57/XI5/MM8_g N_BLN<10>_XI0/XI57/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI5/MM5 N_XI0/XI57/XI5/NET34_XI0/XI57/XI5/MM5_d
+ N_XI0/XI57/XI5/NET33_XI0/XI57/XI5/MM5_g N_VDD_XI0/XI57/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI5/MM4 N_XI0/XI57/XI5/NET33_XI0/XI57/XI5/MM4_d
+ N_XI0/XI57/XI5/NET34_XI0/XI57/XI5/MM4_g N_VDD_XI0/XI57/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI5/MM10 N_XI0/XI57/XI5/NET35_XI0/XI57/XI5/MM10_d
+ N_XI0/XI57/XI5/NET36_XI0/XI57/XI5/MM10_g N_VDD_XI0/XI57/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI5/MM11 N_XI0/XI57/XI5/NET36_XI0/XI57/XI5/MM11_d
+ N_XI0/XI57/XI5/NET35_XI0/XI57/XI5/MM11_g N_VDD_XI0/XI57/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI6/MM2 N_XI0/XI57/XI6/NET34_XI0/XI57/XI6/MM2_d
+ N_XI0/XI57/XI6/NET33_XI0/XI57/XI6/MM2_g N_VSS_XI0/XI57/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM3 N_XI0/XI57/XI6/NET33_XI0/XI57/XI6/MM3_d
+ N_WL<110>_XI0/XI57/XI6/MM3_g N_BLN<9>_XI0/XI57/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM0 N_XI0/XI57/XI6/NET34_XI0/XI57/XI6/MM0_d
+ N_WL<110>_XI0/XI57/XI6/MM0_g N_BL<9>_XI0/XI57/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM1 N_XI0/XI57/XI6/NET33_XI0/XI57/XI6/MM1_d
+ N_XI0/XI57/XI6/NET34_XI0/XI57/XI6/MM1_g N_VSS_XI0/XI57/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM9 N_XI0/XI57/XI6/NET36_XI0/XI57/XI6/MM9_d
+ N_WL<111>_XI0/XI57/XI6/MM9_g N_BL<9>_XI0/XI57/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM6 N_XI0/XI57/XI6/NET35_XI0/XI57/XI6/MM6_d
+ N_XI0/XI57/XI6/NET36_XI0/XI57/XI6/MM6_g N_VSS_XI0/XI57/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM7 N_XI0/XI57/XI6/NET36_XI0/XI57/XI6/MM7_d
+ N_XI0/XI57/XI6/NET35_XI0/XI57/XI6/MM7_g N_VSS_XI0/XI57/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM8 N_XI0/XI57/XI6/NET35_XI0/XI57/XI6/MM8_d
+ N_WL<111>_XI0/XI57/XI6/MM8_g N_BLN<9>_XI0/XI57/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI6/MM5 N_XI0/XI57/XI6/NET34_XI0/XI57/XI6/MM5_d
+ N_XI0/XI57/XI6/NET33_XI0/XI57/XI6/MM5_g N_VDD_XI0/XI57/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI6/MM4 N_XI0/XI57/XI6/NET33_XI0/XI57/XI6/MM4_d
+ N_XI0/XI57/XI6/NET34_XI0/XI57/XI6/MM4_g N_VDD_XI0/XI57/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI6/MM10 N_XI0/XI57/XI6/NET35_XI0/XI57/XI6/MM10_d
+ N_XI0/XI57/XI6/NET36_XI0/XI57/XI6/MM10_g N_VDD_XI0/XI57/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI6/MM11 N_XI0/XI57/XI6/NET36_XI0/XI57/XI6/MM11_d
+ N_XI0/XI57/XI6/NET35_XI0/XI57/XI6/MM11_g N_VDD_XI0/XI57/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI7/MM2 N_XI0/XI57/XI7/NET34_XI0/XI57/XI7/MM2_d
+ N_XI0/XI57/XI7/NET33_XI0/XI57/XI7/MM2_g N_VSS_XI0/XI57/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM3 N_XI0/XI57/XI7/NET33_XI0/XI57/XI7/MM3_d
+ N_WL<110>_XI0/XI57/XI7/MM3_g N_BLN<8>_XI0/XI57/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM0 N_XI0/XI57/XI7/NET34_XI0/XI57/XI7/MM0_d
+ N_WL<110>_XI0/XI57/XI7/MM0_g N_BL<8>_XI0/XI57/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM1 N_XI0/XI57/XI7/NET33_XI0/XI57/XI7/MM1_d
+ N_XI0/XI57/XI7/NET34_XI0/XI57/XI7/MM1_g N_VSS_XI0/XI57/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM9 N_XI0/XI57/XI7/NET36_XI0/XI57/XI7/MM9_d
+ N_WL<111>_XI0/XI57/XI7/MM9_g N_BL<8>_XI0/XI57/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM6 N_XI0/XI57/XI7/NET35_XI0/XI57/XI7/MM6_d
+ N_XI0/XI57/XI7/NET36_XI0/XI57/XI7/MM6_g N_VSS_XI0/XI57/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM7 N_XI0/XI57/XI7/NET36_XI0/XI57/XI7/MM7_d
+ N_XI0/XI57/XI7/NET35_XI0/XI57/XI7/MM7_g N_VSS_XI0/XI57/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM8 N_XI0/XI57/XI7/NET35_XI0/XI57/XI7/MM8_d
+ N_WL<111>_XI0/XI57/XI7/MM8_g N_BLN<8>_XI0/XI57/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI7/MM5 N_XI0/XI57/XI7/NET34_XI0/XI57/XI7/MM5_d
+ N_XI0/XI57/XI7/NET33_XI0/XI57/XI7/MM5_g N_VDD_XI0/XI57/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI7/MM4 N_XI0/XI57/XI7/NET33_XI0/XI57/XI7/MM4_d
+ N_XI0/XI57/XI7/NET34_XI0/XI57/XI7/MM4_g N_VDD_XI0/XI57/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI7/MM10 N_XI0/XI57/XI7/NET35_XI0/XI57/XI7/MM10_d
+ N_XI0/XI57/XI7/NET36_XI0/XI57/XI7/MM10_g N_VDD_XI0/XI57/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI7/MM11 N_XI0/XI57/XI7/NET36_XI0/XI57/XI7/MM11_d
+ N_XI0/XI57/XI7/NET35_XI0/XI57/XI7/MM11_g N_VDD_XI0/XI57/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI8/MM2 N_XI0/XI57/XI8/NET34_XI0/XI57/XI8/MM2_d
+ N_XI0/XI57/XI8/NET33_XI0/XI57/XI8/MM2_g N_VSS_XI0/XI57/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM3 N_XI0/XI57/XI8/NET33_XI0/XI57/XI8/MM3_d
+ N_WL<110>_XI0/XI57/XI8/MM3_g N_BLN<7>_XI0/XI57/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM0 N_XI0/XI57/XI8/NET34_XI0/XI57/XI8/MM0_d
+ N_WL<110>_XI0/XI57/XI8/MM0_g N_BL<7>_XI0/XI57/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM1 N_XI0/XI57/XI8/NET33_XI0/XI57/XI8/MM1_d
+ N_XI0/XI57/XI8/NET34_XI0/XI57/XI8/MM1_g N_VSS_XI0/XI57/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM9 N_XI0/XI57/XI8/NET36_XI0/XI57/XI8/MM9_d
+ N_WL<111>_XI0/XI57/XI8/MM9_g N_BL<7>_XI0/XI57/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM6 N_XI0/XI57/XI8/NET35_XI0/XI57/XI8/MM6_d
+ N_XI0/XI57/XI8/NET36_XI0/XI57/XI8/MM6_g N_VSS_XI0/XI57/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM7 N_XI0/XI57/XI8/NET36_XI0/XI57/XI8/MM7_d
+ N_XI0/XI57/XI8/NET35_XI0/XI57/XI8/MM7_g N_VSS_XI0/XI57/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM8 N_XI0/XI57/XI8/NET35_XI0/XI57/XI8/MM8_d
+ N_WL<111>_XI0/XI57/XI8/MM8_g N_BLN<7>_XI0/XI57/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI8/MM5 N_XI0/XI57/XI8/NET34_XI0/XI57/XI8/MM5_d
+ N_XI0/XI57/XI8/NET33_XI0/XI57/XI8/MM5_g N_VDD_XI0/XI57/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI8/MM4 N_XI0/XI57/XI8/NET33_XI0/XI57/XI8/MM4_d
+ N_XI0/XI57/XI8/NET34_XI0/XI57/XI8/MM4_g N_VDD_XI0/XI57/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI8/MM10 N_XI0/XI57/XI8/NET35_XI0/XI57/XI8/MM10_d
+ N_XI0/XI57/XI8/NET36_XI0/XI57/XI8/MM10_g N_VDD_XI0/XI57/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI8/MM11 N_XI0/XI57/XI8/NET36_XI0/XI57/XI8/MM11_d
+ N_XI0/XI57/XI8/NET35_XI0/XI57/XI8/MM11_g N_VDD_XI0/XI57/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI9/MM2 N_XI0/XI57/XI9/NET34_XI0/XI57/XI9/MM2_d
+ N_XI0/XI57/XI9/NET33_XI0/XI57/XI9/MM2_g N_VSS_XI0/XI57/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM3 N_XI0/XI57/XI9/NET33_XI0/XI57/XI9/MM3_d
+ N_WL<110>_XI0/XI57/XI9/MM3_g N_BLN<6>_XI0/XI57/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM0 N_XI0/XI57/XI9/NET34_XI0/XI57/XI9/MM0_d
+ N_WL<110>_XI0/XI57/XI9/MM0_g N_BL<6>_XI0/XI57/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM1 N_XI0/XI57/XI9/NET33_XI0/XI57/XI9/MM1_d
+ N_XI0/XI57/XI9/NET34_XI0/XI57/XI9/MM1_g N_VSS_XI0/XI57/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM9 N_XI0/XI57/XI9/NET36_XI0/XI57/XI9/MM9_d
+ N_WL<111>_XI0/XI57/XI9/MM9_g N_BL<6>_XI0/XI57/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM6 N_XI0/XI57/XI9/NET35_XI0/XI57/XI9/MM6_d
+ N_XI0/XI57/XI9/NET36_XI0/XI57/XI9/MM6_g N_VSS_XI0/XI57/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM7 N_XI0/XI57/XI9/NET36_XI0/XI57/XI9/MM7_d
+ N_XI0/XI57/XI9/NET35_XI0/XI57/XI9/MM7_g N_VSS_XI0/XI57/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM8 N_XI0/XI57/XI9/NET35_XI0/XI57/XI9/MM8_d
+ N_WL<111>_XI0/XI57/XI9/MM8_g N_BLN<6>_XI0/XI57/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI9/MM5 N_XI0/XI57/XI9/NET34_XI0/XI57/XI9/MM5_d
+ N_XI0/XI57/XI9/NET33_XI0/XI57/XI9/MM5_g N_VDD_XI0/XI57/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI9/MM4 N_XI0/XI57/XI9/NET33_XI0/XI57/XI9/MM4_d
+ N_XI0/XI57/XI9/NET34_XI0/XI57/XI9/MM4_g N_VDD_XI0/XI57/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI9/MM10 N_XI0/XI57/XI9/NET35_XI0/XI57/XI9/MM10_d
+ N_XI0/XI57/XI9/NET36_XI0/XI57/XI9/MM10_g N_VDD_XI0/XI57/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI9/MM11 N_XI0/XI57/XI9/NET36_XI0/XI57/XI9/MM11_d
+ N_XI0/XI57/XI9/NET35_XI0/XI57/XI9/MM11_g N_VDD_XI0/XI57/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI10/MM2 N_XI0/XI57/XI10/NET34_XI0/XI57/XI10/MM2_d
+ N_XI0/XI57/XI10/NET33_XI0/XI57/XI10/MM2_g N_VSS_XI0/XI57/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM3 N_XI0/XI57/XI10/NET33_XI0/XI57/XI10/MM3_d
+ N_WL<110>_XI0/XI57/XI10/MM3_g N_BLN<5>_XI0/XI57/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM0 N_XI0/XI57/XI10/NET34_XI0/XI57/XI10/MM0_d
+ N_WL<110>_XI0/XI57/XI10/MM0_g N_BL<5>_XI0/XI57/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM1 N_XI0/XI57/XI10/NET33_XI0/XI57/XI10/MM1_d
+ N_XI0/XI57/XI10/NET34_XI0/XI57/XI10/MM1_g N_VSS_XI0/XI57/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM9 N_XI0/XI57/XI10/NET36_XI0/XI57/XI10/MM9_d
+ N_WL<111>_XI0/XI57/XI10/MM9_g N_BL<5>_XI0/XI57/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM6 N_XI0/XI57/XI10/NET35_XI0/XI57/XI10/MM6_d
+ N_XI0/XI57/XI10/NET36_XI0/XI57/XI10/MM6_g N_VSS_XI0/XI57/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM7 N_XI0/XI57/XI10/NET36_XI0/XI57/XI10/MM7_d
+ N_XI0/XI57/XI10/NET35_XI0/XI57/XI10/MM7_g N_VSS_XI0/XI57/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM8 N_XI0/XI57/XI10/NET35_XI0/XI57/XI10/MM8_d
+ N_WL<111>_XI0/XI57/XI10/MM8_g N_BLN<5>_XI0/XI57/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI10/MM5 N_XI0/XI57/XI10/NET34_XI0/XI57/XI10/MM5_d
+ N_XI0/XI57/XI10/NET33_XI0/XI57/XI10/MM5_g N_VDD_XI0/XI57/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI10/MM4 N_XI0/XI57/XI10/NET33_XI0/XI57/XI10/MM4_d
+ N_XI0/XI57/XI10/NET34_XI0/XI57/XI10/MM4_g N_VDD_XI0/XI57/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI10/MM10 N_XI0/XI57/XI10/NET35_XI0/XI57/XI10/MM10_d
+ N_XI0/XI57/XI10/NET36_XI0/XI57/XI10/MM10_g N_VDD_XI0/XI57/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI10/MM11 N_XI0/XI57/XI10/NET36_XI0/XI57/XI10/MM11_d
+ N_XI0/XI57/XI10/NET35_XI0/XI57/XI10/MM11_g N_VDD_XI0/XI57/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI11/MM2 N_XI0/XI57/XI11/NET34_XI0/XI57/XI11/MM2_d
+ N_XI0/XI57/XI11/NET33_XI0/XI57/XI11/MM2_g N_VSS_XI0/XI57/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM3 N_XI0/XI57/XI11/NET33_XI0/XI57/XI11/MM3_d
+ N_WL<110>_XI0/XI57/XI11/MM3_g N_BLN<4>_XI0/XI57/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM0 N_XI0/XI57/XI11/NET34_XI0/XI57/XI11/MM0_d
+ N_WL<110>_XI0/XI57/XI11/MM0_g N_BL<4>_XI0/XI57/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM1 N_XI0/XI57/XI11/NET33_XI0/XI57/XI11/MM1_d
+ N_XI0/XI57/XI11/NET34_XI0/XI57/XI11/MM1_g N_VSS_XI0/XI57/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM9 N_XI0/XI57/XI11/NET36_XI0/XI57/XI11/MM9_d
+ N_WL<111>_XI0/XI57/XI11/MM9_g N_BL<4>_XI0/XI57/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM6 N_XI0/XI57/XI11/NET35_XI0/XI57/XI11/MM6_d
+ N_XI0/XI57/XI11/NET36_XI0/XI57/XI11/MM6_g N_VSS_XI0/XI57/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM7 N_XI0/XI57/XI11/NET36_XI0/XI57/XI11/MM7_d
+ N_XI0/XI57/XI11/NET35_XI0/XI57/XI11/MM7_g N_VSS_XI0/XI57/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM8 N_XI0/XI57/XI11/NET35_XI0/XI57/XI11/MM8_d
+ N_WL<111>_XI0/XI57/XI11/MM8_g N_BLN<4>_XI0/XI57/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI11/MM5 N_XI0/XI57/XI11/NET34_XI0/XI57/XI11/MM5_d
+ N_XI0/XI57/XI11/NET33_XI0/XI57/XI11/MM5_g N_VDD_XI0/XI57/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI11/MM4 N_XI0/XI57/XI11/NET33_XI0/XI57/XI11/MM4_d
+ N_XI0/XI57/XI11/NET34_XI0/XI57/XI11/MM4_g N_VDD_XI0/XI57/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI11/MM10 N_XI0/XI57/XI11/NET35_XI0/XI57/XI11/MM10_d
+ N_XI0/XI57/XI11/NET36_XI0/XI57/XI11/MM10_g N_VDD_XI0/XI57/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI11/MM11 N_XI0/XI57/XI11/NET36_XI0/XI57/XI11/MM11_d
+ N_XI0/XI57/XI11/NET35_XI0/XI57/XI11/MM11_g N_VDD_XI0/XI57/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI12/MM2 N_XI0/XI57/XI12/NET34_XI0/XI57/XI12/MM2_d
+ N_XI0/XI57/XI12/NET33_XI0/XI57/XI12/MM2_g N_VSS_XI0/XI57/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM3 N_XI0/XI57/XI12/NET33_XI0/XI57/XI12/MM3_d
+ N_WL<110>_XI0/XI57/XI12/MM3_g N_BLN<3>_XI0/XI57/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM0 N_XI0/XI57/XI12/NET34_XI0/XI57/XI12/MM0_d
+ N_WL<110>_XI0/XI57/XI12/MM0_g N_BL<3>_XI0/XI57/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM1 N_XI0/XI57/XI12/NET33_XI0/XI57/XI12/MM1_d
+ N_XI0/XI57/XI12/NET34_XI0/XI57/XI12/MM1_g N_VSS_XI0/XI57/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM9 N_XI0/XI57/XI12/NET36_XI0/XI57/XI12/MM9_d
+ N_WL<111>_XI0/XI57/XI12/MM9_g N_BL<3>_XI0/XI57/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM6 N_XI0/XI57/XI12/NET35_XI0/XI57/XI12/MM6_d
+ N_XI0/XI57/XI12/NET36_XI0/XI57/XI12/MM6_g N_VSS_XI0/XI57/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM7 N_XI0/XI57/XI12/NET36_XI0/XI57/XI12/MM7_d
+ N_XI0/XI57/XI12/NET35_XI0/XI57/XI12/MM7_g N_VSS_XI0/XI57/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM8 N_XI0/XI57/XI12/NET35_XI0/XI57/XI12/MM8_d
+ N_WL<111>_XI0/XI57/XI12/MM8_g N_BLN<3>_XI0/XI57/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI12/MM5 N_XI0/XI57/XI12/NET34_XI0/XI57/XI12/MM5_d
+ N_XI0/XI57/XI12/NET33_XI0/XI57/XI12/MM5_g N_VDD_XI0/XI57/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI12/MM4 N_XI0/XI57/XI12/NET33_XI0/XI57/XI12/MM4_d
+ N_XI0/XI57/XI12/NET34_XI0/XI57/XI12/MM4_g N_VDD_XI0/XI57/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI12/MM10 N_XI0/XI57/XI12/NET35_XI0/XI57/XI12/MM10_d
+ N_XI0/XI57/XI12/NET36_XI0/XI57/XI12/MM10_g N_VDD_XI0/XI57/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI12/MM11 N_XI0/XI57/XI12/NET36_XI0/XI57/XI12/MM11_d
+ N_XI0/XI57/XI12/NET35_XI0/XI57/XI12/MM11_g N_VDD_XI0/XI57/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI13/MM2 N_XI0/XI57/XI13/NET34_XI0/XI57/XI13/MM2_d
+ N_XI0/XI57/XI13/NET33_XI0/XI57/XI13/MM2_g N_VSS_XI0/XI57/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM3 N_XI0/XI57/XI13/NET33_XI0/XI57/XI13/MM3_d
+ N_WL<110>_XI0/XI57/XI13/MM3_g N_BLN<2>_XI0/XI57/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM0 N_XI0/XI57/XI13/NET34_XI0/XI57/XI13/MM0_d
+ N_WL<110>_XI0/XI57/XI13/MM0_g N_BL<2>_XI0/XI57/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM1 N_XI0/XI57/XI13/NET33_XI0/XI57/XI13/MM1_d
+ N_XI0/XI57/XI13/NET34_XI0/XI57/XI13/MM1_g N_VSS_XI0/XI57/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM9 N_XI0/XI57/XI13/NET36_XI0/XI57/XI13/MM9_d
+ N_WL<111>_XI0/XI57/XI13/MM9_g N_BL<2>_XI0/XI57/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM6 N_XI0/XI57/XI13/NET35_XI0/XI57/XI13/MM6_d
+ N_XI0/XI57/XI13/NET36_XI0/XI57/XI13/MM6_g N_VSS_XI0/XI57/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM7 N_XI0/XI57/XI13/NET36_XI0/XI57/XI13/MM7_d
+ N_XI0/XI57/XI13/NET35_XI0/XI57/XI13/MM7_g N_VSS_XI0/XI57/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM8 N_XI0/XI57/XI13/NET35_XI0/XI57/XI13/MM8_d
+ N_WL<111>_XI0/XI57/XI13/MM8_g N_BLN<2>_XI0/XI57/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI13/MM5 N_XI0/XI57/XI13/NET34_XI0/XI57/XI13/MM5_d
+ N_XI0/XI57/XI13/NET33_XI0/XI57/XI13/MM5_g N_VDD_XI0/XI57/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI13/MM4 N_XI0/XI57/XI13/NET33_XI0/XI57/XI13/MM4_d
+ N_XI0/XI57/XI13/NET34_XI0/XI57/XI13/MM4_g N_VDD_XI0/XI57/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI13/MM10 N_XI0/XI57/XI13/NET35_XI0/XI57/XI13/MM10_d
+ N_XI0/XI57/XI13/NET36_XI0/XI57/XI13/MM10_g N_VDD_XI0/XI57/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI13/MM11 N_XI0/XI57/XI13/NET36_XI0/XI57/XI13/MM11_d
+ N_XI0/XI57/XI13/NET35_XI0/XI57/XI13/MM11_g N_VDD_XI0/XI57/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI14/MM2 N_XI0/XI57/XI14/NET34_XI0/XI57/XI14/MM2_d
+ N_XI0/XI57/XI14/NET33_XI0/XI57/XI14/MM2_g N_VSS_XI0/XI57/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM3 N_XI0/XI57/XI14/NET33_XI0/XI57/XI14/MM3_d
+ N_WL<110>_XI0/XI57/XI14/MM3_g N_BLN<1>_XI0/XI57/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM0 N_XI0/XI57/XI14/NET34_XI0/XI57/XI14/MM0_d
+ N_WL<110>_XI0/XI57/XI14/MM0_g N_BL<1>_XI0/XI57/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM1 N_XI0/XI57/XI14/NET33_XI0/XI57/XI14/MM1_d
+ N_XI0/XI57/XI14/NET34_XI0/XI57/XI14/MM1_g N_VSS_XI0/XI57/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM9 N_XI0/XI57/XI14/NET36_XI0/XI57/XI14/MM9_d
+ N_WL<111>_XI0/XI57/XI14/MM9_g N_BL<1>_XI0/XI57/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM6 N_XI0/XI57/XI14/NET35_XI0/XI57/XI14/MM6_d
+ N_XI0/XI57/XI14/NET36_XI0/XI57/XI14/MM6_g N_VSS_XI0/XI57/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM7 N_XI0/XI57/XI14/NET36_XI0/XI57/XI14/MM7_d
+ N_XI0/XI57/XI14/NET35_XI0/XI57/XI14/MM7_g N_VSS_XI0/XI57/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM8 N_XI0/XI57/XI14/NET35_XI0/XI57/XI14/MM8_d
+ N_WL<111>_XI0/XI57/XI14/MM8_g N_BLN<1>_XI0/XI57/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI14/MM5 N_XI0/XI57/XI14/NET34_XI0/XI57/XI14/MM5_d
+ N_XI0/XI57/XI14/NET33_XI0/XI57/XI14/MM5_g N_VDD_XI0/XI57/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI14/MM4 N_XI0/XI57/XI14/NET33_XI0/XI57/XI14/MM4_d
+ N_XI0/XI57/XI14/NET34_XI0/XI57/XI14/MM4_g N_VDD_XI0/XI57/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI14/MM10 N_XI0/XI57/XI14/NET35_XI0/XI57/XI14/MM10_d
+ N_XI0/XI57/XI14/NET36_XI0/XI57/XI14/MM10_g N_VDD_XI0/XI57/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI14/MM11 N_XI0/XI57/XI14/NET36_XI0/XI57/XI14/MM11_d
+ N_XI0/XI57/XI14/NET35_XI0/XI57/XI14/MM11_g N_VDD_XI0/XI57/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI15/MM2 N_XI0/XI57/XI15/NET34_XI0/XI57/XI15/MM2_d
+ N_XI0/XI57/XI15/NET33_XI0/XI57/XI15/MM2_g N_VSS_XI0/XI57/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM3 N_XI0/XI57/XI15/NET33_XI0/XI57/XI15/MM3_d
+ N_WL<110>_XI0/XI57/XI15/MM3_g N_BLN<0>_XI0/XI57/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM0 N_XI0/XI57/XI15/NET34_XI0/XI57/XI15/MM0_d
+ N_WL<110>_XI0/XI57/XI15/MM0_g N_BL<0>_XI0/XI57/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM1 N_XI0/XI57/XI15/NET33_XI0/XI57/XI15/MM1_d
+ N_XI0/XI57/XI15/NET34_XI0/XI57/XI15/MM1_g N_VSS_XI0/XI57/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM9 N_XI0/XI57/XI15/NET36_XI0/XI57/XI15/MM9_d
+ N_WL<111>_XI0/XI57/XI15/MM9_g N_BL<0>_XI0/XI57/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM6 N_XI0/XI57/XI15/NET35_XI0/XI57/XI15/MM6_d
+ N_XI0/XI57/XI15/NET36_XI0/XI57/XI15/MM6_g N_VSS_XI0/XI57/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM7 N_XI0/XI57/XI15/NET36_XI0/XI57/XI15/MM7_d
+ N_XI0/XI57/XI15/NET35_XI0/XI57/XI15/MM7_g N_VSS_XI0/XI57/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM8 N_XI0/XI57/XI15/NET35_XI0/XI57/XI15/MM8_d
+ N_WL<111>_XI0/XI57/XI15/MM8_g N_BLN<0>_XI0/XI57/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI57/XI15/MM5 N_XI0/XI57/XI15/NET34_XI0/XI57/XI15/MM5_d
+ N_XI0/XI57/XI15/NET33_XI0/XI57/XI15/MM5_g N_VDD_XI0/XI57/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI15/MM4 N_XI0/XI57/XI15/NET33_XI0/XI57/XI15/MM4_d
+ N_XI0/XI57/XI15/NET34_XI0/XI57/XI15/MM4_g N_VDD_XI0/XI57/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI15/MM10 N_XI0/XI57/XI15/NET35_XI0/XI57/XI15/MM10_d
+ N_XI0/XI57/XI15/NET36_XI0/XI57/XI15/MM10_g N_VDD_XI0/XI57/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI57/XI15/MM11 N_XI0/XI57/XI15/NET36_XI0/XI57/XI15/MM11_d
+ N_XI0/XI57/XI15/NET35_XI0/XI57/XI15/MM11_g N_VDD_XI0/XI57/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI0/MM2 N_XI0/XI58/XI0/NET34_XI0/XI58/XI0/MM2_d
+ N_XI0/XI58/XI0/NET33_XI0/XI58/XI0/MM2_g N_VSS_XI0/XI58/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM3 N_XI0/XI58/XI0/NET33_XI0/XI58/XI0/MM3_d
+ N_WL<112>_XI0/XI58/XI0/MM3_g N_BLN<15>_XI0/XI58/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM0 N_XI0/XI58/XI0/NET34_XI0/XI58/XI0/MM0_d
+ N_WL<112>_XI0/XI58/XI0/MM0_g N_BL<15>_XI0/XI58/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM1 N_XI0/XI58/XI0/NET33_XI0/XI58/XI0/MM1_d
+ N_XI0/XI58/XI0/NET34_XI0/XI58/XI0/MM1_g N_VSS_XI0/XI58/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM9 N_XI0/XI58/XI0/NET36_XI0/XI58/XI0/MM9_d
+ N_WL<113>_XI0/XI58/XI0/MM9_g N_BL<15>_XI0/XI58/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM6 N_XI0/XI58/XI0/NET35_XI0/XI58/XI0/MM6_d
+ N_XI0/XI58/XI0/NET36_XI0/XI58/XI0/MM6_g N_VSS_XI0/XI58/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM7 N_XI0/XI58/XI0/NET36_XI0/XI58/XI0/MM7_d
+ N_XI0/XI58/XI0/NET35_XI0/XI58/XI0/MM7_g N_VSS_XI0/XI58/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM8 N_XI0/XI58/XI0/NET35_XI0/XI58/XI0/MM8_d
+ N_WL<113>_XI0/XI58/XI0/MM8_g N_BLN<15>_XI0/XI58/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI0/MM5 N_XI0/XI58/XI0/NET34_XI0/XI58/XI0/MM5_d
+ N_XI0/XI58/XI0/NET33_XI0/XI58/XI0/MM5_g N_VDD_XI0/XI58/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI0/MM4 N_XI0/XI58/XI0/NET33_XI0/XI58/XI0/MM4_d
+ N_XI0/XI58/XI0/NET34_XI0/XI58/XI0/MM4_g N_VDD_XI0/XI58/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI0/MM10 N_XI0/XI58/XI0/NET35_XI0/XI58/XI0/MM10_d
+ N_XI0/XI58/XI0/NET36_XI0/XI58/XI0/MM10_g N_VDD_XI0/XI58/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI0/MM11 N_XI0/XI58/XI0/NET36_XI0/XI58/XI0/MM11_d
+ N_XI0/XI58/XI0/NET35_XI0/XI58/XI0/MM11_g N_VDD_XI0/XI58/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI1/MM2 N_XI0/XI58/XI1/NET34_XI0/XI58/XI1/MM2_d
+ N_XI0/XI58/XI1/NET33_XI0/XI58/XI1/MM2_g N_VSS_XI0/XI58/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM3 N_XI0/XI58/XI1/NET33_XI0/XI58/XI1/MM3_d
+ N_WL<112>_XI0/XI58/XI1/MM3_g N_BLN<14>_XI0/XI58/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM0 N_XI0/XI58/XI1/NET34_XI0/XI58/XI1/MM0_d
+ N_WL<112>_XI0/XI58/XI1/MM0_g N_BL<14>_XI0/XI58/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM1 N_XI0/XI58/XI1/NET33_XI0/XI58/XI1/MM1_d
+ N_XI0/XI58/XI1/NET34_XI0/XI58/XI1/MM1_g N_VSS_XI0/XI58/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM9 N_XI0/XI58/XI1/NET36_XI0/XI58/XI1/MM9_d
+ N_WL<113>_XI0/XI58/XI1/MM9_g N_BL<14>_XI0/XI58/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM6 N_XI0/XI58/XI1/NET35_XI0/XI58/XI1/MM6_d
+ N_XI0/XI58/XI1/NET36_XI0/XI58/XI1/MM6_g N_VSS_XI0/XI58/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM7 N_XI0/XI58/XI1/NET36_XI0/XI58/XI1/MM7_d
+ N_XI0/XI58/XI1/NET35_XI0/XI58/XI1/MM7_g N_VSS_XI0/XI58/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM8 N_XI0/XI58/XI1/NET35_XI0/XI58/XI1/MM8_d
+ N_WL<113>_XI0/XI58/XI1/MM8_g N_BLN<14>_XI0/XI58/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI1/MM5 N_XI0/XI58/XI1/NET34_XI0/XI58/XI1/MM5_d
+ N_XI0/XI58/XI1/NET33_XI0/XI58/XI1/MM5_g N_VDD_XI0/XI58/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI1/MM4 N_XI0/XI58/XI1/NET33_XI0/XI58/XI1/MM4_d
+ N_XI0/XI58/XI1/NET34_XI0/XI58/XI1/MM4_g N_VDD_XI0/XI58/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI1/MM10 N_XI0/XI58/XI1/NET35_XI0/XI58/XI1/MM10_d
+ N_XI0/XI58/XI1/NET36_XI0/XI58/XI1/MM10_g N_VDD_XI0/XI58/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI1/MM11 N_XI0/XI58/XI1/NET36_XI0/XI58/XI1/MM11_d
+ N_XI0/XI58/XI1/NET35_XI0/XI58/XI1/MM11_g N_VDD_XI0/XI58/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI2/MM2 N_XI0/XI58/XI2/NET34_XI0/XI58/XI2/MM2_d
+ N_XI0/XI58/XI2/NET33_XI0/XI58/XI2/MM2_g N_VSS_XI0/XI58/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM3 N_XI0/XI58/XI2/NET33_XI0/XI58/XI2/MM3_d
+ N_WL<112>_XI0/XI58/XI2/MM3_g N_BLN<13>_XI0/XI58/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM0 N_XI0/XI58/XI2/NET34_XI0/XI58/XI2/MM0_d
+ N_WL<112>_XI0/XI58/XI2/MM0_g N_BL<13>_XI0/XI58/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM1 N_XI0/XI58/XI2/NET33_XI0/XI58/XI2/MM1_d
+ N_XI0/XI58/XI2/NET34_XI0/XI58/XI2/MM1_g N_VSS_XI0/XI58/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM9 N_XI0/XI58/XI2/NET36_XI0/XI58/XI2/MM9_d
+ N_WL<113>_XI0/XI58/XI2/MM9_g N_BL<13>_XI0/XI58/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM6 N_XI0/XI58/XI2/NET35_XI0/XI58/XI2/MM6_d
+ N_XI0/XI58/XI2/NET36_XI0/XI58/XI2/MM6_g N_VSS_XI0/XI58/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM7 N_XI0/XI58/XI2/NET36_XI0/XI58/XI2/MM7_d
+ N_XI0/XI58/XI2/NET35_XI0/XI58/XI2/MM7_g N_VSS_XI0/XI58/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM8 N_XI0/XI58/XI2/NET35_XI0/XI58/XI2/MM8_d
+ N_WL<113>_XI0/XI58/XI2/MM8_g N_BLN<13>_XI0/XI58/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI2/MM5 N_XI0/XI58/XI2/NET34_XI0/XI58/XI2/MM5_d
+ N_XI0/XI58/XI2/NET33_XI0/XI58/XI2/MM5_g N_VDD_XI0/XI58/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI2/MM4 N_XI0/XI58/XI2/NET33_XI0/XI58/XI2/MM4_d
+ N_XI0/XI58/XI2/NET34_XI0/XI58/XI2/MM4_g N_VDD_XI0/XI58/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI2/MM10 N_XI0/XI58/XI2/NET35_XI0/XI58/XI2/MM10_d
+ N_XI0/XI58/XI2/NET36_XI0/XI58/XI2/MM10_g N_VDD_XI0/XI58/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI2/MM11 N_XI0/XI58/XI2/NET36_XI0/XI58/XI2/MM11_d
+ N_XI0/XI58/XI2/NET35_XI0/XI58/XI2/MM11_g N_VDD_XI0/XI58/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI3/MM2 N_XI0/XI58/XI3/NET34_XI0/XI58/XI3/MM2_d
+ N_XI0/XI58/XI3/NET33_XI0/XI58/XI3/MM2_g N_VSS_XI0/XI58/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM3 N_XI0/XI58/XI3/NET33_XI0/XI58/XI3/MM3_d
+ N_WL<112>_XI0/XI58/XI3/MM3_g N_BLN<12>_XI0/XI58/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM0 N_XI0/XI58/XI3/NET34_XI0/XI58/XI3/MM0_d
+ N_WL<112>_XI0/XI58/XI3/MM0_g N_BL<12>_XI0/XI58/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM1 N_XI0/XI58/XI3/NET33_XI0/XI58/XI3/MM1_d
+ N_XI0/XI58/XI3/NET34_XI0/XI58/XI3/MM1_g N_VSS_XI0/XI58/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM9 N_XI0/XI58/XI3/NET36_XI0/XI58/XI3/MM9_d
+ N_WL<113>_XI0/XI58/XI3/MM9_g N_BL<12>_XI0/XI58/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM6 N_XI0/XI58/XI3/NET35_XI0/XI58/XI3/MM6_d
+ N_XI0/XI58/XI3/NET36_XI0/XI58/XI3/MM6_g N_VSS_XI0/XI58/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM7 N_XI0/XI58/XI3/NET36_XI0/XI58/XI3/MM7_d
+ N_XI0/XI58/XI3/NET35_XI0/XI58/XI3/MM7_g N_VSS_XI0/XI58/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM8 N_XI0/XI58/XI3/NET35_XI0/XI58/XI3/MM8_d
+ N_WL<113>_XI0/XI58/XI3/MM8_g N_BLN<12>_XI0/XI58/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI3/MM5 N_XI0/XI58/XI3/NET34_XI0/XI58/XI3/MM5_d
+ N_XI0/XI58/XI3/NET33_XI0/XI58/XI3/MM5_g N_VDD_XI0/XI58/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI3/MM4 N_XI0/XI58/XI3/NET33_XI0/XI58/XI3/MM4_d
+ N_XI0/XI58/XI3/NET34_XI0/XI58/XI3/MM4_g N_VDD_XI0/XI58/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI3/MM10 N_XI0/XI58/XI3/NET35_XI0/XI58/XI3/MM10_d
+ N_XI0/XI58/XI3/NET36_XI0/XI58/XI3/MM10_g N_VDD_XI0/XI58/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI3/MM11 N_XI0/XI58/XI3/NET36_XI0/XI58/XI3/MM11_d
+ N_XI0/XI58/XI3/NET35_XI0/XI58/XI3/MM11_g N_VDD_XI0/XI58/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI4/MM2 N_XI0/XI58/XI4/NET34_XI0/XI58/XI4/MM2_d
+ N_XI0/XI58/XI4/NET33_XI0/XI58/XI4/MM2_g N_VSS_XI0/XI58/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM3 N_XI0/XI58/XI4/NET33_XI0/XI58/XI4/MM3_d
+ N_WL<112>_XI0/XI58/XI4/MM3_g N_BLN<11>_XI0/XI58/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM0 N_XI0/XI58/XI4/NET34_XI0/XI58/XI4/MM0_d
+ N_WL<112>_XI0/XI58/XI4/MM0_g N_BL<11>_XI0/XI58/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM1 N_XI0/XI58/XI4/NET33_XI0/XI58/XI4/MM1_d
+ N_XI0/XI58/XI4/NET34_XI0/XI58/XI4/MM1_g N_VSS_XI0/XI58/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM9 N_XI0/XI58/XI4/NET36_XI0/XI58/XI4/MM9_d
+ N_WL<113>_XI0/XI58/XI4/MM9_g N_BL<11>_XI0/XI58/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM6 N_XI0/XI58/XI4/NET35_XI0/XI58/XI4/MM6_d
+ N_XI0/XI58/XI4/NET36_XI0/XI58/XI4/MM6_g N_VSS_XI0/XI58/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM7 N_XI0/XI58/XI4/NET36_XI0/XI58/XI4/MM7_d
+ N_XI0/XI58/XI4/NET35_XI0/XI58/XI4/MM7_g N_VSS_XI0/XI58/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM8 N_XI0/XI58/XI4/NET35_XI0/XI58/XI4/MM8_d
+ N_WL<113>_XI0/XI58/XI4/MM8_g N_BLN<11>_XI0/XI58/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI4/MM5 N_XI0/XI58/XI4/NET34_XI0/XI58/XI4/MM5_d
+ N_XI0/XI58/XI4/NET33_XI0/XI58/XI4/MM5_g N_VDD_XI0/XI58/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI4/MM4 N_XI0/XI58/XI4/NET33_XI0/XI58/XI4/MM4_d
+ N_XI0/XI58/XI4/NET34_XI0/XI58/XI4/MM4_g N_VDD_XI0/XI58/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI4/MM10 N_XI0/XI58/XI4/NET35_XI0/XI58/XI4/MM10_d
+ N_XI0/XI58/XI4/NET36_XI0/XI58/XI4/MM10_g N_VDD_XI0/XI58/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI4/MM11 N_XI0/XI58/XI4/NET36_XI0/XI58/XI4/MM11_d
+ N_XI0/XI58/XI4/NET35_XI0/XI58/XI4/MM11_g N_VDD_XI0/XI58/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI5/MM2 N_XI0/XI58/XI5/NET34_XI0/XI58/XI5/MM2_d
+ N_XI0/XI58/XI5/NET33_XI0/XI58/XI5/MM2_g N_VSS_XI0/XI58/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM3 N_XI0/XI58/XI5/NET33_XI0/XI58/XI5/MM3_d
+ N_WL<112>_XI0/XI58/XI5/MM3_g N_BLN<10>_XI0/XI58/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM0 N_XI0/XI58/XI5/NET34_XI0/XI58/XI5/MM0_d
+ N_WL<112>_XI0/XI58/XI5/MM0_g N_BL<10>_XI0/XI58/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM1 N_XI0/XI58/XI5/NET33_XI0/XI58/XI5/MM1_d
+ N_XI0/XI58/XI5/NET34_XI0/XI58/XI5/MM1_g N_VSS_XI0/XI58/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM9 N_XI0/XI58/XI5/NET36_XI0/XI58/XI5/MM9_d
+ N_WL<113>_XI0/XI58/XI5/MM9_g N_BL<10>_XI0/XI58/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM6 N_XI0/XI58/XI5/NET35_XI0/XI58/XI5/MM6_d
+ N_XI0/XI58/XI5/NET36_XI0/XI58/XI5/MM6_g N_VSS_XI0/XI58/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM7 N_XI0/XI58/XI5/NET36_XI0/XI58/XI5/MM7_d
+ N_XI0/XI58/XI5/NET35_XI0/XI58/XI5/MM7_g N_VSS_XI0/XI58/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM8 N_XI0/XI58/XI5/NET35_XI0/XI58/XI5/MM8_d
+ N_WL<113>_XI0/XI58/XI5/MM8_g N_BLN<10>_XI0/XI58/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI5/MM5 N_XI0/XI58/XI5/NET34_XI0/XI58/XI5/MM5_d
+ N_XI0/XI58/XI5/NET33_XI0/XI58/XI5/MM5_g N_VDD_XI0/XI58/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI5/MM4 N_XI0/XI58/XI5/NET33_XI0/XI58/XI5/MM4_d
+ N_XI0/XI58/XI5/NET34_XI0/XI58/XI5/MM4_g N_VDD_XI0/XI58/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI5/MM10 N_XI0/XI58/XI5/NET35_XI0/XI58/XI5/MM10_d
+ N_XI0/XI58/XI5/NET36_XI0/XI58/XI5/MM10_g N_VDD_XI0/XI58/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI5/MM11 N_XI0/XI58/XI5/NET36_XI0/XI58/XI5/MM11_d
+ N_XI0/XI58/XI5/NET35_XI0/XI58/XI5/MM11_g N_VDD_XI0/XI58/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI6/MM2 N_XI0/XI58/XI6/NET34_XI0/XI58/XI6/MM2_d
+ N_XI0/XI58/XI6/NET33_XI0/XI58/XI6/MM2_g N_VSS_XI0/XI58/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM3 N_XI0/XI58/XI6/NET33_XI0/XI58/XI6/MM3_d
+ N_WL<112>_XI0/XI58/XI6/MM3_g N_BLN<9>_XI0/XI58/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM0 N_XI0/XI58/XI6/NET34_XI0/XI58/XI6/MM0_d
+ N_WL<112>_XI0/XI58/XI6/MM0_g N_BL<9>_XI0/XI58/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM1 N_XI0/XI58/XI6/NET33_XI0/XI58/XI6/MM1_d
+ N_XI0/XI58/XI6/NET34_XI0/XI58/XI6/MM1_g N_VSS_XI0/XI58/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM9 N_XI0/XI58/XI6/NET36_XI0/XI58/XI6/MM9_d
+ N_WL<113>_XI0/XI58/XI6/MM9_g N_BL<9>_XI0/XI58/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM6 N_XI0/XI58/XI6/NET35_XI0/XI58/XI6/MM6_d
+ N_XI0/XI58/XI6/NET36_XI0/XI58/XI6/MM6_g N_VSS_XI0/XI58/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM7 N_XI0/XI58/XI6/NET36_XI0/XI58/XI6/MM7_d
+ N_XI0/XI58/XI6/NET35_XI0/XI58/XI6/MM7_g N_VSS_XI0/XI58/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM8 N_XI0/XI58/XI6/NET35_XI0/XI58/XI6/MM8_d
+ N_WL<113>_XI0/XI58/XI6/MM8_g N_BLN<9>_XI0/XI58/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI6/MM5 N_XI0/XI58/XI6/NET34_XI0/XI58/XI6/MM5_d
+ N_XI0/XI58/XI6/NET33_XI0/XI58/XI6/MM5_g N_VDD_XI0/XI58/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI6/MM4 N_XI0/XI58/XI6/NET33_XI0/XI58/XI6/MM4_d
+ N_XI0/XI58/XI6/NET34_XI0/XI58/XI6/MM4_g N_VDD_XI0/XI58/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI6/MM10 N_XI0/XI58/XI6/NET35_XI0/XI58/XI6/MM10_d
+ N_XI0/XI58/XI6/NET36_XI0/XI58/XI6/MM10_g N_VDD_XI0/XI58/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI6/MM11 N_XI0/XI58/XI6/NET36_XI0/XI58/XI6/MM11_d
+ N_XI0/XI58/XI6/NET35_XI0/XI58/XI6/MM11_g N_VDD_XI0/XI58/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI7/MM2 N_XI0/XI58/XI7/NET34_XI0/XI58/XI7/MM2_d
+ N_XI0/XI58/XI7/NET33_XI0/XI58/XI7/MM2_g N_VSS_XI0/XI58/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM3 N_XI0/XI58/XI7/NET33_XI0/XI58/XI7/MM3_d
+ N_WL<112>_XI0/XI58/XI7/MM3_g N_BLN<8>_XI0/XI58/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM0 N_XI0/XI58/XI7/NET34_XI0/XI58/XI7/MM0_d
+ N_WL<112>_XI0/XI58/XI7/MM0_g N_BL<8>_XI0/XI58/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM1 N_XI0/XI58/XI7/NET33_XI0/XI58/XI7/MM1_d
+ N_XI0/XI58/XI7/NET34_XI0/XI58/XI7/MM1_g N_VSS_XI0/XI58/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM9 N_XI0/XI58/XI7/NET36_XI0/XI58/XI7/MM9_d
+ N_WL<113>_XI0/XI58/XI7/MM9_g N_BL<8>_XI0/XI58/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM6 N_XI0/XI58/XI7/NET35_XI0/XI58/XI7/MM6_d
+ N_XI0/XI58/XI7/NET36_XI0/XI58/XI7/MM6_g N_VSS_XI0/XI58/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM7 N_XI0/XI58/XI7/NET36_XI0/XI58/XI7/MM7_d
+ N_XI0/XI58/XI7/NET35_XI0/XI58/XI7/MM7_g N_VSS_XI0/XI58/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM8 N_XI0/XI58/XI7/NET35_XI0/XI58/XI7/MM8_d
+ N_WL<113>_XI0/XI58/XI7/MM8_g N_BLN<8>_XI0/XI58/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI7/MM5 N_XI0/XI58/XI7/NET34_XI0/XI58/XI7/MM5_d
+ N_XI0/XI58/XI7/NET33_XI0/XI58/XI7/MM5_g N_VDD_XI0/XI58/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI7/MM4 N_XI0/XI58/XI7/NET33_XI0/XI58/XI7/MM4_d
+ N_XI0/XI58/XI7/NET34_XI0/XI58/XI7/MM4_g N_VDD_XI0/XI58/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI7/MM10 N_XI0/XI58/XI7/NET35_XI0/XI58/XI7/MM10_d
+ N_XI0/XI58/XI7/NET36_XI0/XI58/XI7/MM10_g N_VDD_XI0/XI58/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI7/MM11 N_XI0/XI58/XI7/NET36_XI0/XI58/XI7/MM11_d
+ N_XI0/XI58/XI7/NET35_XI0/XI58/XI7/MM11_g N_VDD_XI0/XI58/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI8/MM2 N_XI0/XI58/XI8/NET34_XI0/XI58/XI8/MM2_d
+ N_XI0/XI58/XI8/NET33_XI0/XI58/XI8/MM2_g N_VSS_XI0/XI58/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM3 N_XI0/XI58/XI8/NET33_XI0/XI58/XI8/MM3_d
+ N_WL<112>_XI0/XI58/XI8/MM3_g N_BLN<7>_XI0/XI58/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM0 N_XI0/XI58/XI8/NET34_XI0/XI58/XI8/MM0_d
+ N_WL<112>_XI0/XI58/XI8/MM0_g N_BL<7>_XI0/XI58/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM1 N_XI0/XI58/XI8/NET33_XI0/XI58/XI8/MM1_d
+ N_XI0/XI58/XI8/NET34_XI0/XI58/XI8/MM1_g N_VSS_XI0/XI58/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM9 N_XI0/XI58/XI8/NET36_XI0/XI58/XI8/MM9_d
+ N_WL<113>_XI0/XI58/XI8/MM9_g N_BL<7>_XI0/XI58/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM6 N_XI0/XI58/XI8/NET35_XI0/XI58/XI8/MM6_d
+ N_XI0/XI58/XI8/NET36_XI0/XI58/XI8/MM6_g N_VSS_XI0/XI58/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM7 N_XI0/XI58/XI8/NET36_XI0/XI58/XI8/MM7_d
+ N_XI0/XI58/XI8/NET35_XI0/XI58/XI8/MM7_g N_VSS_XI0/XI58/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM8 N_XI0/XI58/XI8/NET35_XI0/XI58/XI8/MM8_d
+ N_WL<113>_XI0/XI58/XI8/MM8_g N_BLN<7>_XI0/XI58/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI8/MM5 N_XI0/XI58/XI8/NET34_XI0/XI58/XI8/MM5_d
+ N_XI0/XI58/XI8/NET33_XI0/XI58/XI8/MM5_g N_VDD_XI0/XI58/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI8/MM4 N_XI0/XI58/XI8/NET33_XI0/XI58/XI8/MM4_d
+ N_XI0/XI58/XI8/NET34_XI0/XI58/XI8/MM4_g N_VDD_XI0/XI58/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI8/MM10 N_XI0/XI58/XI8/NET35_XI0/XI58/XI8/MM10_d
+ N_XI0/XI58/XI8/NET36_XI0/XI58/XI8/MM10_g N_VDD_XI0/XI58/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI8/MM11 N_XI0/XI58/XI8/NET36_XI0/XI58/XI8/MM11_d
+ N_XI0/XI58/XI8/NET35_XI0/XI58/XI8/MM11_g N_VDD_XI0/XI58/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI9/MM2 N_XI0/XI58/XI9/NET34_XI0/XI58/XI9/MM2_d
+ N_XI0/XI58/XI9/NET33_XI0/XI58/XI9/MM2_g N_VSS_XI0/XI58/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM3 N_XI0/XI58/XI9/NET33_XI0/XI58/XI9/MM3_d
+ N_WL<112>_XI0/XI58/XI9/MM3_g N_BLN<6>_XI0/XI58/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM0 N_XI0/XI58/XI9/NET34_XI0/XI58/XI9/MM0_d
+ N_WL<112>_XI0/XI58/XI9/MM0_g N_BL<6>_XI0/XI58/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM1 N_XI0/XI58/XI9/NET33_XI0/XI58/XI9/MM1_d
+ N_XI0/XI58/XI9/NET34_XI0/XI58/XI9/MM1_g N_VSS_XI0/XI58/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM9 N_XI0/XI58/XI9/NET36_XI0/XI58/XI9/MM9_d
+ N_WL<113>_XI0/XI58/XI9/MM9_g N_BL<6>_XI0/XI58/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM6 N_XI0/XI58/XI9/NET35_XI0/XI58/XI9/MM6_d
+ N_XI0/XI58/XI9/NET36_XI0/XI58/XI9/MM6_g N_VSS_XI0/XI58/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM7 N_XI0/XI58/XI9/NET36_XI0/XI58/XI9/MM7_d
+ N_XI0/XI58/XI9/NET35_XI0/XI58/XI9/MM7_g N_VSS_XI0/XI58/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM8 N_XI0/XI58/XI9/NET35_XI0/XI58/XI9/MM8_d
+ N_WL<113>_XI0/XI58/XI9/MM8_g N_BLN<6>_XI0/XI58/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI9/MM5 N_XI0/XI58/XI9/NET34_XI0/XI58/XI9/MM5_d
+ N_XI0/XI58/XI9/NET33_XI0/XI58/XI9/MM5_g N_VDD_XI0/XI58/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI9/MM4 N_XI0/XI58/XI9/NET33_XI0/XI58/XI9/MM4_d
+ N_XI0/XI58/XI9/NET34_XI0/XI58/XI9/MM4_g N_VDD_XI0/XI58/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI9/MM10 N_XI0/XI58/XI9/NET35_XI0/XI58/XI9/MM10_d
+ N_XI0/XI58/XI9/NET36_XI0/XI58/XI9/MM10_g N_VDD_XI0/XI58/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI9/MM11 N_XI0/XI58/XI9/NET36_XI0/XI58/XI9/MM11_d
+ N_XI0/XI58/XI9/NET35_XI0/XI58/XI9/MM11_g N_VDD_XI0/XI58/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI10/MM2 N_XI0/XI58/XI10/NET34_XI0/XI58/XI10/MM2_d
+ N_XI0/XI58/XI10/NET33_XI0/XI58/XI10/MM2_g N_VSS_XI0/XI58/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM3 N_XI0/XI58/XI10/NET33_XI0/XI58/XI10/MM3_d
+ N_WL<112>_XI0/XI58/XI10/MM3_g N_BLN<5>_XI0/XI58/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM0 N_XI0/XI58/XI10/NET34_XI0/XI58/XI10/MM0_d
+ N_WL<112>_XI0/XI58/XI10/MM0_g N_BL<5>_XI0/XI58/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM1 N_XI0/XI58/XI10/NET33_XI0/XI58/XI10/MM1_d
+ N_XI0/XI58/XI10/NET34_XI0/XI58/XI10/MM1_g N_VSS_XI0/XI58/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM9 N_XI0/XI58/XI10/NET36_XI0/XI58/XI10/MM9_d
+ N_WL<113>_XI0/XI58/XI10/MM9_g N_BL<5>_XI0/XI58/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM6 N_XI0/XI58/XI10/NET35_XI0/XI58/XI10/MM6_d
+ N_XI0/XI58/XI10/NET36_XI0/XI58/XI10/MM6_g N_VSS_XI0/XI58/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM7 N_XI0/XI58/XI10/NET36_XI0/XI58/XI10/MM7_d
+ N_XI0/XI58/XI10/NET35_XI0/XI58/XI10/MM7_g N_VSS_XI0/XI58/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM8 N_XI0/XI58/XI10/NET35_XI0/XI58/XI10/MM8_d
+ N_WL<113>_XI0/XI58/XI10/MM8_g N_BLN<5>_XI0/XI58/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI10/MM5 N_XI0/XI58/XI10/NET34_XI0/XI58/XI10/MM5_d
+ N_XI0/XI58/XI10/NET33_XI0/XI58/XI10/MM5_g N_VDD_XI0/XI58/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI10/MM4 N_XI0/XI58/XI10/NET33_XI0/XI58/XI10/MM4_d
+ N_XI0/XI58/XI10/NET34_XI0/XI58/XI10/MM4_g N_VDD_XI0/XI58/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI10/MM10 N_XI0/XI58/XI10/NET35_XI0/XI58/XI10/MM10_d
+ N_XI0/XI58/XI10/NET36_XI0/XI58/XI10/MM10_g N_VDD_XI0/XI58/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI10/MM11 N_XI0/XI58/XI10/NET36_XI0/XI58/XI10/MM11_d
+ N_XI0/XI58/XI10/NET35_XI0/XI58/XI10/MM11_g N_VDD_XI0/XI58/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI11/MM2 N_XI0/XI58/XI11/NET34_XI0/XI58/XI11/MM2_d
+ N_XI0/XI58/XI11/NET33_XI0/XI58/XI11/MM2_g N_VSS_XI0/XI58/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM3 N_XI0/XI58/XI11/NET33_XI0/XI58/XI11/MM3_d
+ N_WL<112>_XI0/XI58/XI11/MM3_g N_BLN<4>_XI0/XI58/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM0 N_XI0/XI58/XI11/NET34_XI0/XI58/XI11/MM0_d
+ N_WL<112>_XI0/XI58/XI11/MM0_g N_BL<4>_XI0/XI58/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM1 N_XI0/XI58/XI11/NET33_XI0/XI58/XI11/MM1_d
+ N_XI0/XI58/XI11/NET34_XI0/XI58/XI11/MM1_g N_VSS_XI0/XI58/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM9 N_XI0/XI58/XI11/NET36_XI0/XI58/XI11/MM9_d
+ N_WL<113>_XI0/XI58/XI11/MM9_g N_BL<4>_XI0/XI58/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM6 N_XI0/XI58/XI11/NET35_XI0/XI58/XI11/MM6_d
+ N_XI0/XI58/XI11/NET36_XI0/XI58/XI11/MM6_g N_VSS_XI0/XI58/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM7 N_XI0/XI58/XI11/NET36_XI0/XI58/XI11/MM7_d
+ N_XI0/XI58/XI11/NET35_XI0/XI58/XI11/MM7_g N_VSS_XI0/XI58/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM8 N_XI0/XI58/XI11/NET35_XI0/XI58/XI11/MM8_d
+ N_WL<113>_XI0/XI58/XI11/MM8_g N_BLN<4>_XI0/XI58/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI11/MM5 N_XI0/XI58/XI11/NET34_XI0/XI58/XI11/MM5_d
+ N_XI0/XI58/XI11/NET33_XI0/XI58/XI11/MM5_g N_VDD_XI0/XI58/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI11/MM4 N_XI0/XI58/XI11/NET33_XI0/XI58/XI11/MM4_d
+ N_XI0/XI58/XI11/NET34_XI0/XI58/XI11/MM4_g N_VDD_XI0/XI58/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI11/MM10 N_XI0/XI58/XI11/NET35_XI0/XI58/XI11/MM10_d
+ N_XI0/XI58/XI11/NET36_XI0/XI58/XI11/MM10_g N_VDD_XI0/XI58/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI11/MM11 N_XI0/XI58/XI11/NET36_XI0/XI58/XI11/MM11_d
+ N_XI0/XI58/XI11/NET35_XI0/XI58/XI11/MM11_g N_VDD_XI0/XI58/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI12/MM2 N_XI0/XI58/XI12/NET34_XI0/XI58/XI12/MM2_d
+ N_XI0/XI58/XI12/NET33_XI0/XI58/XI12/MM2_g N_VSS_XI0/XI58/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM3 N_XI0/XI58/XI12/NET33_XI0/XI58/XI12/MM3_d
+ N_WL<112>_XI0/XI58/XI12/MM3_g N_BLN<3>_XI0/XI58/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM0 N_XI0/XI58/XI12/NET34_XI0/XI58/XI12/MM0_d
+ N_WL<112>_XI0/XI58/XI12/MM0_g N_BL<3>_XI0/XI58/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM1 N_XI0/XI58/XI12/NET33_XI0/XI58/XI12/MM1_d
+ N_XI0/XI58/XI12/NET34_XI0/XI58/XI12/MM1_g N_VSS_XI0/XI58/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM9 N_XI0/XI58/XI12/NET36_XI0/XI58/XI12/MM9_d
+ N_WL<113>_XI0/XI58/XI12/MM9_g N_BL<3>_XI0/XI58/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM6 N_XI0/XI58/XI12/NET35_XI0/XI58/XI12/MM6_d
+ N_XI0/XI58/XI12/NET36_XI0/XI58/XI12/MM6_g N_VSS_XI0/XI58/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM7 N_XI0/XI58/XI12/NET36_XI0/XI58/XI12/MM7_d
+ N_XI0/XI58/XI12/NET35_XI0/XI58/XI12/MM7_g N_VSS_XI0/XI58/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM8 N_XI0/XI58/XI12/NET35_XI0/XI58/XI12/MM8_d
+ N_WL<113>_XI0/XI58/XI12/MM8_g N_BLN<3>_XI0/XI58/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI12/MM5 N_XI0/XI58/XI12/NET34_XI0/XI58/XI12/MM5_d
+ N_XI0/XI58/XI12/NET33_XI0/XI58/XI12/MM5_g N_VDD_XI0/XI58/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI12/MM4 N_XI0/XI58/XI12/NET33_XI0/XI58/XI12/MM4_d
+ N_XI0/XI58/XI12/NET34_XI0/XI58/XI12/MM4_g N_VDD_XI0/XI58/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI12/MM10 N_XI0/XI58/XI12/NET35_XI0/XI58/XI12/MM10_d
+ N_XI0/XI58/XI12/NET36_XI0/XI58/XI12/MM10_g N_VDD_XI0/XI58/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI12/MM11 N_XI0/XI58/XI12/NET36_XI0/XI58/XI12/MM11_d
+ N_XI0/XI58/XI12/NET35_XI0/XI58/XI12/MM11_g N_VDD_XI0/XI58/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI13/MM2 N_XI0/XI58/XI13/NET34_XI0/XI58/XI13/MM2_d
+ N_XI0/XI58/XI13/NET33_XI0/XI58/XI13/MM2_g N_VSS_XI0/XI58/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM3 N_XI0/XI58/XI13/NET33_XI0/XI58/XI13/MM3_d
+ N_WL<112>_XI0/XI58/XI13/MM3_g N_BLN<2>_XI0/XI58/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM0 N_XI0/XI58/XI13/NET34_XI0/XI58/XI13/MM0_d
+ N_WL<112>_XI0/XI58/XI13/MM0_g N_BL<2>_XI0/XI58/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM1 N_XI0/XI58/XI13/NET33_XI0/XI58/XI13/MM1_d
+ N_XI0/XI58/XI13/NET34_XI0/XI58/XI13/MM1_g N_VSS_XI0/XI58/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM9 N_XI0/XI58/XI13/NET36_XI0/XI58/XI13/MM9_d
+ N_WL<113>_XI0/XI58/XI13/MM9_g N_BL<2>_XI0/XI58/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM6 N_XI0/XI58/XI13/NET35_XI0/XI58/XI13/MM6_d
+ N_XI0/XI58/XI13/NET36_XI0/XI58/XI13/MM6_g N_VSS_XI0/XI58/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM7 N_XI0/XI58/XI13/NET36_XI0/XI58/XI13/MM7_d
+ N_XI0/XI58/XI13/NET35_XI0/XI58/XI13/MM7_g N_VSS_XI0/XI58/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM8 N_XI0/XI58/XI13/NET35_XI0/XI58/XI13/MM8_d
+ N_WL<113>_XI0/XI58/XI13/MM8_g N_BLN<2>_XI0/XI58/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI13/MM5 N_XI0/XI58/XI13/NET34_XI0/XI58/XI13/MM5_d
+ N_XI0/XI58/XI13/NET33_XI0/XI58/XI13/MM5_g N_VDD_XI0/XI58/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI13/MM4 N_XI0/XI58/XI13/NET33_XI0/XI58/XI13/MM4_d
+ N_XI0/XI58/XI13/NET34_XI0/XI58/XI13/MM4_g N_VDD_XI0/XI58/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI13/MM10 N_XI0/XI58/XI13/NET35_XI0/XI58/XI13/MM10_d
+ N_XI0/XI58/XI13/NET36_XI0/XI58/XI13/MM10_g N_VDD_XI0/XI58/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI13/MM11 N_XI0/XI58/XI13/NET36_XI0/XI58/XI13/MM11_d
+ N_XI0/XI58/XI13/NET35_XI0/XI58/XI13/MM11_g N_VDD_XI0/XI58/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI14/MM2 N_XI0/XI58/XI14/NET34_XI0/XI58/XI14/MM2_d
+ N_XI0/XI58/XI14/NET33_XI0/XI58/XI14/MM2_g N_VSS_XI0/XI58/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM3 N_XI0/XI58/XI14/NET33_XI0/XI58/XI14/MM3_d
+ N_WL<112>_XI0/XI58/XI14/MM3_g N_BLN<1>_XI0/XI58/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM0 N_XI0/XI58/XI14/NET34_XI0/XI58/XI14/MM0_d
+ N_WL<112>_XI0/XI58/XI14/MM0_g N_BL<1>_XI0/XI58/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM1 N_XI0/XI58/XI14/NET33_XI0/XI58/XI14/MM1_d
+ N_XI0/XI58/XI14/NET34_XI0/XI58/XI14/MM1_g N_VSS_XI0/XI58/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM9 N_XI0/XI58/XI14/NET36_XI0/XI58/XI14/MM9_d
+ N_WL<113>_XI0/XI58/XI14/MM9_g N_BL<1>_XI0/XI58/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM6 N_XI0/XI58/XI14/NET35_XI0/XI58/XI14/MM6_d
+ N_XI0/XI58/XI14/NET36_XI0/XI58/XI14/MM6_g N_VSS_XI0/XI58/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM7 N_XI0/XI58/XI14/NET36_XI0/XI58/XI14/MM7_d
+ N_XI0/XI58/XI14/NET35_XI0/XI58/XI14/MM7_g N_VSS_XI0/XI58/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM8 N_XI0/XI58/XI14/NET35_XI0/XI58/XI14/MM8_d
+ N_WL<113>_XI0/XI58/XI14/MM8_g N_BLN<1>_XI0/XI58/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI14/MM5 N_XI0/XI58/XI14/NET34_XI0/XI58/XI14/MM5_d
+ N_XI0/XI58/XI14/NET33_XI0/XI58/XI14/MM5_g N_VDD_XI0/XI58/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI14/MM4 N_XI0/XI58/XI14/NET33_XI0/XI58/XI14/MM4_d
+ N_XI0/XI58/XI14/NET34_XI0/XI58/XI14/MM4_g N_VDD_XI0/XI58/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI14/MM10 N_XI0/XI58/XI14/NET35_XI0/XI58/XI14/MM10_d
+ N_XI0/XI58/XI14/NET36_XI0/XI58/XI14/MM10_g N_VDD_XI0/XI58/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI14/MM11 N_XI0/XI58/XI14/NET36_XI0/XI58/XI14/MM11_d
+ N_XI0/XI58/XI14/NET35_XI0/XI58/XI14/MM11_g N_VDD_XI0/XI58/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI15/MM2 N_XI0/XI58/XI15/NET34_XI0/XI58/XI15/MM2_d
+ N_XI0/XI58/XI15/NET33_XI0/XI58/XI15/MM2_g N_VSS_XI0/XI58/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM3 N_XI0/XI58/XI15/NET33_XI0/XI58/XI15/MM3_d
+ N_WL<112>_XI0/XI58/XI15/MM3_g N_BLN<0>_XI0/XI58/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM0 N_XI0/XI58/XI15/NET34_XI0/XI58/XI15/MM0_d
+ N_WL<112>_XI0/XI58/XI15/MM0_g N_BL<0>_XI0/XI58/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM1 N_XI0/XI58/XI15/NET33_XI0/XI58/XI15/MM1_d
+ N_XI0/XI58/XI15/NET34_XI0/XI58/XI15/MM1_g N_VSS_XI0/XI58/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM9 N_XI0/XI58/XI15/NET36_XI0/XI58/XI15/MM9_d
+ N_WL<113>_XI0/XI58/XI15/MM9_g N_BL<0>_XI0/XI58/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM6 N_XI0/XI58/XI15/NET35_XI0/XI58/XI15/MM6_d
+ N_XI0/XI58/XI15/NET36_XI0/XI58/XI15/MM6_g N_VSS_XI0/XI58/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM7 N_XI0/XI58/XI15/NET36_XI0/XI58/XI15/MM7_d
+ N_XI0/XI58/XI15/NET35_XI0/XI58/XI15/MM7_g N_VSS_XI0/XI58/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM8 N_XI0/XI58/XI15/NET35_XI0/XI58/XI15/MM8_d
+ N_WL<113>_XI0/XI58/XI15/MM8_g N_BLN<0>_XI0/XI58/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI58/XI15/MM5 N_XI0/XI58/XI15/NET34_XI0/XI58/XI15/MM5_d
+ N_XI0/XI58/XI15/NET33_XI0/XI58/XI15/MM5_g N_VDD_XI0/XI58/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI15/MM4 N_XI0/XI58/XI15/NET33_XI0/XI58/XI15/MM4_d
+ N_XI0/XI58/XI15/NET34_XI0/XI58/XI15/MM4_g N_VDD_XI0/XI58/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI15/MM10 N_XI0/XI58/XI15/NET35_XI0/XI58/XI15/MM10_d
+ N_XI0/XI58/XI15/NET36_XI0/XI58/XI15/MM10_g N_VDD_XI0/XI58/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI58/XI15/MM11 N_XI0/XI58/XI15/NET36_XI0/XI58/XI15/MM11_d
+ N_XI0/XI58/XI15/NET35_XI0/XI58/XI15/MM11_g N_VDD_XI0/XI58/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI0/MM2 N_XI0/XI59/XI0/NET34_XI0/XI59/XI0/MM2_d
+ N_XI0/XI59/XI0/NET33_XI0/XI59/XI0/MM2_g N_VSS_XI0/XI59/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM3 N_XI0/XI59/XI0/NET33_XI0/XI59/XI0/MM3_d
+ N_WL<114>_XI0/XI59/XI0/MM3_g N_BLN<15>_XI0/XI59/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM0 N_XI0/XI59/XI0/NET34_XI0/XI59/XI0/MM0_d
+ N_WL<114>_XI0/XI59/XI0/MM0_g N_BL<15>_XI0/XI59/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM1 N_XI0/XI59/XI0/NET33_XI0/XI59/XI0/MM1_d
+ N_XI0/XI59/XI0/NET34_XI0/XI59/XI0/MM1_g N_VSS_XI0/XI59/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM9 N_XI0/XI59/XI0/NET36_XI0/XI59/XI0/MM9_d
+ N_WL<115>_XI0/XI59/XI0/MM9_g N_BL<15>_XI0/XI59/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM6 N_XI0/XI59/XI0/NET35_XI0/XI59/XI0/MM6_d
+ N_XI0/XI59/XI0/NET36_XI0/XI59/XI0/MM6_g N_VSS_XI0/XI59/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM7 N_XI0/XI59/XI0/NET36_XI0/XI59/XI0/MM7_d
+ N_XI0/XI59/XI0/NET35_XI0/XI59/XI0/MM7_g N_VSS_XI0/XI59/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM8 N_XI0/XI59/XI0/NET35_XI0/XI59/XI0/MM8_d
+ N_WL<115>_XI0/XI59/XI0/MM8_g N_BLN<15>_XI0/XI59/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI0/MM5 N_XI0/XI59/XI0/NET34_XI0/XI59/XI0/MM5_d
+ N_XI0/XI59/XI0/NET33_XI0/XI59/XI0/MM5_g N_VDD_XI0/XI59/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI0/MM4 N_XI0/XI59/XI0/NET33_XI0/XI59/XI0/MM4_d
+ N_XI0/XI59/XI0/NET34_XI0/XI59/XI0/MM4_g N_VDD_XI0/XI59/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI0/MM10 N_XI0/XI59/XI0/NET35_XI0/XI59/XI0/MM10_d
+ N_XI0/XI59/XI0/NET36_XI0/XI59/XI0/MM10_g N_VDD_XI0/XI59/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI0/MM11 N_XI0/XI59/XI0/NET36_XI0/XI59/XI0/MM11_d
+ N_XI0/XI59/XI0/NET35_XI0/XI59/XI0/MM11_g N_VDD_XI0/XI59/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI1/MM2 N_XI0/XI59/XI1/NET34_XI0/XI59/XI1/MM2_d
+ N_XI0/XI59/XI1/NET33_XI0/XI59/XI1/MM2_g N_VSS_XI0/XI59/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM3 N_XI0/XI59/XI1/NET33_XI0/XI59/XI1/MM3_d
+ N_WL<114>_XI0/XI59/XI1/MM3_g N_BLN<14>_XI0/XI59/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM0 N_XI0/XI59/XI1/NET34_XI0/XI59/XI1/MM0_d
+ N_WL<114>_XI0/XI59/XI1/MM0_g N_BL<14>_XI0/XI59/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM1 N_XI0/XI59/XI1/NET33_XI0/XI59/XI1/MM1_d
+ N_XI0/XI59/XI1/NET34_XI0/XI59/XI1/MM1_g N_VSS_XI0/XI59/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM9 N_XI0/XI59/XI1/NET36_XI0/XI59/XI1/MM9_d
+ N_WL<115>_XI0/XI59/XI1/MM9_g N_BL<14>_XI0/XI59/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM6 N_XI0/XI59/XI1/NET35_XI0/XI59/XI1/MM6_d
+ N_XI0/XI59/XI1/NET36_XI0/XI59/XI1/MM6_g N_VSS_XI0/XI59/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM7 N_XI0/XI59/XI1/NET36_XI0/XI59/XI1/MM7_d
+ N_XI0/XI59/XI1/NET35_XI0/XI59/XI1/MM7_g N_VSS_XI0/XI59/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM8 N_XI0/XI59/XI1/NET35_XI0/XI59/XI1/MM8_d
+ N_WL<115>_XI0/XI59/XI1/MM8_g N_BLN<14>_XI0/XI59/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI1/MM5 N_XI0/XI59/XI1/NET34_XI0/XI59/XI1/MM5_d
+ N_XI0/XI59/XI1/NET33_XI0/XI59/XI1/MM5_g N_VDD_XI0/XI59/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI1/MM4 N_XI0/XI59/XI1/NET33_XI0/XI59/XI1/MM4_d
+ N_XI0/XI59/XI1/NET34_XI0/XI59/XI1/MM4_g N_VDD_XI0/XI59/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI1/MM10 N_XI0/XI59/XI1/NET35_XI0/XI59/XI1/MM10_d
+ N_XI0/XI59/XI1/NET36_XI0/XI59/XI1/MM10_g N_VDD_XI0/XI59/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI1/MM11 N_XI0/XI59/XI1/NET36_XI0/XI59/XI1/MM11_d
+ N_XI0/XI59/XI1/NET35_XI0/XI59/XI1/MM11_g N_VDD_XI0/XI59/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI2/MM2 N_XI0/XI59/XI2/NET34_XI0/XI59/XI2/MM2_d
+ N_XI0/XI59/XI2/NET33_XI0/XI59/XI2/MM2_g N_VSS_XI0/XI59/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM3 N_XI0/XI59/XI2/NET33_XI0/XI59/XI2/MM3_d
+ N_WL<114>_XI0/XI59/XI2/MM3_g N_BLN<13>_XI0/XI59/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM0 N_XI0/XI59/XI2/NET34_XI0/XI59/XI2/MM0_d
+ N_WL<114>_XI0/XI59/XI2/MM0_g N_BL<13>_XI0/XI59/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM1 N_XI0/XI59/XI2/NET33_XI0/XI59/XI2/MM1_d
+ N_XI0/XI59/XI2/NET34_XI0/XI59/XI2/MM1_g N_VSS_XI0/XI59/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM9 N_XI0/XI59/XI2/NET36_XI0/XI59/XI2/MM9_d
+ N_WL<115>_XI0/XI59/XI2/MM9_g N_BL<13>_XI0/XI59/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM6 N_XI0/XI59/XI2/NET35_XI0/XI59/XI2/MM6_d
+ N_XI0/XI59/XI2/NET36_XI0/XI59/XI2/MM6_g N_VSS_XI0/XI59/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM7 N_XI0/XI59/XI2/NET36_XI0/XI59/XI2/MM7_d
+ N_XI0/XI59/XI2/NET35_XI0/XI59/XI2/MM7_g N_VSS_XI0/XI59/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM8 N_XI0/XI59/XI2/NET35_XI0/XI59/XI2/MM8_d
+ N_WL<115>_XI0/XI59/XI2/MM8_g N_BLN<13>_XI0/XI59/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI2/MM5 N_XI0/XI59/XI2/NET34_XI0/XI59/XI2/MM5_d
+ N_XI0/XI59/XI2/NET33_XI0/XI59/XI2/MM5_g N_VDD_XI0/XI59/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI2/MM4 N_XI0/XI59/XI2/NET33_XI0/XI59/XI2/MM4_d
+ N_XI0/XI59/XI2/NET34_XI0/XI59/XI2/MM4_g N_VDD_XI0/XI59/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI2/MM10 N_XI0/XI59/XI2/NET35_XI0/XI59/XI2/MM10_d
+ N_XI0/XI59/XI2/NET36_XI0/XI59/XI2/MM10_g N_VDD_XI0/XI59/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI2/MM11 N_XI0/XI59/XI2/NET36_XI0/XI59/XI2/MM11_d
+ N_XI0/XI59/XI2/NET35_XI0/XI59/XI2/MM11_g N_VDD_XI0/XI59/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI3/MM2 N_XI0/XI59/XI3/NET34_XI0/XI59/XI3/MM2_d
+ N_XI0/XI59/XI3/NET33_XI0/XI59/XI3/MM2_g N_VSS_XI0/XI59/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM3 N_XI0/XI59/XI3/NET33_XI0/XI59/XI3/MM3_d
+ N_WL<114>_XI0/XI59/XI3/MM3_g N_BLN<12>_XI0/XI59/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM0 N_XI0/XI59/XI3/NET34_XI0/XI59/XI3/MM0_d
+ N_WL<114>_XI0/XI59/XI3/MM0_g N_BL<12>_XI0/XI59/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM1 N_XI0/XI59/XI3/NET33_XI0/XI59/XI3/MM1_d
+ N_XI0/XI59/XI3/NET34_XI0/XI59/XI3/MM1_g N_VSS_XI0/XI59/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM9 N_XI0/XI59/XI3/NET36_XI0/XI59/XI3/MM9_d
+ N_WL<115>_XI0/XI59/XI3/MM9_g N_BL<12>_XI0/XI59/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM6 N_XI0/XI59/XI3/NET35_XI0/XI59/XI3/MM6_d
+ N_XI0/XI59/XI3/NET36_XI0/XI59/XI3/MM6_g N_VSS_XI0/XI59/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM7 N_XI0/XI59/XI3/NET36_XI0/XI59/XI3/MM7_d
+ N_XI0/XI59/XI3/NET35_XI0/XI59/XI3/MM7_g N_VSS_XI0/XI59/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM8 N_XI0/XI59/XI3/NET35_XI0/XI59/XI3/MM8_d
+ N_WL<115>_XI0/XI59/XI3/MM8_g N_BLN<12>_XI0/XI59/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI3/MM5 N_XI0/XI59/XI3/NET34_XI0/XI59/XI3/MM5_d
+ N_XI0/XI59/XI3/NET33_XI0/XI59/XI3/MM5_g N_VDD_XI0/XI59/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI3/MM4 N_XI0/XI59/XI3/NET33_XI0/XI59/XI3/MM4_d
+ N_XI0/XI59/XI3/NET34_XI0/XI59/XI3/MM4_g N_VDD_XI0/XI59/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI3/MM10 N_XI0/XI59/XI3/NET35_XI0/XI59/XI3/MM10_d
+ N_XI0/XI59/XI3/NET36_XI0/XI59/XI3/MM10_g N_VDD_XI0/XI59/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI3/MM11 N_XI0/XI59/XI3/NET36_XI0/XI59/XI3/MM11_d
+ N_XI0/XI59/XI3/NET35_XI0/XI59/XI3/MM11_g N_VDD_XI0/XI59/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI4/MM2 N_XI0/XI59/XI4/NET34_XI0/XI59/XI4/MM2_d
+ N_XI0/XI59/XI4/NET33_XI0/XI59/XI4/MM2_g N_VSS_XI0/XI59/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM3 N_XI0/XI59/XI4/NET33_XI0/XI59/XI4/MM3_d
+ N_WL<114>_XI0/XI59/XI4/MM3_g N_BLN<11>_XI0/XI59/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM0 N_XI0/XI59/XI4/NET34_XI0/XI59/XI4/MM0_d
+ N_WL<114>_XI0/XI59/XI4/MM0_g N_BL<11>_XI0/XI59/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM1 N_XI0/XI59/XI4/NET33_XI0/XI59/XI4/MM1_d
+ N_XI0/XI59/XI4/NET34_XI0/XI59/XI4/MM1_g N_VSS_XI0/XI59/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM9 N_XI0/XI59/XI4/NET36_XI0/XI59/XI4/MM9_d
+ N_WL<115>_XI0/XI59/XI4/MM9_g N_BL<11>_XI0/XI59/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM6 N_XI0/XI59/XI4/NET35_XI0/XI59/XI4/MM6_d
+ N_XI0/XI59/XI4/NET36_XI0/XI59/XI4/MM6_g N_VSS_XI0/XI59/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM7 N_XI0/XI59/XI4/NET36_XI0/XI59/XI4/MM7_d
+ N_XI0/XI59/XI4/NET35_XI0/XI59/XI4/MM7_g N_VSS_XI0/XI59/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM8 N_XI0/XI59/XI4/NET35_XI0/XI59/XI4/MM8_d
+ N_WL<115>_XI0/XI59/XI4/MM8_g N_BLN<11>_XI0/XI59/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI4/MM5 N_XI0/XI59/XI4/NET34_XI0/XI59/XI4/MM5_d
+ N_XI0/XI59/XI4/NET33_XI0/XI59/XI4/MM5_g N_VDD_XI0/XI59/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI4/MM4 N_XI0/XI59/XI4/NET33_XI0/XI59/XI4/MM4_d
+ N_XI0/XI59/XI4/NET34_XI0/XI59/XI4/MM4_g N_VDD_XI0/XI59/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI4/MM10 N_XI0/XI59/XI4/NET35_XI0/XI59/XI4/MM10_d
+ N_XI0/XI59/XI4/NET36_XI0/XI59/XI4/MM10_g N_VDD_XI0/XI59/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI4/MM11 N_XI0/XI59/XI4/NET36_XI0/XI59/XI4/MM11_d
+ N_XI0/XI59/XI4/NET35_XI0/XI59/XI4/MM11_g N_VDD_XI0/XI59/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI5/MM2 N_XI0/XI59/XI5/NET34_XI0/XI59/XI5/MM2_d
+ N_XI0/XI59/XI5/NET33_XI0/XI59/XI5/MM2_g N_VSS_XI0/XI59/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM3 N_XI0/XI59/XI5/NET33_XI0/XI59/XI5/MM3_d
+ N_WL<114>_XI0/XI59/XI5/MM3_g N_BLN<10>_XI0/XI59/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM0 N_XI0/XI59/XI5/NET34_XI0/XI59/XI5/MM0_d
+ N_WL<114>_XI0/XI59/XI5/MM0_g N_BL<10>_XI0/XI59/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM1 N_XI0/XI59/XI5/NET33_XI0/XI59/XI5/MM1_d
+ N_XI0/XI59/XI5/NET34_XI0/XI59/XI5/MM1_g N_VSS_XI0/XI59/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM9 N_XI0/XI59/XI5/NET36_XI0/XI59/XI5/MM9_d
+ N_WL<115>_XI0/XI59/XI5/MM9_g N_BL<10>_XI0/XI59/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM6 N_XI0/XI59/XI5/NET35_XI0/XI59/XI5/MM6_d
+ N_XI0/XI59/XI5/NET36_XI0/XI59/XI5/MM6_g N_VSS_XI0/XI59/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM7 N_XI0/XI59/XI5/NET36_XI0/XI59/XI5/MM7_d
+ N_XI0/XI59/XI5/NET35_XI0/XI59/XI5/MM7_g N_VSS_XI0/XI59/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM8 N_XI0/XI59/XI5/NET35_XI0/XI59/XI5/MM8_d
+ N_WL<115>_XI0/XI59/XI5/MM8_g N_BLN<10>_XI0/XI59/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI5/MM5 N_XI0/XI59/XI5/NET34_XI0/XI59/XI5/MM5_d
+ N_XI0/XI59/XI5/NET33_XI0/XI59/XI5/MM5_g N_VDD_XI0/XI59/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI5/MM4 N_XI0/XI59/XI5/NET33_XI0/XI59/XI5/MM4_d
+ N_XI0/XI59/XI5/NET34_XI0/XI59/XI5/MM4_g N_VDD_XI0/XI59/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI5/MM10 N_XI0/XI59/XI5/NET35_XI0/XI59/XI5/MM10_d
+ N_XI0/XI59/XI5/NET36_XI0/XI59/XI5/MM10_g N_VDD_XI0/XI59/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI5/MM11 N_XI0/XI59/XI5/NET36_XI0/XI59/XI5/MM11_d
+ N_XI0/XI59/XI5/NET35_XI0/XI59/XI5/MM11_g N_VDD_XI0/XI59/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI6/MM2 N_XI0/XI59/XI6/NET34_XI0/XI59/XI6/MM2_d
+ N_XI0/XI59/XI6/NET33_XI0/XI59/XI6/MM2_g N_VSS_XI0/XI59/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM3 N_XI0/XI59/XI6/NET33_XI0/XI59/XI6/MM3_d
+ N_WL<114>_XI0/XI59/XI6/MM3_g N_BLN<9>_XI0/XI59/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM0 N_XI0/XI59/XI6/NET34_XI0/XI59/XI6/MM0_d
+ N_WL<114>_XI0/XI59/XI6/MM0_g N_BL<9>_XI0/XI59/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM1 N_XI0/XI59/XI6/NET33_XI0/XI59/XI6/MM1_d
+ N_XI0/XI59/XI6/NET34_XI0/XI59/XI6/MM1_g N_VSS_XI0/XI59/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM9 N_XI0/XI59/XI6/NET36_XI0/XI59/XI6/MM9_d
+ N_WL<115>_XI0/XI59/XI6/MM9_g N_BL<9>_XI0/XI59/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM6 N_XI0/XI59/XI6/NET35_XI0/XI59/XI6/MM6_d
+ N_XI0/XI59/XI6/NET36_XI0/XI59/XI6/MM6_g N_VSS_XI0/XI59/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM7 N_XI0/XI59/XI6/NET36_XI0/XI59/XI6/MM7_d
+ N_XI0/XI59/XI6/NET35_XI0/XI59/XI6/MM7_g N_VSS_XI0/XI59/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM8 N_XI0/XI59/XI6/NET35_XI0/XI59/XI6/MM8_d
+ N_WL<115>_XI0/XI59/XI6/MM8_g N_BLN<9>_XI0/XI59/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI6/MM5 N_XI0/XI59/XI6/NET34_XI0/XI59/XI6/MM5_d
+ N_XI0/XI59/XI6/NET33_XI0/XI59/XI6/MM5_g N_VDD_XI0/XI59/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI6/MM4 N_XI0/XI59/XI6/NET33_XI0/XI59/XI6/MM4_d
+ N_XI0/XI59/XI6/NET34_XI0/XI59/XI6/MM4_g N_VDD_XI0/XI59/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI6/MM10 N_XI0/XI59/XI6/NET35_XI0/XI59/XI6/MM10_d
+ N_XI0/XI59/XI6/NET36_XI0/XI59/XI6/MM10_g N_VDD_XI0/XI59/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI6/MM11 N_XI0/XI59/XI6/NET36_XI0/XI59/XI6/MM11_d
+ N_XI0/XI59/XI6/NET35_XI0/XI59/XI6/MM11_g N_VDD_XI0/XI59/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI7/MM2 N_XI0/XI59/XI7/NET34_XI0/XI59/XI7/MM2_d
+ N_XI0/XI59/XI7/NET33_XI0/XI59/XI7/MM2_g N_VSS_XI0/XI59/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM3 N_XI0/XI59/XI7/NET33_XI0/XI59/XI7/MM3_d
+ N_WL<114>_XI0/XI59/XI7/MM3_g N_BLN<8>_XI0/XI59/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM0 N_XI0/XI59/XI7/NET34_XI0/XI59/XI7/MM0_d
+ N_WL<114>_XI0/XI59/XI7/MM0_g N_BL<8>_XI0/XI59/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM1 N_XI0/XI59/XI7/NET33_XI0/XI59/XI7/MM1_d
+ N_XI0/XI59/XI7/NET34_XI0/XI59/XI7/MM1_g N_VSS_XI0/XI59/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM9 N_XI0/XI59/XI7/NET36_XI0/XI59/XI7/MM9_d
+ N_WL<115>_XI0/XI59/XI7/MM9_g N_BL<8>_XI0/XI59/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM6 N_XI0/XI59/XI7/NET35_XI0/XI59/XI7/MM6_d
+ N_XI0/XI59/XI7/NET36_XI0/XI59/XI7/MM6_g N_VSS_XI0/XI59/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM7 N_XI0/XI59/XI7/NET36_XI0/XI59/XI7/MM7_d
+ N_XI0/XI59/XI7/NET35_XI0/XI59/XI7/MM7_g N_VSS_XI0/XI59/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM8 N_XI0/XI59/XI7/NET35_XI0/XI59/XI7/MM8_d
+ N_WL<115>_XI0/XI59/XI7/MM8_g N_BLN<8>_XI0/XI59/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI7/MM5 N_XI0/XI59/XI7/NET34_XI0/XI59/XI7/MM5_d
+ N_XI0/XI59/XI7/NET33_XI0/XI59/XI7/MM5_g N_VDD_XI0/XI59/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI7/MM4 N_XI0/XI59/XI7/NET33_XI0/XI59/XI7/MM4_d
+ N_XI0/XI59/XI7/NET34_XI0/XI59/XI7/MM4_g N_VDD_XI0/XI59/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI7/MM10 N_XI0/XI59/XI7/NET35_XI0/XI59/XI7/MM10_d
+ N_XI0/XI59/XI7/NET36_XI0/XI59/XI7/MM10_g N_VDD_XI0/XI59/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI7/MM11 N_XI0/XI59/XI7/NET36_XI0/XI59/XI7/MM11_d
+ N_XI0/XI59/XI7/NET35_XI0/XI59/XI7/MM11_g N_VDD_XI0/XI59/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI8/MM2 N_XI0/XI59/XI8/NET34_XI0/XI59/XI8/MM2_d
+ N_XI0/XI59/XI8/NET33_XI0/XI59/XI8/MM2_g N_VSS_XI0/XI59/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM3 N_XI0/XI59/XI8/NET33_XI0/XI59/XI8/MM3_d
+ N_WL<114>_XI0/XI59/XI8/MM3_g N_BLN<7>_XI0/XI59/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM0 N_XI0/XI59/XI8/NET34_XI0/XI59/XI8/MM0_d
+ N_WL<114>_XI0/XI59/XI8/MM0_g N_BL<7>_XI0/XI59/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM1 N_XI0/XI59/XI8/NET33_XI0/XI59/XI8/MM1_d
+ N_XI0/XI59/XI8/NET34_XI0/XI59/XI8/MM1_g N_VSS_XI0/XI59/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM9 N_XI0/XI59/XI8/NET36_XI0/XI59/XI8/MM9_d
+ N_WL<115>_XI0/XI59/XI8/MM9_g N_BL<7>_XI0/XI59/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM6 N_XI0/XI59/XI8/NET35_XI0/XI59/XI8/MM6_d
+ N_XI0/XI59/XI8/NET36_XI0/XI59/XI8/MM6_g N_VSS_XI0/XI59/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM7 N_XI0/XI59/XI8/NET36_XI0/XI59/XI8/MM7_d
+ N_XI0/XI59/XI8/NET35_XI0/XI59/XI8/MM7_g N_VSS_XI0/XI59/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM8 N_XI0/XI59/XI8/NET35_XI0/XI59/XI8/MM8_d
+ N_WL<115>_XI0/XI59/XI8/MM8_g N_BLN<7>_XI0/XI59/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI8/MM5 N_XI0/XI59/XI8/NET34_XI0/XI59/XI8/MM5_d
+ N_XI0/XI59/XI8/NET33_XI0/XI59/XI8/MM5_g N_VDD_XI0/XI59/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI8/MM4 N_XI0/XI59/XI8/NET33_XI0/XI59/XI8/MM4_d
+ N_XI0/XI59/XI8/NET34_XI0/XI59/XI8/MM4_g N_VDD_XI0/XI59/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI8/MM10 N_XI0/XI59/XI8/NET35_XI0/XI59/XI8/MM10_d
+ N_XI0/XI59/XI8/NET36_XI0/XI59/XI8/MM10_g N_VDD_XI0/XI59/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI8/MM11 N_XI0/XI59/XI8/NET36_XI0/XI59/XI8/MM11_d
+ N_XI0/XI59/XI8/NET35_XI0/XI59/XI8/MM11_g N_VDD_XI0/XI59/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI9/MM2 N_XI0/XI59/XI9/NET34_XI0/XI59/XI9/MM2_d
+ N_XI0/XI59/XI9/NET33_XI0/XI59/XI9/MM2_g N_VSS_XI0/XI59/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM3 N_XI0/XI59/XI9/NET33_XI0/XI59/XI9/MM3_d
+ N_WL<114>_XI0/XI59/XI9/MM3_g N_BLN<6>_XI0/XI59/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM0 N_XI0/XI59/XI9/NET34_XI0/XI59/XI9/MM0_d
+ N_WL<114>_XI0/XI59/XI9/MM0_g N_BL<6>_XI0/XI59/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM1 N_XI0/XI59/XI9/NET33_XI0/XI59/XI9/MM1_d
+ N_XI0/XI59/XI9/NET34_XI0/XI59/XI9/MM1_g N_VSS_XI0/XI59/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM9 N_XI0/XI59/XI9/NET36_XI0/XI59/XI9/MM9_d
+ N_WL<115>_XI0/XI59/XI9/MM9_g N_BL<6>_XI0/XI59/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM6 N_XI0/XI59/XI9/NET35_XI0/XI59/XI9/MM6_d
+ N_XI0/XI59/XI9/NET36_XI0/XI59/XI9/MM6_g N_VSS_XI0/XI59/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM7 N_XI0/XI59/XI9/NET36_XI0/XI59/XI9/MM7_d
+ N_XI0/XI59/XI9/NET35_XI0/XI59/XI9/MM7_g N_VSS_XI0/XI59/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM8 N_XI0/XI59/XI9/NET35_XI0/XI59/XI9/MM8_d
+ N_WL<115>_XI0/XI59/XI9/MM8_g N_BLN<6>_XI0/XI59/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI9/MM5 N_XI0/XI59/XI9/NET34_XI0/XI59/XI9/MM5_d
+ N_XI0/XI59/XI9/NET33_XI0/XI59/XI9/MM5_g N_VDD_XI0/XI59/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI9/MM4 N_XI0/XI59/XI9/NET33_XI0/XI59/XI9/MM4_d
+ N_XI0/XI59/XI9/NET34_XI0/XI59/XI9/MM4_g N_VDD_XI0/XI59/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI9/MM10 N_XI0/XI59/XI9/NET35_XI0/XI59/XI9/MM10_d
+ N_XI0/XI59/XI9/NET36_XI0/XI59/XI9/MM10_g N_VDD_XI0/XI59/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI9/MM11 N_XI0/XI59/XI9/NET36_XI0/XI59/XI9/MM11_d
+ N_XI0/XI59/XI9/NET35_XI0/XI59/XI9/MM11_g N_VDD_XI0/XI59/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI10/MM2 N_XI0/XI59/XI10/NET34_XI0/XI59/XI10/MM2_d
+ N_XI0/XI59/XI10/NET33_XI0/XI59/XI10/MM2_g N_VSS_XI0/XI59/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM3 N_XI0/XI59/XI10/NET33_XI0/XI59/XI10/MM3_d
+ N_WL<114>_XI0/XI59/XI10/MM3_g N_BLN<5>_XI0/XI59/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM0 N_XI0/XI59/XI10/NET34_XI0/XI59/XI10/MM0_d
+ N_WL<114>_XI0/XI59/XI10/MM0_g N_BL<5>_XI0/XI59/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM1 N_XI0/XI59/XI10/NET33_XI0/XI59/XI10/MM1_d
+ N_XI0/XI59/XI10/NET34_XI0/XI59/XI10/MM1_g N_VSS_XI0/XI59/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM9 N_XI0/XI59/XI10/NET36_XI0/XI59/XI10/MM9_d
+ N_WL<115>_XI0/XI59/XI10/MM9_g N_BL<5>_XI0/XI59/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM6 N_XI0/XI59/XI10/NET35_XI0/XI59/XI10/MM6_d
+ N_XI0/XI59/XI10/NET36_XI0/XI59/XI10/MM6_g N_VSS_XI0/XI59/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM7 N_XI0/XI59/XI10/NET36_XI0/XI59/XI10/MM7_d
+ N_XI0/XI59/XI10/NET35_XI0/XI59/XI10/MM7_g N_VSS_XI0/XI59/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM8 N_XI0/XI59/XI10/NET35_XI0/XI59/XI10/MM8_d
+ N_WL<115>_XI0/XI59/XI10/MM8_g N_BLN<5>_XI0/XI59/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI10/MM5 N_XI0/XI59/XI10/NET34_XI0/XI59/XI10/MM5_d
+ N_XI0/XI59/XI10/NET33_XI0/XI59/XI10/MM5_g N_VDD_XI0/XI59/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI10/MM4 N_XI0/XI59/XI10/NET33_XI0/XI59/XI10/MM4_d
+ N_XI0/XI59/XI10/NET34_XI0/XI59/XI10/MM4_g N_VDD_XI0/XI59/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI10/MM10 N_XI0/XI59/XI10/NET35_XI0/XI59/XI10/MM10_d
+ N_XI0/XI59/XI10/NET36_XI0/XI59/XI10/MM10_g N_VDD_XI0/XI59/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI10/MM11 N_XI0/XI59/XI10/NET36_XI0/XI59/XI10/MM11_d
+ N_XI0/XI59/XI10/NET35_XI0/XI59/XI10/MM11_g N_VDD_XI0/XI59/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI11/MM2 N_XI0/XI59/XI11/NET34_XI0/XI59/XI11/MM2_d
+ N_XI0/XI59/XI11/NET33_XI0/XI59/XI11/MM2_g N_VSS_XI0/XI59/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM3 N_XI0/XI59/XI11/NET33_XI0/XI59/XI11/MM3_d
+ N_WL<114>_XI0/XI59/XI11/MM3_g N_BLN<4>_XI0/XI59/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM0 N_XI0/XI59/XI11/NET34_XI0/XI59/XI11/MM0_d
+ N_WL<114>_XI0/XI59/XI11/MM0_g N_BL<4>_XI0/XI59/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM1 N_XI0/XI59/XI11/NET33_XI0/XI59/XI11/MM1_d
+ N_XI0/XI59/XI11/NET34_XI0/XI59/XI11/MM1_g N_VSS_XI0/XI59/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM9 N_XI0/XI59/XI11/NET36_XI0/XI59/XI11/MM9_d
+ N_WL<115>_XI0/XI59/XI11/MM9_g N_BL<4>_XI0/XI59/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM6 N_XI0/XI59/XI11/NET35_XI0/XI59/XI11/MM6_d
+ N_XI0/XI59/XI11/NET36_XI0/XI59/XI11/MM6_g N_VSS_XI0/XI59/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM7 N_XI0/XI59/XI11/NET36_XI0/XI59/XI11/MM7_d
+ N_XI0/XI59/XI11/NET35_XI0/XI59/XI11/MM7_g N_VSS_XI0/XI59/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM8 N_XI0/XI59/XI11/NET35_XI0/XI59/XI11/MM8_d
+ N_WL<115>_XI0/XI59/XI11/MM8_g N_BLN<4>_XI0/XI59/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI11/MM5 N_XI0/XI59/XI11/NET34_XI0/XI59/XI11/MM5_d
+ N_XI0/XI59/XI11/NET33_XI0/XI59/XI11/MM5_g N_VDD_XI0/XI59/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI11/MM4 N_XI0/XI59/XI11/NET33_XI0/XI59/XI11/MM4_d
+ N_XI0/XI59/XI11/NET34_XI0/XI59/XI11/MM4_g N_VDD_XI0/XI59/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI11/MM10 N_XI0/XI59/XI11/NET35_XI0/XI59/XI11/MM10_d
+ N_XI0/XI59/XI11/NET36_XI0/XI59/XI11/MM10_g N_VDD_XI0/XI59/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI11/MM11 N_XI0/XI59/XI11/NET36_XI0/XI59/XI11/MM11_d
+ N_XI0/XI59/XI11/NET35_XI0/XI59/XI11/MM11_g N_VDD_XI0/XI59/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI12/MM2 N_XI0/XI59/XI12/NET34_XI0/XI59/XI12/MM2_d
+ N_XI0/XI59/XI12/NET33_XI0/XI59/XI12/MM2_g N_VSS_XI0/XI59/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM3 N_XI0/XI59/XI12/NET33_XI0/XI59/XI12/MM3_d
+ N_WL<114>_XI0/XI59/XI12/MM3_g N_BLN<3>_XI0/XI59/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM0 N_XI0/XI59/XI12/NET34_XI0/XI59/XI12/MM0_d
+ N_WL<114>_XI0/XI59/XI12/MM0_g N_BL<3>_XI0/XI59/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM1 N_XI0/XI59/XI12/NET33_XI0/XI59/XI12/MM1_d
+ N_XI0/XI59/XI12/NET34_XI0/XI59/XI12/MM1_g N_VSS_XI0/XI59/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM9 N_XI0/XI59/XI12/NET36_XI0/XI59/XI12/MM9_d
+ N_WL<115>_XI0/XI59/XI12/MM9_g N_BL<3>_XI0/XI59/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM6 N_XI0/XI59/XI12/NET35_XI0/XI59/XI12/MM6_d
+ N_XI0/XI59/XI12/NET36_XI0/XI59/XI12/MM6_g N_VSS_XI0/XI59/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM7 N_XI0/XI59/XI12/NET36_XI0/XI59/XI12/MM7_d
+ N_XI0/XI59/XI12/NET35_XI0/XI59/XI12/MM7_g N_VSS_XI0/XI59/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM8 N_XI0/XI59/XI12/NET35_XI0/XI59/XI12/MM8_d
+ N_WL<115>_XI0/XI59/XI12/MM8_g N_BLN<3>_XI0/XI59/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI12/MM5 N_XI0/XI59/XI12/NET34_XI0/XI59/XI12/MM5_d
+ N_XI0/XI59/XI12/NET33_XI0/XI59/XI12/MM5_g N_VDD_XI0/XI59/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI12/MM4 N_XI0/XI59/XI12/NET33_XI0/XI59/XI12/MM4_d
+ N_XI0/XI59/XI12/NET34_XI0/XI59/XI12/MM4_g N_VDD_XI0/XI59/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI12/MM10 N_XI0/XI59/XI12/NET35_XI0/XI59/XI12/MM10_d
+ N_XI0/XI59/XI12/NET36_XI0/XI59/XI12/MM10_g N_VDD_XI0/XI59/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI12/MM11 N_XI0/XI59/XI12/NET36_XI0/XI59/XI12/MM11_d
+ N_XI0/XI59/XI12/NET35_XI0/XI59/XI12/MM11_g N_VDD_XI0/XI59/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI13/MM2 N_XI0/XI59/XI13/NET34_XI0/XI59/XI13/MM2_d
+ N_XI0/XI59/XI13/NET33_XI0/XI59/XI13/MM2_g N_VSS_XI0/XI59/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM3 N_XI0/XI59/XI13/NET33_XI0/XI59/XI13/MM3_d
+ N_WL<114>_XI0/XI59/XI13/MM3_g N_BLN<2>_XI0/XI59/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM0 N_XI0/XI59/XI13/NET34_XI0/XI59/XI13/MM0_d
+ N_WL<114>_XI0/XI59/XI13/MM0_g N_BL<2>_XI0/XI59/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM1 N_XI0/XI59/XI13/NET33_XI0/XI59/XI13/MM1_d
+ N_XI0/XI59/XI13/NET34_XI0/XI59/XI13/MM1_g N_VSS_XI0/XI59/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM9 N_XI0/XI59/XI13/NET36_XI0/XI59/XI13/MM9_d
+ N_WL<115>_XI0/XI59/XI13/MM9_g N_BL<2>_XI0/XI59/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM6 N_XI0/XI59/XI13/NET35_XI0/XI59/XI13/MM6_d
+ N_XI0/XI59/XI13/NET36_XI0/XI59/XI13/MM6_g N_VSS_XI0/XI59/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM7 N_XI0/XI59/XI13/NET36_XI0/XI59/XI13/MM7_d
+ N_XI0/XI59/XI13/NET35_XI0/XI59/XI13/MM7_g N_VSS_XI0/XI59/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM8 N_XI0/XI59/XI13/NET35_XI0/XI59/XI13/MM8_d
+ N_WL<115>_XI0/XI59/XI13/MM8_g N_BLN<2>_XI0/XI59/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI13/MM5 N_XI0/XI59/XI13/NET34_XI0/XI59/XI13/MM5_d
+ N_XI0/XI59/XI13/NET33_XI0/XI59/XI13/MM5_g N_VDD_XI0/XI59/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI13/MM4 N_XI0/XI59/XI13/NET33_XI0/XI59/XI13/MM4_d
+ N_XI0/XI59/XI13/NET34_XI0/XI59/XI13/MM4_g N_VDD_XI0/XI59/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI13/MM10 N_XI0/XI59/XI13/NET35_XI0/XI59/XI13/MM10_d
+ N_XI0/XI59/XI13/NET36_XI0/XI59/XI13/MM10_g N_VDD_XI0/XI59/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI13/MM11 N_XI0/XI59/XI13/NET36_XI0/XI59/XI13/MM11_d
+ N_XI0/XI59/XI13/NET35_XI0/XI59/XI13/MM11_g N_VDD_XI0/XI59/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI14/MM2 N_XI0/XI59/XI14/NET34_XI0/XI59/XI14/MM2_d
+ N_XI0/XI59/XI14/NET33_XI0/XI59/XI14/MM2_g N_VSS_XI0/XI59/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM3 N_XI0/XI59/XI14/NET33_XI0/XI59/XI14/MM3_d
+ N_WL<114>_XI0/XI59/XI14/MM3_g N_BLN<1>_XI0/XI59/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM0 N_XI0/XI59/XI14/NET34_XI0/XI59/XI14/MM0_d
+ N_WL<114>_XI0/XI59/XI14/MM0_g N_BL<1>_XI0/XI59/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM1 N_XI0/XI59/XI14/NET33_XI0/XI59/XI14/MM1_d
+ N_XI0/XI59/XI14/NET34_XI0/XI59/XI14/MM1_g N_VSS_XI0/XI59/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM9 N_XI0/XI59/XI14/NET36_XI0/XI59/XI14/MM9_d
+ N_WL<115>_XI0/XI59/XI14/MM9_g N_BL<1>_XI0/XI59/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM6 N_XI0/XI59/XI14/NET35_XI0/XI59/XI14/MM6_d
+ N_XI0/XI59/XI14/NET36_XI0/XI59/XI14/MM6_g N_VSS_XI0/XI59/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM7 N_XI0/XI59/XI14/NET36_XI0/XI59/XI14/MM7_d
+ N_XI0/XI59/XI14/NET35_XI0/XI59/XI14/MM7_g N_VSS_XI0/XI59/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM8 N_XI0/XI59/XI14/NET35_XI0/XI59/XI14/MM8_d
+ N_WL<115>_XI0/XI59/XI14/MM8_g N_BLN<1>_XI0/XI59/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI14/MM5 N_XI0/XI59/XI14/NET34_XI0/XI59/XI14/MM5_d
+ N_XI0/XI59/XI14/NET33_XI0/XI59/XI14/MM5_g N_VDD_XI0/XI59/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI14/MM4 N_XI0/XI59/XI14/NET33_XI0/XI59/XI14/MM4_d
+ N_XI0/XI59/XI14/NET34_XI0/XI59/XI14/MM4_g N_VDD_XI0/XI59/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI14/MM10 N_XI0/XI59/XI14/NET35_XI0/XI59/XI14/MM10_d
+ N_XI0/XI59/XI14/NET36_XI0/XI59/XI14/MM10_g N_VDD_XI0/XI59/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI14/MM11 N_XI0/XI59/XI14/NET36_XI0/XI59/XI14/MM11_d
+ N_XI0/XI59/XI14/NET35_XI0/XI59/XI14/MM11_g N_VDD_XI0/XI59/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI15/MM2 N_XI0/XI59/XI15/NET34_XI0/XI59/XI15/MM2_d
+ N_XI0/XI59/XI15/NET33_XI0/XI59/XI15/MM2_g N_VSS_XI0/XI59/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM3 N_XI0/XI59/XI15/NET33_XI0/XI59/XI15/MM3_d
+ N_WL<114>_XI0/XI59/XI15/MM3_g N_BLN<0>_XI0/XI59/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM0 N_XI0/XI59/XI15/NET34_XI0/XI59/XI15/MM0_d
+ N_WL<114>_XI0/XI59/XI15/MM0_g N_BL<0>_XI0/XI59/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM1 N_XI0/XI59/XI15/NET33_XI0/XI59/XI15/MM1_d
+ N_XI0/XI59/XI15/NET34_XI0/XI59/XI15/MM1_g N_VSS_XI0/XI59/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM9 N_XI0/XI59/XI15/NET36_XI0/XI59/XI15/MM9_d
+ N_WL<115>_XI0/XI59/XI15/MM9_g N_BL<0>_XI0/XI59/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM6 N_XI0/XI59/XI15/NET35_XI0/XI59/XI15/MM6_d
+ N_XI0/XI59/XI15/NET36_XI0/XI59/XI15/MM6_g N_VSS_XI0/XI59/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM7 N_XI0/XI59/XI15/NET36_XI0/XI59/XI15/MM7_d
+ N_XI0/XI59/XI15/NET35_XI0/XI59/XI15/MM7_g N_VSS_XI0/XI59/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM8 N_XI0/XI59/XI15/NET35_XI0/XI59/XI15/MM8_d
+ N_WL<115>_XI0/XI59/XI15/MM8_g N_BLN<0>_XI0/XI59/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI59/XI15/MM5 N_XI0/XI59/XI15/NET34_XI0/XI59/XI15/MM5_d
+ N_XI0/XI59/XI15/NET33_XI0/XI59/XI15/MM5_g N_VDD_XI0/XI59/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI15/MM4 N_XI0/XI59/XI15/NET33_XI0/XI59/XI15/MM4_d
+ N_XI0/XI59/XI15/NET34_XI0/XI59/XI15/MM4_g N_VDD_XI0/XI59/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI15/MM10 N_XI0/XI59/XI15/NET35_XI0/XI59/XI15/MM10_d
+ N_XI0/XI59/XI15/NET36_XI0/XI59/XI15/MM10_g N_VDD_XI0/XI59/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI59/XI15/MM11 N_XI0/XI59/XI15/NET36_XI0/XI59/XI15/MM11_d
+ N_XI0/XI59/XI15/NET35_XI0/XI59/XI15/MM11_g N_VDD_XI0/XI59/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI0/MM2 N_XI0/XI60/XI0/NET34_XI0/XI60/XI0/MM2_d
+ N_XI0/XI60/XI0/NET33_XI0/XI60/XI0/MM2_g N_VSS_XI0/XI60/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM3 N_XI0/XI60/XI0/NET33_XI0/XI60/XI0/MM3_d
+ N_WL<116>_XI0/XI60/XI0/MM3_g N_BLN<15>_XI0/XI60/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM0 N_XI0/XI60/XI0/NET34_XI0/XI60/XI0/MM0_d
+ N_WL<116>_XI0/XI60/XI0/MM0_g N_BL<15>_XI0/XI60/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM1 N_XI0/XI60/XI0/NET33_XI0/XI60/XI0/MM1_d
+ N_XI0/XI60/XI0/NET34_XI0/XI60/XI0/MM1_g N_VSS_XI0/XI60/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM9 N_XI0/XI60/XI0/NET36_XI0/XI60/XI0/MM9_d
+ N_WL<117>_XI0/XI60/XI0/MM9_g N_BL<15>_XI0/XI60/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM6 N_XI0/XI60/XI0/NET35_XI0/XI60/XI0/MM6_d
+ N_XI0/XI60/XI0/NET36_XI0/XI60/XI0/MM6_g N_VSS_XI0/XI60/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM7 N_XI0/XI60/XI0/NET36_XI0/XI60/XI0/MM7_d
+ N_XI0/XI60/XI0/NET35_XI0/XI60/XI0/MM7_g N_VSS_XI0/XI60/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM8 N_XI0/XI60/XI0/NET35_XI0/XI60/XI0/MM8_d
+ N_WL<117>_XI0/XI60/XI0/MM8_g N_BLN<15>_XI0/XI60/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI0/MM5 N_XI0/XI60/XI0/NET34_XI0/XI60/XI0/MM5_d
+ N_XI0/XI60/XI0/NET33_XI0/XI60/XI0/MM5_g N_VDD_XI0/XI60/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI0/MM4 N_XI0/XI60/XI0/NET33_XI0/XI60/XI0/MM4_d
+ N_XI0/XI60/XI0/NET34_XI0/XI60/XI0/MM4_g N_VDD_XI0/XI60/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI0/MM10 N_XI0/XI60/XI0/NET35_XI0/XI60/XI0/MM10_d
+ N_XI0/XI60/XI0/NET36_XI0/XI60/XI0/MM10_g N_VDD_XI0/XI60/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI0/MM11 N_XI0/XI60/XI0/NET36_XI0/XI60/XI0/MM11_d
+ N_XI0/XI60/XI0/NET35_XI0/XI60/XI0/MM11_g N_VDD_XI0/XI60/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI1/MM2 N_XI0/XI60/XI1/NET34_XI0/XI60/XI1/MM2_d
+ N_XI0/XI60/XI1/NET33_XI0/XI60/XI1/MM2_g N_VSS_XI0/XI60/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM3 N_XI0/XI60/XI1/NET33_XI0/XI60/XI1/MM3_d
+ N_WL<116>_XI0/XI60/XI1/MM3_g N_BLN<14>_XI0/XI60/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM0 N_XI0/XI60/XI1/NET34_XI0/XI60/XI1/MM0_d
+ N_WL<116>_XI0/XI60/XI1/MM0_g N_BL<14>_XI0/XI60/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM1 N_XI0/XI60/XI1/NET33_XI0/XI60/XI1/MM1_d
+ N_XI0/XI60/XI1/NET34_XI0/XI60/XI1/MM1_g N_VSS_XI0/XI60/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM9 N_XI0/XI60/XI1/NET36_XI0/XI60/XI1/MM9_d
+ N_WL<117>_XI0/XI60/XI1/MM9_g N_BL<14>_XI0/XI60/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM6 N_XI0/XI60/XI1/NET35_XI0/XI60/XI1/MM6_d
+ N_XI0/XI60/XI1/NET36_XI0/XI60/XI1/MM6_g N_VSS_XI0/XI60/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM7 N_XI0/XI60/XI1/NET36_XI0/XI60/XI1/MM7_d
+ N_XI0/XI60/XI1/NET35_XI0/XI60/XI1/MM7_g N_VSS_XI0/XI60/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM8 N_XI0/XI60/XI1/NET35_XI0/XI60/XI1/MM8_d
+ N_WL<117>_XI0/XI60/XI1/MM8_g N_BLN<14>_XI0/XI60/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI1/MM5 N_XI0/XI60/XI1/NET34_XI0/XI60/XI1/MM5_d
+ N_XI0/XI60/XI1/NET33_XI0/XI60/XI1/MM5_g N_VDD_XI0/XI60/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI1/MM4 N_XI0/XI60/XI1/NET33_XI0/XI60/XI1/MM4_d
+ N_XI0/XI60/XI1/NET34_XI0/XI60/XI1/MM4_g N_VDD_XI0/XI60/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI1/MM10 N_XI0/XI60/XI1/NET35_XI0/XI60/XI1/MM10_d
+ N_XI0/XI60/XI1/NET36_XI0/XI60/XI1/MM10_g N_VDD_XI0/XI60/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI1/MM11 N_XI0/XI60/XI1/NET36_XI0/XI60/XI1/MM11_d
+ N_XI0/XI60/XI1/NET35_XI0/XI60/XI1/MM11_g N_VDD_XI0/XI60/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI2/MM2 N_XI0/XI60/XI2/NET34_XI0/XI60/XI2/MM2_d
+ N_XI0/XI60/XI2/NET33_XI0/XI60/XI2/MM2_g N_VSS_XI0/XI60/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM3 N_XI0/XI60/XI2/NET33_XI0/XI60/XI2/MM3_d
+ N_WL<116>_XI0/XI60/XI2/MM3_g N_BLN<13>_XI0/XI60/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM0 N_XI0/XI60/XI2/NET34_XI0/XI60/XI2/MM0_d
+ N_WL<116>_XI0/XI60/XI2/MM0_g N_BL<13>_XI0/XI60/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM1 N_XI0/XI60/XI2/NET33_XI0/XI60/XI2/MM1_d
+ N_XI0/XI60/XI2/NET34_XI0/XI60/XI2/MM1_g N_VSS_XI0/XI60/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM9 N_XI0/XI60/XI2/NET36_XI0/XI60/XI2/MM9_d
+ N_WL<117>_XI0/XI60/XI2/MM9_g N_BL<13>_XI0/XI60/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM6 N_XI0/XI60/XI2/NET35_XI0/XI60/XI2/MM6_d
+ N_XI0/XI60/XI2/NET36_XI0/XI60/XI2/MM6_g N_VSS_XI0/XI60/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM7 N_XI0/XI60/XI2/NET36_XI0/XI60/XI2/MM7_d
+ N_XI0/XI60/XI2/NET35_XI0/XI60/XI2/MM7_g N_VSS_XI0/XI60/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM8 N_XI0/XI60/XI2/NET35_XI0/XI60/XI2/MM8_d
+ N_WL<117>_XI0/XI60/XI2/MM8_g N_BLN<13>_XI0/XI60/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI2/MM5 N_XI0/XI60/XI2/NET34_XI0/XI60/XI2/MM5_d
+ N_XI0/XI60/XI2/NET33_XI0/XI60/XI2/MM5_g N_VDD_XI0/XI60/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI2/MM4 N_XI0/XI60/XI2/NET33_XI0/XI60/XI2/MM4_d
+ N_XI0/XI60/XI2/NET34_XI0/XI60/XI2/MM4_g N_VDD_XI0/XI60/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI2/MM10 N_XI0/XI60/XI2/NET35_XI0/XI60/XI2/MM10_d
+ N_XI0/XI60/XI2/NET36_XI0/XI60/XI2/MM10_g N_VDD_XI0/XI60/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI2/MM11 N_XI0/XI60/XI2/NET36_XI0/XI60/XI2/MM11_d
+ N_XI0/XI60/XI2/NET35_XI0/XI60/XI2/MM11_g N_VDD_XI0/XI60/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI3/MM2 N_XI0/XI60/XI3/NET34_XI0/XI60/XI3/MM2_d
+ N_XI0/XI60/XI3/NET33_XI0/XI60/XI3/MM2_g N_VSS_XI0/XI60/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM3 N_XI0/XI60/XI3/NET33_XI0/XI60/XI3/MM3_d
+ N_WL<116>_XI0/XI60/XI3/MM3_g N_BLN<12>_XI0/XI60/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM0 N_XI0/XI60/XI3/NET34_XI0/XI60/XI3/MM0_d
+ N_WL<116>_XI0/XI60/XI3/MM0_g N_BL<12>_XI0/XI60/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM1 N_XI0/XI60/XI3/NET33_XI0/XI60/XI3/MM1_d
+ N_XI0/XI60/XI3/NET34_XI0/XI60/XI3/MM1_g N_VSS_XI0/XI60/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM9 N_XI0/XI60/XI3/NET36_XI0/XI60/XI3/MM9_d
+ N_WL<117>_XI0/XI60/XI3/MM9_g N_BL<12>_XI0/XI60/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM6 N_XI0/XI60/XI3/NET35_XI0/XI60/XI3/MM6_d
+ N_XI0/XI60/XI3/NET36_XI0/XI60/XI3/MM6_g N_VSS_XI0/XI60/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM7 N_XI0/XI60/XI3/NET36_XI0/XI60/XI3/MM7_d
+ N_XI0/XI60/XI3/NET35_XI0/XI60/XI3/MM7_g N_VSS_XI0/XI60/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM8 N_XI0/XI60/XI3/NET35_XI0/XI60/XI3/MM8_d
+ N_WL<117>_XI0/XI60/XI3/MM8_g N_BLN<12>_XI0/XI60/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI3/MM5 N_XI0/XI60/XI3/NET34_XI0/XI60/XI3/MM5_d
+ N_XI0/XI60/XI3/NET33_XI0/XI60/XI3/MM5_g N_VDD_XI0/XI60/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI3/MM4 N_XI0/XI60/XI3/NET33_XI0/XI60/XI3/MM4_d
+ N_XI0/XI60/XI3/NET34_XI0/XI60/XI3/MM4_g N_VDD_XI0/XI60/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI3/MM10 N_XI0/XI60/XI3/NET35_XI0/XI60/XI3/MM10_d
+ N_XI0/XI60/XI3/NET36_XI0/XI60/XI3/MM10_g N_VDD_XI0/XI60/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI3/MM11 N_XI0/XI60/XI3/NET36_XI0/XI60/XI3/MM11_d
+ N_XI0/XI60/XI3/NET35_XI0/XI60/XI3/MM11_g N_VDD_XI0/XI60/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI4/MM2 N_XI0/XI60/XI4/NET34_XI0/XI60/XI4/MM2_d
+ N_XI0/XI60/XI4/NET33_XI0/XI60/XI4/MM2_g N_VSS_XI0/XI60/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM3 N_XI0/XI60/XI4/NET33_XI0/XI60/XI4/MM3_d
+ N_WL<116>_XI0/XI60/XI4/MM3_g N_BLN<11>_XI0/XI60/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM0 N_XI0/XI60/XI4/NET34_XI0/XI60/XI4/MM0_d
+ N_WL<116>_XI0/XI60/XI4/MM0_g N_BL<11>_XI0/XI60/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM1 N_XI0/XI60/XI4/NET33_XI0/XI60/XI4/MM1_d
+ N_XI0/XI60/XI4/NET34_XI0/XI60/XI4/MM1_g N_VSS_XI0/XI60/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM9 N_XI0/XI60/XI4/NET36_XI0/XI60/XI4/MM9_d
+ N_WL<117>_XI0/XI60/XI4/MM9_g N_BL<11>_XI0/XI60/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM6 N_XI0/XI60/XI4/NET35_XI0/XI60/XI4/MM6_d
+ N_XI0/XI60/XI4/NET36_XI0/XI60/XI4/MM6_g N_VSS_XI0/XI60/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM7 N_XI0/XI60/XI4/NET36_XI0/XI60/XI4/MM7_d
+ N_XI0/XI60/XI4/NET35_XI0/XI60/XI4/MM7_g N_VSS_XI0/XI60/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM8 N_XI0/XI60/XI4/NET35_XI0/XI60/XI4/MM8_d
+ N_WL<117>_XI0/XI60/XI4/MM8_g N_BLN<11>_XI0/XI60/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI4/MM5 N_XI0/XI60/XI4/NET34_XI0/XI60/XI4/MM5_d
+ N_XI0/XI60/XI4/NET33_XI0/XI60/XI4/MM5_g N_VDD_XI0/XI60/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI4/MM4 N_XI0/XI60/XI4/NET33_XI0/XI60/XI4/MM4_d
+ N_XI0/XI60/XI4/NET34_XI0/XI60/XI4/MM4_g N_VDD_XI0/XI60/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI4/MM10 N_XI0/XI60/XI4/NET35_XI0/XI60/XI4/MM10_d
+ N_XI0/XI60/XI4/NET36_XI0/XI60/XI4/MM10_g N_VDD_XI0/XI60/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI4/MM11 N_XI0/XI60/XI4/NET36_XI0/XI60/XI4/MM11_d
+ N_XI0/XI60/XI4/NET35_XI0/XI60/XI4/MM11_g N_VDD_XI0/XI60/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI5/MM2 N_XI0/XI60/XI5/NET34_XI0/XI60/XI5/MM2_d
+ N_XI0/XI60/XI5/NET33_XI0/XI60/XI5/MM2_g N_VSS_XI0/XI60/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM3 N_XI0/XI60/XI5/NET33_XI0/XI60/XI5/MM3_d
+ N_WL<116>_XI0/XI60/XI5/MM3_g N_BLN<10>_XI0/XI60/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM0 N_XI0/XI60/XI5/NET34_XI0/XI60/XI5/MM0_d
+ N_WL<116>_XI0/XI60/XI5/MM0_g N_BL<10>_XI0/XI60/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM1 N_XI0/XI60/XI5/NET33_XI0/XI60/XI5/MM1_d
+ N_XI0/XI60/XI5/NET34_XI0/XI60/XI5/MM1_g N_VSS_XI0/XI60/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM9 N_XI0/XI60/XI5/NET36_XI0/XI60/XI5/MM9_d
+ N_WL<117>_XI0/XI60/XI5/MM9_g N_BL<10>_XI0/XI60/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM6 N_XI0/XI60/XI5/NET35_XI0/XI60/XI5/MM6_d
+ N_XI0/XI60/XI5/NET36_XI0/XI60/XI5/MM6_g N_VSS_XI0/XI60/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM7 N_XI0/XI60/XI5/NET36_XI0/XI60/XI5/MM7_d
+ N_XI0/XI60/XI5/NET35_XI0/XI60/XI5/MM7_g N_VSS_XI0/XI60/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM8 N_XI0/XI60/XI5/NET35_XI0/XI60/XI5/MM8_d
+ N_WL<117>_XI0/XI60/XI5/MM8_g N_BLN<10>_XI0/XI60/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI5/MM5 N_XI0/XI60/XI5/NET34_XI0/XI60/XI5/MM5_d
+ N_XI0/XI60/XI5/NET33_XI0/XI60/XI5/MM5_g N_VDD_XI0/XI60/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI5/MM4 N_XI0/XI60/XI5/NET33_XI0/XI60/XI5/MM4_d
+ N_XI0/XI60/XI5/NET34_XI0/XI60/XI5/MM4_g N_VDD_XI0/XI60/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI5/MM10 N_XI0/XI60/XI5/NET35_XI0/XI60/XI5/MM10_d
+ N_XI0/XI60/XI5/NET36_XI0/XI60/XI5/MM10_g N_VDD_XI0/XI60/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI5/MM11 N_XI0/XI60/XI5/NET36_XI0/XI60/XI5/MM11_d
+ N_XI0/XI60/XI5/NET35_XI0/XI60/XI5/MM11_g N_VDD_XI0/XI60/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI6/MM2 N_XI0/XI60/XI6/NET34_XI0/XI60/XI6/MM2_d
+ N_XI0/XI60/XI6/NET33_XI0/XI60/XI6/MM2_g N_VSS_XI0/XI60/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM3 N_XI0/XI60/XI6/NET33_XI0/XI60/XI6/MM3_d
+ N_WL<116>_XI0/XI60/XI6/MM3_g N_BLN<9>_XI0/XI60/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM0 N_XI0/XI60/XI6/NET34_XI0/XI60/XI6/MM0_d
+ N_WL<116>_XI0/XI60/XI6/MM0_g N_BL<9>_XI0/XI60/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM1 N_XI0/XI60/XI6/NET33_XI0/XI60/XI6/MM1_d
+ N_XI0/XI60/XI6/NET34_XI0/XI60/XI6/MM1_g N_VSS_XI0/XI60/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM9 N_XI0/XI60/XI6/NET36_XI0/XI60/XI6/MM9_d
+ N_WL<117>_XI0/XI60/XI6/MM9_g N_BL<9>_XI0/XI60/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM6 N_XI0/XI60/XI6/NET35_XI0/XI60/XI6/MM6_d
+ N_XI0/XI60/XI6/NET36_XI0/XI60/XI6/MM6_g N_VSS_XI0/XI60/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM7 N_XI0/XI60/XI6/NET36_XI0/XI60/XI6/MM7_d
+ N_XI0/XI60/XI6/NET35_XI0/XI60/XI6/MM7_g N_VSS_XI0/XI60/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM8 N_XI0/XI60/XI6/NET35_XI0/XI60/XI6/MM8_d
+ N_WL<117>_XI0/XI60/XI6/MM8_g N_BLN<9>_XI0/XI60/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI6/MM5 N_XI0/XI60/XI6/NET34_XI0/XI60/XI6/MM5_d
+ N_XI0/XI60/XI6/NET33_XI0/XI60/XI6/MM5_g N_VDD_XI0/XI60/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI6/MM4 N_XI0/XI60/XI6/NET33_XI0/XI60/XI6/MM4_d
+ N_XI0/XI60/XI6/NET34_XI0/XI60/XI6/MM4_g N_VDD_XI0/XI60/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI6/MM10 N_XI0/XI60/XI6/NET35_XI0/XI60/XI6/MM10_d
+ N_XI0/XI60/XI6/NET36_XI0/XI60/XI6/MM10_g N_VDD_XI0/XI60/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI6/MM11 N_XI0/XI60/XI6/NET36_XI0/XI60/XI6/MM11_d
+ N_XI0/XI60/XI6/NET35_XI0/XI60/XI6/MM11_g N_VDD_XI0/XI60/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI7/MM2 N_XI0/XI60/XI7/NET34_XI0/XI60/XI7/MM2_d
+ N_XI0/XI60/XI7/NET33_XI0/XI60/XI7/MM2_g N_VSS_XI0/XI60/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM3 N_XI0/XI60/XI7/NET33_XI0/XI60/XI7/MM3_d
+ N_WL<116>_XI0/XI60/XI7/MM3_g N_BLN<8>_XI0/XI60/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM0 N_XI0/XI60/XI7/NET34_XI0/XI60/XI7/MM0_d
+ N_WL<116>_XI0/XI60/XI7/MM0_g N_BL<8>_XI0/XI60/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM1 N_XI0/XI60/XI7/NET33_XI0/XI60/XI7/MM1_d
+ N_XI0/XI60/XI7/NET34_XI0/XI60/XI7/MM1_g N_VSS_XI0/XI60/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM9 N_XI0/XI60/XI7/NET36_XI0/XI60/XI7/MM9_d
+ N_WL<117>_XI0/XI60/XI7/MM9_g N_BL<8>_XI0/XI60/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM6 N_XI0/XI60/XI7/NET35_XI0/XI60/XI7/MM6_d
+ N_XI0/XI60/XI7/NET36_XI0/XI60/XI7/MM6_g N_VSS_XI0/XI60/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM7 N_XI0/XI60/XI7/NET36_XI0/XI60/XI7/MM7_d
+ N_XI0/XI60/XI7/NET35_XI0/XI60/XI7/MM7_g N_VSS_XI0/XI60/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM8 N_XI0/XI60/XI7/NET35_XI0/XI60/XI7/MM8_d
+ N_WL<117>_XI0/XI60/XI7/MM8_g N_BLN<8>_XI0/XI60/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI7/MM5 N_XI0/XI60/XI7/NET34_XI0/XI60/XI7/MM5_d
+ N_XI0/XI60/XI7/NET33_XI0/XI60/XI7/MM5_g N_VDD_XI0/XI60/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI7/MM4 N_XI0/XI60/XI7/NET33_XI0/XI60/XI7/MM4_d
+ N_XI0/XI60/XI7/NET34_XI0/XI60/XI7/MM4_g N_VDD_XI0/XI60/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI7/MM10 N_XI0/XI60/XI7/NET35_XI0/XI60/XI7/MM10_d
+ N_XI0/XI60/XI7/NET36_XI0/XI60/XI7/MM10_g N_VDD_XI0/XI60/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI7/MM11 N_XI0/XI60/XI7/NET36_XI0/XI60/XI7/MM11_d
+ N_XI0/XI60/XI7/NET35_XI0/XI60/XI7/MM11_g N_VDD_XI0/XI60/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI8/MM2 N_XI0/XI60/XI8/NET34_XI0/XI60/XI8/MM2_d
+ N_XI0/XI60/XI8/NET33_XI0/XI60/XI8/MM2_g N_VSS_XI0/XI60/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM3 N_XI0/XI60/XI8/NET33_XI0/XI60/XI8/MM3_d
+ N_WL<116>_XI0/XI60/XI8/MM3_g N_BLN<7>_XI0/XI60/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM0 N_XI0/XI60/XI8/NET34_XI0/XI60/XI8/MM0_d
+ N_WL<116>_XI0/XI60/XI8/MM0_g N_BL<7>_XI0/XI60/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM1 N_XI0/XI60/XI8/NET33_XI0/XI60/XI8/MM1_d
+ N_XI0/XI60/XI8/NET34_XI0/XI60/XI8/MM1_g N_VSS_XI0/XI60/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM9 N_XI0/XI60/XI8/NET36_XI0/XI60/XI8/MM9_d
+ N_WL<117>_XI0/XI60/XI8/MM9_g N_BL<7>_XI0/XI60/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM6 N_XI0/XI60/XI8/NET35_XI0/XI60/XI8/MM6_d
+ N_XI0/XI60/XI8/NET36_XI0/XI60/XI8/MM6_g N_VSS_XI0/XI60/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM7 N_XI0/XI60/XI8/NET36_XI0/XI60/XI8/MM7_d
+ N_XI0/XI60/XI8/NET35_XI0/XI60/XI8/MM7_g N_VSS_XI0/XI60/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM8 N_XI0/XI60/XI8/NET35_XI0/XI60/XI8/MM8_d
+ N_WL<117>_XI0/XI60/XI8/MM8_g N_BLN<7>_XI0/XI60/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI8/MM5 N_XI0/XI60/XI8/NET34_XI0/XI60/XI8/MM5_d
+ N_XI0/XI60/XI8/NET33_XI0/XI60/XI8/MM5_g N_VDD_XI0/XI60/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI8/MM4 N_XI0/XI60/XI8/NET33_XI0/XI60/XI8/MM4_d
+ N_XI0/XI60/XI8/NET34_XI0/XI60/XI8/MM4_g N_VDD_XI0/XI60/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI8/MM10 N_XI0/XI60/XI8/NET35_XI0/XI60/XI8/MM10_d
+ N_XI0/XI60/XI8/NET36_XI0/XI60/XI8/MM10_g N_VDD_XI0/XI60/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI8/MM11 N_XI0/XI60/XI8/NET36_XI0/XI60/XI8/MM11_d
+ N_XI0/XI60/XI8/NET35_XI0/XI60/XI8/MM11_g N_VDD_XI0/XI60/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI9/MM2 N_XI0/XI60/XI9/NET34_XI0/XI60/XI9/MM2_d
+ N_XI0/XI60/XI9/NET33_XI0/XI60/XI9/MM2_g N_VSS_XI0/XI60/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM3 N_XI0/XI60/XI9/NET33_XI0/XI60/XI9/MM3_d
+ N_WL<116>_XI0/XI60/XI9/MM3_g N_BLN<6>_XI0/XI60/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM0 N_XI0/XI60/XI9/NET34_XI0/XI60/XI9/MM0_d
+ N_WL<116>_XI0/XI60/XI9/MM0_g N_BL<6>_XI0/XI60/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM1 N_XI0/XI60/XI9/NET33_XI0/XI60/XI9/MM1_d
+ N_XI0/XI60/XI9/NET34_XI0/XI60/XI9/MM1_g N_VSS_XI0/XI60/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM9 N_XI0/XI60/XI9/NET36_XI0/XI60/XI9/MM9_d
+ N_WL<117>_XI0/XI60/XI9/MM9_g N_BL<6>_XI0/XI60/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM6 N_XI0/XI60/XI9/NET35_XI0/XI60/XI9/MM6_d
+ N_XI0/XI60/XI9/NET36_XI0/XI60/XI9/MM6_g N_VSS_XI0/XI60/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM7 N_XI0/XI60/XI9/NET36_XI0/XI60/XI9/MM7_d
+ N_XI0/XI60/XI9/NET35_XI0/XI60/XI9/MM7_g N_VSS_XI0/XI60/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM8 N_XI0/XI60/XI9/NET35_XI0/XI60/XI9/MM8_d
+ N_WL<117>_XI0/XI60/XI9/MM8_g N_BLN<6>_XI0/XI60/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI9/MM5 N_XI0/XI60/XI9/NET34_XI0/XI60/XI9/MM5_d
+ N_XI0/XI60/XI9/NET33_XI0/XI60/XI9/MM5_g N_VDD_XI0/XI60/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI9/MM4 N_XI0/XI60/XI9/NET33_XI0/XI60/XI9/MM4_d
+ N_XI0/XI60/XI9/NET34_XI0/XI60/XI9/MM4_g N_VDD_XI0/XI60/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI9/MM10 N_XI0/XI60/XI9/NET35_XI0/XI60/XI9/MM10_d
+ N_XI0/XI60/XI9/NET36_XI0/XI60/XI9/MM10_g N_VDD_XI0/XI60/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI9/MM11 N_XI0/XI60/XI9/NET36_XI0/XI60/XI9/MM11_d
+ N_XI0/XI60/XI9/NET35_XI0/XI60/XI9/MM11_g N_VDD_XI0/XI60/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI10/MM2 N_XI0/XI60/XI10/NET34_XI0/XI60/XI10/MM2_d
+ N_XI0/XI60/XI10/NET33_XI0/XI60/XI10/MM2_g N_VSS_XI0/XI60/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM3 N_XI0/XI60/XI10/NET33_XI0/XI60/XI10/MM3_d
+ N_WL<116>_XI0/XI60/XI10/MM3_g N_BLN<5>_XI0/XI60/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM0 N_XI0/XI60/XI10/NET34_XI0/XI60/XI10/MM0_d
+ N_WL<116>_XI0/XI60/XI10/MM0_g N_BL<5>_XI0/XI60/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM1 N_XI0/XI60/XI10/NET33_XI0/XI60/XI10/MM1_d
+ N_XI0/XI60/XI10/NET34_XI0/XI60/XI10/MM1_g N_VSS_XI0/XI60/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM9 N_XI0/XI60/XI10/NET36_XI0/XI60/XI10/MM9_d
+ N_WL<117>_XI0/XI60/XI10/MM9_g N_BL<5>_XI0/XI60/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM6 N_XI0/XI60/XI10/NET35_XI0/XI60/XI10/MM6_d
+ N_XI0/XI60/XI10/NET36_XI0/XI60/XI10/MM6_g N_VSS_XI0/XI60/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM7 N_XI0/XI60/XI10/NET36_XI0/XI60/XI10/MM7_d
+ N_XI0/XI60/XI10/NET35_XI0/XI60/XI10/MM7_g N_VSS_XI0/XI60/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM8 N_XI0/XI60/XI10/NET35_XI0/XI60/XI10/MM8_d
+ N_WL<117>_XI0/XI60/XI10/MM8_g N_BLN<5>_XI0/XI60/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI10/MM5 N_XI0/XI60/XI10/NET34_XI0/XI60/XI10/MM5_d
+ N_XI0/XI60/XI10/NET33_XI0/XI60/XI10/MM5_g N_VDD_XI0/XI60/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI10/MM4 N_XI0/XI60/XI10/NET33_XI0/XI60/XI10/MM4_d
+ N_XI0/XI60/XI10/NET34_XI0/XI60/XI10/MM4_g N_VDD_XI0/XI60/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI10/MM10 N_XI0/XI60/XI10/NET35_XI0/XI60/XI10/MM10_d
+ N_XI0/XI60/XI10/NET36_XI0/XI60/XI10/MM10_g N_VDD_XI0/XI60/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI10/MM11 N_XI0/XI60/XI10/NET36_XI0/XI60/XI10/MM11_d
+ N_XI0/XI60/XI10/NET35_XI0/XI60/XI10/MM11_g N_VDD_XI0/XI60/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI11/MM2 N_XI0/XI60/XI11/NET34_XI0/XI60/XI11/MM2_d
+ N_XI0/XI60/XI11/NET33_XI0/XI60/XI11/MM2_g N_VSS_XI0/XI60/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM3 N_XI0/XI60/XI11/NET33_XI0/XI60/XI11/MM3_d
+ N_WL<116>_XI0/XI60/XI11/MM3_g N_BLN<4>_XI0/XI60/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM0 N_XI0/XI60/XI11/NET34_XI0/XI60/XI11/MM0_d
+ N_WL<116>_XI0/XI60/XI11/MM0_g N_BL<4>_XI0/XI60/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM1 N_XI0/XI60/XI11/NET33_XI0/XI60/XI11/MM1_d
+ N_XI0/XI60/XI11/NET34_XI0/XI60/XI11/MM1_g N_VSS_XI0/XI60/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM9 N_XI0/XI60/XI11/NET36_XI0/XI60/XI11/MM9_d
+ N_WL<117>_XI0/XI60/XI11/MM9_g N_BL<4>_XI0/XI60/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM6 N_XI0/XI60/XI11/NET35_XI0/XI60/XI11/MM6_d
+ N_XI0/XI60/XI11/NET36_XI0/XI60/XI11/MM6_g N_VSS_XI0/XI60/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM7 N_XI0/XI60/XI11/NET36_XI0/XI60/XI11/MM7_d
+ N_XI0/XI60/XI11/NET35_XI0/XI60/XI11/MM7_g N_VSS_XI0/XI60/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM8 N_XI0/XI60/XI11/NET35_XI0/XI60/XI11/MM8_d
+ N_WL<117>_XI0/XI60/XI11/MM8_g N_BLN<4>_XI0/XI60/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI11/MM5 N_XI0/XI60/XI11/NET34_XI0/XI60/XI11/MM5_d
+ N_XI0/XI60/XI11/NET33_XI0/XI60/XI11/MM5_g N_VDD_XI0/XI60/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI11/MM4 N_XI0/XI60/XI11/NET33_XI0/XI60/XI11/MM4_d
+ N_XI0/XI60/XI11/NET34_XI0/XI60/XI11/MM4_g N_VDD_XI0/XI60/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI11/MM10 N_XI0/XI60/XI11/NET35_XI0/XI60/XI11/MM10_d
+ N_XI0/XI60/XI11/NET36_XI0/XI60/XI11/MM10_g N_VDD_XI0/XI60/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI11/MM11 N_XI0/XI60/XI11/NET36_XI0/XI60/XI11/MM11_d
+ N_XI0/XI60/XI11/NET35_XI0/XI60/XI11/MM11_g N_VDD_XI0/XI60/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI12/MM2 N_XI0/XI60/XI12/NET34_XI0/XI60/XI12/MM2_d
+ N_XI0/XI60/XI12/NET33_XI0/XI60/XI12/MM2_g N_VSS_XI0/XI60/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM3 N_XI0/XI60/XI12/NET33_XI0/XI60/XI12/MM3_d
+ N_WL<116>_XI0/XI60/XI12/MM3_g N_BLN<3>_XI0/XI60/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM0 N_XI0/XI60/XI12/NET34_XI0/XI60/XI12/MM0_d
+ N_WL<116>_XI0/XI60/XI12/MM0_g N_BL<3>_XI0/XI60/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM1 N_XI0/XI60/XI12/NET33_XI0/XI60/XI12/MM1_d
+ N_XI0/XI60/XI12/NET34_XI0/XI60/XI12/MM1_g N_VSS_XI0/XI60/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM9 N_XI0/XI60/XI12/NET36_XI0/XI60/XI12/MM9_d
+ N_WL<117>_XI0/XI60/XI12/MM9_g N_BL<3>_XI0/XI60/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM6 N_XI0/XI60/XI12/NET35_XI0/XI60/XI12/MM6_d
+ N_XI0/XI60/XI12/NET36_XI0/XI60/XI12/MM6_g N_VSS_XI0/XI60/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM7 N_XI0/XI60/XI12/NET36_XI0/XI60/XI12/MM7_d
+ N_XI0/XI60/XI12/NET35_XI0/XI60/XI12/MM7_g N_VSS_XI0/XI60/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM8 N_XI0/XI60/XI12/NET35_XI0/XI60/XI12/MM8_d
+ N_WL<117>_XI0/XI60/XI12/MM8_g N_BLN<3>_XI0/XI60/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI12/MM5 N_XI0/XI60/XI12/NET34_XI0/XI60/XI12/MM5_d
+ N_XI0/XI60/XI12/NET33_XI0/XI60/XI12/MM5_g N_VDD_XI0/XI60/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI12/MM4 N_XI0/XI60/XI12/NET33_XI0/XI60/XI12/MM4_d
+ N_XI0/XI60/XI12/NET34_XI0/XI60/XI12/MM4_g N_VDD_XI0/XI60/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI12/MM10 N_XI0/XI60/XI12/NET35_XI0/XI60/XI12/MM10_d
+ N_XI0/XI60/XI12/NET36_XI0/XI60/XI12/MM10_g N_VDD_XI0/XI60/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI12/MM11 N_XI0/XI60/XI12/NET36_XI0/XI60/XI12/MM11_d
+ N_XI0/XI60/XI12/NET35_XI0/XI60/XI12/MM11_g N_VDD_XI0/XI60/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI13/MM2 N_XI0/XI60/XI13/NET34_XI0/XI60/XI13/MM2_d
+ N_XI0/XI60/XI13/NET33_XI0/XI60/XI13/MM2_g N_VSS_XI0/XI60/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM3 N_XI0/XI60/XI13/NET33_XI0/XI60/XI13/MM3_d
+ N_WL<116>_XI0/XI60/XI13/MM3_g N_BLN<2>_XI0/XI60/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM0 N_XI0/XI60/XI13/NET34_XI0/XI60/XI13/MM0_d
+ N_WL<116>_XI0/XI60/XI13/MM0_g N_BL<2>_XI0/XI60/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM1 N_XI0/XI60/XI13/NET33_XI0/XI60/XI13/MM1_d
+ N_XI0/XI60/XI13/NET34_XI0/XI60/XI13/MM1_g N_VSS_XI0/XI60/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM9 N_XI0/XI60/XI13/NET36_XI0/XI60/XI13/MM9_d
+ N_WL<117>_XI0/XI60/XI13/MM9_g N_BL<2>_XI0/XI60/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM6 N_XI0/XI60/XI13/NET35_XI0/XI60/XI13/MM6_d
+ N_XI0/XI60/XI13/NET36_XI0/XI60/XI13/MM6_g N_VSS_XI0/XI60/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM7 N_XI0/XI60/XI13/NET36_XI0/XI60/XI13/MM7_d
+ N_XI0/XI60/XI13/NET35_XI0/XI60/XI13/MM7_g N_VSS_XI0/XI60/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM8 N_XI0/XI60/XI13/NET35_XI0/XI60/XI13/MM8_d
+ N_WL<117>_XI0/XI60/XI13/MM8_g N_BLN<2>_XI0/XI60/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI13/MM5 N_XI0/XI60/XI13/NET34_XI0/XI60/XI13/MM5_d
+ N_XI0/XI60/XI13/NET33_XI0/XI60/XI13/MM5_g N_VDD_XI0/XI60/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI13/MM4 N_XI0/XI60/XI13/NET33_XI0/XI60/XI13/MM4_d
+ N_XI0/XI60/XI13/NET34_XI0/XI60/XI13/MM4_g N_VDD_XI0/XI60/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI13/MM10 N_XI0/XI60/XI13/NET35_XI0/XI60/XI13/MM10_d
+ N_XI0/XI60/XI13/NET36_XI0/XI60/XI13/MM10_g N_VDD_XI0/XI60/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI13/MM11 N_XI0/XI60/XI13/NET36_XI0/XI60/XI13/MM11_d
+ N_XI0/XI60/XI13/NET35_XI0/XI60/XI13/MM11_g N_VDD_XI0/XI60/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI14/MM2 N_XI0/XI60/XI14/NET34_XI0/XI60/XI14/MM2_d
+ N_XI0/XI60/XI14/NET33_XI0/XI60/XI14/MM2_g N_VSS_XI0/XI60/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM3 N_XI0/XI60/XI14/NET33_XI0/XI60/XI14/MM3_d
+ N_WL<116>_XI0/XI60/XI14/MM3_g N_BLN<1>_XI0/XI60/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM0 N_XI0/XI60/XI14/NET34_XI0/XI60/XI14/MM0_d
+ N_WL<116>_XI0/XI60/XI14/MM0_g N_BL<1>_XI0/XI60/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM1 N_XI0/XI60/XI14/NET33_XI0/XI60/XI14/MM1_d
+ N_XI0/XI60/XI14/NET34_XI0/XI60/XI14/MM1_g N_VSS_XI0/XI60/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM9 N_XI0/XI60/XI14/NET36_XI0/XI60/XI14/MM9_d
+ N_WL<117>_XI0/XI60/XI14/MM9_g N_BL<1>_XI0/XI60/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM6 N_XI0/XI60/XI14/NET35_XI0/XI60/XI14/MM6_d
+ N_XI0/XI60/XI14/NET36_XI0/XI60/XI14/MM6_g N_VSS_XI0/XI60/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM7 N_XI0/XI60/XI14/NET36_XI0/XI60/XI14/MM7_d
+ N_XI0/XI60/XI14/NET35_XI0/XI60/XI14/MM7_g N_VSS_XI0/XI60/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM8 N_XI0/XI60/XI14/NET35_XI0/XI60/XI14/MM8_d
+ N_WL<117>_XI0/XI60/XI14/MM8_g N_BLN<1>_XI0/XI60/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI14/MM5 N_XI0/XI60/XI14/NET34_XI0/XI60/XI14/MM5_d
+ N_XI0/XI60/XI14/NET33_XI0/XI60/XI14/MM5_g N_VDD_XI0/XI60/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI14/MM4 N_XI0/XI60/XI14/NET33_XI0/XI60/XI14/MM4_d
+ N_XI0/XI60/XI14/NET34_XI0/XI60/XI14/MM4_g N_VDD_XI0/XI60/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI14/MM10 N_XI0/XI60/XI14/NET35_XI0/XI60/XI14/MM10_d
+ N_XI0/XI60/XI14/NET36_XI0/XI60/XI14/MM10_g N_VDD_XI0/XI60/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI14/MM11 N_XI0/XI60/XI14/NET36_XI0/XI60/XI14/MM11_d
+ N_XI0/XI60/XI14/NET35_XI0/XI60/XI14/MM11_g N_VDD_XI0/XI60/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI15/MM2 N_XI0/XI60/XI15/NET34_XI0/XI60/XI15/MM2_d
+ N_XI0/XI60/XI15/NET33_XI0/XI60/XI15/MM2_g N_VSS_XI0/XI60/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM3 N_XI0/XI60/XI15/NET33_XI0/XI60/XI15/MM3_d
+ N_WL<116>_XI0/XI60/XI15/MM3_g N_BLN<0>_XI0/XI60/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM0 N_XI0/XI60/XI15/NET34_XI0/XI60/XI15/MM0_d
+ N_WL<116>_XI0/XI60/XI15/MM0_g N_BL<0>_XI0/XI60/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM1 N_XI0/XI60/XI15/NET33_XI0/XI60/XI15/MM1_d
+ N_XI0/XI60/XI15/NET34_XI0/XI60/XI15/MM1_g N_VSS_XI0/XI60/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM9 N_XI0/XI60/XI15/NET36_XI0/XI60/XI15/MM9_d
+ N_WL<117>_XI0/XI60/XI15/MM9_g N_BL<0>_XI0/XI60/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM6 N_XI0/XI60/XI15/NET35_XI0/XI60/XI15/MM6_d
+ N_XI0/XI60/XI15/NET36_XI0/XI60/XI15/MM6_g N_VSS_XI0/XI60/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM7 N_XI0/XI60/XI15/NET36_XI0/XI60/XI15/MM7_d
+ N_XI0/XI60/XI15/NET35_XI0/XI60/XI15/MM7_g N_VSS_XI0/XI60/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM8 N_XI0/XI60/XI15/NET35_XI0/XI60/XI15/MM8_d
+ N_WL<117>_XI0/XI60/XI15/MM8_g N_BLN<0>_XI0/XI60/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI60/XI15/MM5 N_XI0/XI60/XI15/NET34_XI0/XI60/XI15/MM5_d
+ N_XI0/XI60/XI15/NET33_XI0/XI60/XI15/MM5_g N_VDD_XI0/XI60/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI15/MM4 N_XI0/XI60/XI15/NET33_XI0/XI60/XI15/MM4_d
+ N_XI0/XI60/XI15/NET34_XI0/XI60/XI15/MM4_g N_VDD_XI0/XI60/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI15/MM10 N_XI0/XI60/XI15/NET35_XI0/XI60/XI15/MM10_d
+ N_XI0/XI60/XI15/NET36_XI0/XI60/XI15/MM10_g N_VDD_XI0/XI60/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI60/XI15/MM11 N_XI0/XI60/XI15/NET36_XI0/XI60/XI15/MM11_d
+ N_XI0/XI60/XI15/NET35_XI0/XI60/XI15/MM11_g N_VDD_XI0/XI60/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI0/MM2 N_XI0/XI61/XI0/NET34_XI0/XI61/XI0/MM2_d
+ N_XI0/XI61/XI0/NET33_XI0/XI61/XI0/MM2_g N_VSS_XI0/XI61/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM3 N_XI0/XI61/XI0/NET33_XI0/XI61/XI0/MM3_d
+ N_WL<118>_XI0/XI61/XI0/MM3_g N_BLN<15>_XI0/XI61/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM0 N_XI0/XI61/XI0/NET34_XI0/XI61/XI0/MM0_d
+ N_WL<118>_XI0/XI61/XI0/MM0_g N_BL<15>_XI0/XI61/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM1 N_XI0/XI61/XI0/NET33_XI0/XI61/XI0/MM1_d
+ N_XI0/XI61/XI0/NET34_XI0/XI61/XI0/MM1_g N_VSS_XI0/XI61/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM9 N_XI0/XI61/XI0/NET36_XI0/XI61/XI0/MM9_d
+ N_WL<119>_XI0/XI61/XI0/MM9_g N_BL<15>_XI0/XI61/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM6 N_XI0/XI61/XI0/NET35_XI0/XI61/XI0/MM6_d
+ N_XI0/XI61/XI0/NET36_XI0/XI61/XI0/MM6_g N_VSS_XI0/XI61/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM7 N_XI0/XI61/XI0/NET36_XI0/XI61/XI0/MM7_d
+ N_XI0/XI61/XI0/NET35_XI0/XI61/XI0/MM7_g N_VSS_XI0/XI61/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM8 N_XI0/XI61/XI0/NET35_XI0/XI61/XI0/MM8_d
+ N_WL<119>_XI0/XI61/XI0/MM8_g N_BLN<15>_XI0/XI61/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI0/MM5 N_XI0/XI61/XI0/NET34_XI0/XI61/XI0/MM5_d
+ N_XI0/XI61/XI0/NET33_XI0/XI61/XI0/MM5_g N_VDD_XI0/XI61/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI0/MM4 N_XI0/XI61/XI0/NET33_XI0/XI61/XI0/MM4_d
+ N_XI0/XI61/XI0/NET34_XI0/XI61/XI0/MM4_g N_VDD_XI0/XI61/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI0/MM10 N_XI0/XI61/XI0/NET35_XI0/XI61/XI0/MM10_d
+ N_XI0/XI61/XI0/NET36_XI0/XI61/XI0/MM10_g N_VDD_XI0/XI61/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI0/MM11 N_XI0/XI61/XI0/NET36_XI0/XI61/XI0/MM11_d
+ N_XI0/XI61/XI0/NET35_XI0/XI61/XI0/MM11_g N_VDD_XI0/XI61/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI1/MM2 N_XI0/XI61/XI1/NET34_XI0/XI61/XI1/MM2_d
+ N_XI0/XI61/XI1/NET33_XI0/XI61/XI1/MM2_g N_VSS_XI0/XI61/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM3 N_XI0/XI61/XI1/NET33_XI0/XI61/XI1/MM3_d
+ N_WL<118>_XI0/XI61/XI1/MM3_g N_BLN<14>_XI0/XI61/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM0 N_XI0/XI61/XI1/NET34_XI0/XI61/XI1/MM0_d
+ N_WL<118>_XI0/XI61/XI1/MM0_g N_BL<14>_XI0/XI61/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM1 N_XI0/XI61/XI1/NET33_XI0/XI61/XI1/MM1_d
+ N_XI0/XI61/XI1/NET34_XI0/XI61/XI1/MM1_g N_VSS_XI0/XI61/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM9 N_XI0/XI61/XI1/NET36_XI0/XI61/XI1/MM9_d
+ N_WL<119>_XI0/XI61/XI1/MM9_g N_BL<14>_XI0/XI61/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM6 N_XI0/XI61/XI1/NET35_XI0/XI61/XI1/MM6_d
+ N_XI0/XI61/XI1/NET36_XI0/XI61/XI1/MM6_g N_VSS_XI0/XI61/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM7 N_XI0/XI61/XI1/NET36_XI0/XI61/XI1/MM7_d
+ N_XI0/XI61/XI1/NET35_XI0/XI61/XI1/MM7_g N_VSS_XI0/XI61/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM8 N_XI0/XI61/XI1/NET35_XI0/XI61/XI1/MM8_d
+ N_WL<119>_XI0/XI61/XI1/MM8_g N_BLN<14>_XI0/XI61/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI1/MM5 N_XI0/XI61/XI1/NET34_XI0/XI61/XI1/MM5_d
+ N_XI0/XI61/XI1/NET33_XI0/XI61/XI1/MM5_g N_VDD_XI0/XI61/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI1/MM4 N_XI0/XI61/XI1/NET33_XI0/XI61/XI1/MM4_d
+ N_XI0/XI61/XI1/NET34_XI0/XI61/XI1/MM4_g N_VDD_XI0/XI61/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI1/MM10 N_XI0/XI61/XI1/NET35_XI0/XI61/XI1/MM10_d
+ N_XI0/XI61/XI1/NET36_XI0/XI61/XI1/MM10_g N_VDD_XI0/XI61/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI1/MM11 N_XI0/XI61/XI1/NET36_XI0/XI61/XI1/MM11_d
+ N_XI0/XI61/XI1/NET35_XI0/XI61/XI1/MM11_g N_VDD_XI0/XI61/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI2/MM2 N_XI0/XI61/XI2/NET34_XI0/XI61/XI2/MM2_d
+ N_XI0/XI61/XI2/NET33_XI0/XI61/XI2/MM2_g N_VSS_XI0/XI61/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM3 N_XI0/XI61/XI2/NET33_XI0/XI61/XI2/MM3_d
+ N_WL<118>_XI0/XI61/XI2/MM3_g N_BLN<13>_XI0/XI61/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM0 N_XI0/XI61/XI2/NET34_XI0/XI61/XI2/MM0_d
+ N_WL<118>_XI0/XI61/XI2/MM0_g N_BL<13>_XI0/XI61/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM1 N_XI0/XI61/XI2/NET33_XI0/XI61/XI2/MM1_d
+ N_XI0/XI61/XI2/NET34_XI0/XI61/XI2/MM1_g N_VSS_XI0/XI61/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM9 N_XI0/XI61/XI2/NET36_XI0/XI61/XI2/MM9_d
+ N_WL<119>_XI0/XI61/XI2/MM9_g N_BL<13>_XI0/XI61/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM6 N_XI0/XI61/XI2/NET35_XI0/XI61/XI2/MM6_d
+ N_XI0/XI61/XI2/NET36_XI0/XI61/XI2/MM6_g N_VSS_XI0/XI61/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM7 N_XI0/XI61/XI2/NET36_XI0/XI61/XI2/MM7_d
+ N_XI0/XI61/XI2/NET35_XI0/XI61/XI2/MM7_g N_VSS_XI0/XI61/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM8 N_XI0/XI61/XI2/NET35_XI0/XI61/XI2/MM8_d
+ N_WL<119>_XI0/XI61/XI2/MM8_g N_BLN<13>_XI0/XI61/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI2/MM5 N_XI0/XI61/XI2/NET34_XI0/XI61/XI2/MM5_d
+ N_XI0/XI61/XI2/NET33_XI0/XI61/XI2/MM5_g N_VDD_XI0/XI61/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI2/MM4 N_XI0/XI61/XI2/NET33_XI0/XI61/XI2/MM4_d
+ N_XI0/XI61/XI2/NET34_XI0/XI61/XI2/MM4_g N_VDD_XI0/XI61/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI2/MM10 N_XI0/XI61/XI2/NET35_XI0/XI61/XI2/MM10_d
+ N_XI0/XI61/XI2/NET36_XI0/XI61/XI2/MM10_g N_VDD_XI0/XI61/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI2/MM11 N_XI0/XI61/XI2/NET36_XI0/XI61/XI2/MM11_d
+ N_XI0/XI61/XI2/NET35_XI0/XI61/XI2/MM11_g N_VDD_XI0/XI61/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI3/MM2 N_XI0/XI61/XI3/NET34_XI0/XI61/XI3/MM2_d
+ N_XI0/XI61/XI3/NET33_XI0/XI61/XI3/MM2_g N_VSS_XI0/XI61/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM3 N_XI0/XI61/XI3/NET33_XI0/XI61/XI3/MM3_d
+ N_WL<118>_XI0/XI61/XI3/MM3_g N_BLN<12>_XI0/XI61/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM0 N_XI0/XI61/XI3/NET34_XI0/XI61/XI3/MM0_d
+ N_WL<118>_XI0/XI61/XI3/MM0_g N_BL<12>_XI0/XI61/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM1 N_XI0/XI61/XI3/NET33_XI0/XI61/XI3/MM1_d
+ N_XI0/XI61/XI3/NET34_XI0/XI61/XI3/MM1_g N_VSS_XI0/XI61/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM9 N_XI0/XI61/XI3/NET36_XI0/XI61/XI3/MM9_d
+ N_WL<119>_XI0/XI61/XI3/MM9_g N_BL<12>_XI0/XI61/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM6 N_XI0/XI61/XI3/NET35_XI0/XI61/XI3/MM6_d
+ N_XI0/XI61/XI3/NET36_XI0/XI61/XI3/MM6_g N_VSS_XI0/XI61/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM7 N_XI0/XI61/XI3/NET36_XI0/XI61/XI3/MM7_d
+ N_XI0/XI61/XI3/NET35_XI0/XI61/XI3/MM7_g N_VSS_XI0/XI61/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM8 N_XI0/XI61/XI3/NET35_XI0/XI61/XI3/MM8_d
+ N_WL<119>_XI0/XI61/XI3/MM8_g N_BLN<12>_XI0/XI61/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI3/MM5 N_XI0/XI61/XI3/NET34_XI0/XI61/XI3/MM5_d
+ N_XI0/XI61/XI3/NET33_XI0/XI61/XI3/MM5_g N_VDD_XI0/XI61/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI3/MM4 N_XI0/XI61/XI3/NET33_XI0/XI61/XI3/MM4_d
+ N_XI0/XI61/XI3/NET34_XI0/XI61/XI3/MM4_g N_VDD_XI0/XI61/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI3/MM10 N_XI0/XI61/XI3/NET35_XI0/XI61/XI3/MM10_d
+ N_XI0/XI61/XI3/NET36_XI0/XI61/XI3/MM10_g N_VDD_XI0/XI61/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI3/MM11 N_XI0/XI61/XI3/NET36_XI0/XI61/XI3/MM11_d
+ N_XI0/XI61/XI3/NET35_XI0/XI61/XI3/MM11_g N_VDD_XI0/XI61/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI4/MM2 N_XI0/XI61/XI4/NET34_XI0/XI61/XI4/MM2_d
+ N_XI0/XI61/XI4/NET33_XI0/XI61/XI4/MM2_g N_VSS_XI0/XI61/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM3 N_XI0/XI61/XI4/NET33_XI0/XI61/XI4/MM3_d
+ N_WL<118>_XI0/XI61/XI4/MM3_g N_BLN<11>_XI0/XI61/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM0 N_XI0/XI61/XI4/NET34_XI0/XI61/XI4/MM0_d
+ N_WL<118>_XI0/XI61/XI4/MM0_g N_BL<11>_XI0/XI61/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM1 N_XI0/XI61/XI4/NET33_XI0/XI61/XI4/MM1_d
+ N_XI0/XI61/XI4/NET34_XI0/XI61/XI4/MM1_g N_VSS_XI0/XI61/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM9 N_XI0/XI61/XI4/NET36_XI0/XI61/XI4/MM9_d
+ N_WL<119>_XI0/XI61/XI4/MM9_g N_BL<11>_XI0/XI61/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM6 N_XI0/XI61/XI4/NET35_XI0/XI61/XI4/MM6_d
+ N_XI0/XI61/XI4/NET36_XI0/XI61/XI4/MM6_g N_VSS_XI0/XI61/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM7 N_XI0/XI61/XI4/NET36_XI0/XI61/XI4/MM7_d
+ N_XI0/XI61/XI4/NET35_XI0/XI61/XI4/MM7_g N_VSS_XI0/XI61/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM8 N_XI0/XI61/XI4/NET35_XI0/XI61/XI4/MM8_d
+ N_WL<119>_XI0/XI61/XI4/MM8_g N_BLN<11>_XI0/XI61/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI4/MM5 N_XI0/XI61/XI4/NET34_XI0/XI61/XI4/MM5_d
+ N_XI0/XI61/XI4/NET33_XI0/XI61/XI4/MM5_g N_VDD_XI0/XI61/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI4/MM4 N_XI0/XI61/XI4/NET33_XI0/XI61/XI4/MM4_d
+ N_XI0/XI61/XI4/NET34_XI0/XI61/XI4/MM4_g N_VDD_XI0/XI61/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI4/MM10 N_XI0/XI61/XI4/NET35_XI0/XI61/XI4/MM10_d
+ N_XI0/XI61/XI4/NET36_XI0/XI61/XI4/MM10_g N_VDD_XI0/XI61/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI4/MM11 N_XI0/XI61/XI4/NET36_XI0/XI61/XI4/MM11_d
+ N_XI0/XI61/XI4/NET35_XI0/XI61/XI4/MM11_g N_VDD_XI0/XI61/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI5/MM2 N_XI0/XI61/XI5/NET34_XI0/XI61/XI5/MM2_d
+ N_XI0/XI61/XI5/NET33_XI0/XI61/XI5/MM2_g N_VSS_XI0/XI61/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM3 N_XI0/XI61/XI5/NET33_XI0/XI61/XI5/MM3_d
+ N_WL<118>_XI0/XI61/XI5/MM3_g N_BLN<10>_XI0/XI61/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM0 N_XI0/XI61/XI5/NET34_XI0/XI61/XI5/MM0_d
+ N_WL<118>_XI0/XI61/XI5/MM0_g N_BL<10>_XI0/XI61/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM1 N_XI0/XI61/XI5/NET33_XI0/XI61/XI5/MM1_d
+ N_XI0/XI61/XI5/NET34_XI0/XI61/XI5/MM1_g N_VSS_XI0/XI61/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM9 N_XI0/XI61/XI5/NET36_XI0/XI61/XI5/MM9_d
+ N_WL<119>_XI0/XI61/XI5/MM9_g N_BL<10>_XI0/XI61/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM6 N_XI0/XI61/XI5/NET35_XI0/XI61/XI5/MM6_d
+ N_XI0/XI61/XI5/NET36_XI0/XI61/XI5/MM6_g N_VSS_XI0/XI61/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM7 N_XI0/XI61/XI5/NET36_XI0/XI61/XI5/MM7_d
+ N_XI0/XI61/XI5/NET35_XI0/XI61/XI5/MM7_g N_VSS_XI0/XI61/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM8 N_XI0/XI61/XI5/NET35_XI0/XI61/XI5/MM8_d
+ N_WL<119>_XI0/XI61/XI5/MM8_g N_BLN<10>_XI0/XI61/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI5/MM5 N_XI0/XI61/XI5/NET34_XI0/XI61/XI5/MM5_d
+ N_XI0/XI61/XI5/NET33_XI0/XI61/XI5/MM5_g N_VDD_XI0/XI61/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI5/MM4 N_XI0/XI61/XI5/NET33_XI0/XI61/XI5/MM4_d
+ N_XI0/XI61/XI5/NET34_XI0/XI61/XI5/MM4_g N_VDD_XI0/XI61/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI5/MM10 N_XI0/XI61/XI5/NET35_XI0/XI61/XI5/MM10_d
+ N_XI0/XI61/XI5/NET36_XI0/XI61/XI5/MM10_g N_VDD_XI0/XI61/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI5/MM11 N_XI0/XI61/XI5/NET36_XI0/XI61/XI5/MM11_d
+ N_XI0/XI61/XI5/NET35_XI0/XI61/XI5/MM11_g N_VDD_XI0/XI61/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI6/MM2 N_XI0/XI61/XI6/NET34_XI0/XI61/XI6/MM2_d
+ N_XI0/XI61/XI6/NET33_XI0/XI61/XI6/MM2_g N_VSS_XI0/XI61/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM3 N_XI0/XI61/XI6/NET33_XI0/XI61/XI6/MM3_d
+ N_WL<118>_XI0/XI61/XI6/MM3_g N_BLN<9>_XI0/XI61/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM0 N_XI0/XI61/XI6/NET34_XI0/XI61/XI6/MM0_d
+ N_WL<118>_XI0/XI61/XI6/MM0_g N_BL<9>_XI0/XI61/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM1 N_XI0/XI61/XI6/NET33_XI0/XI61/XI6/MM1_d
+ N_XI0/XI61/XI6/NET34_XI0/XI61/XI6/MM1_g N_VSS_XI0/XI61/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM9 N_XI0/XI61/XI6/NET36_XI0/XI61/XI6/MM9_d
+ N_WL<119>_XI0/XI61/XI6/MM9_g N_BL<9>_XI0/XI61/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM6 N_XI0/XI61/XI6/NET35_XI0/XI61/XI6/MM6_d
+ N_XI0/XI61/XI6/NET36_XI0/XI61/XI6/MM6_g N_VSS_XI0/XI61/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM7 N_XI0/XI61/XI6/NET36_XI0/XI61/XI6/MM7_d
+ N_XI0/XI61/XI6/NET35_XI0/XI61/XI6/MM7_g N_VSS_XI0/XI61/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM8 N_XI0/XI61/XI6/NET35_XI0/XI61/XI6/MM8_d
+ N_WL<119>_XI0/XI61/XI6/MM8_g N_BLN<9>_XI0/XI61/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI6/MM5 N_XI0/XI61/XI6/NET34_XI0/XI61/XI6/MM5_d
+ N_XI0/XI61/XI6/NET33_XI0/XI61/XI6/MM5_g N_VDD_XI0/XI61/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI6/MM4 N_XI0/XI61/XI6/NET33_XI0/XI61/XI6/MM4_d
+ N_XI0/XI61/XI6/NET34_XI0/XI61/XI6/MM4_g N_VDD_XI0/XI61/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI6/MM10 N_XI0/XI61/XI6/NET35_XI0/XI61/XI6/MM10_d
+ N_XI0/XI61/XI6/NET36_XI0/XI61/XI6/MM10_g N_VDD_XI0/XI61/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI6/MM11 N_XI0/XI61/XI6/NET36_XI0/XI61/XI6/MM11_d
+ N_XI0/XI61/XI6/NET35_XI0/XI61/XI6/MM11_g N_VDD_XI0/XI61/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI7/MM2 N_XI0/XI61/XI7/NET34_XI0/XI61/XI7/MM2_d
+ N_XI0/XI61/XI7/NET33_XI0/XI61/XI7/MM2_g N_VSS_XI0/XI61/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM3 N_XI0/XI61/XI7/NET33_XI0/XI61/XI7/MM3_d
+ N_WL<118>_XI0/XI61/XI7/MM3_g N_BLN<8>_XI0/XI61/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM0 N_XI0/XI61/XI7/NET34_XI0/XI61/XI7/MM0_d
+ N_WL<118>_XI0/XI61/XI7/MM0_g N_BL<8>_XI0/XI61/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM1 N_XI0/XI61/XI7/NET33_XI0/XI61/XI7/MM1_d
+ N_XI0/XI61/XI7/NET34_XI0/XI61/XI7/MM1_g N_VSS_XI0/XI61/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM9 N_XI0/XI61/XI7/NET36_XI0/XI61/XI7/MM9_d
+ N_WL<119>_XI0/XI61/XI7/MM9_g N_BL<8>_XI0/XI61/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM6 N_XI0/XI61/XI7/NET35_XI0/XI61/XI7/MM6_d
+ N_XI0/XI61/XI7/NET36_XI0/XI61/XI7/MM6_g N_VSS_XI0/XI61/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM7 N_XI0/XI61/XI7/NET36_XI0/XI61/XI7/MM7_d
+ N_XI0/XI61/XI7/NET35_XI0/XI61/XI7/MM7_g N_VSS_XI0/XI61/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM8 N_XI0/XI61/XI7/NET35_XI0/XI61/XI7/MM8_d
+ N_WL<119>_XI0/XI61/XI7/MM8_g N_BLN<8>_XI0/XI61/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI7/MM5 N_XI0/XI61/XI7/NET34_XI0/XI61/XI7/MM5_d
+ N_XI0/XI61/XI7/NET33_XI0/XI61/XI7/MM5_g N_VDD_XI0/XI61/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI7/MM4 N_XI0/XI61/XI7/NET33_XI0/XI61/XI7/MM4_d
+ N_XI0/XI61/XI7/NET34_XI0/XI61/XI7/MM4_g N_VDD_XI0/XI61/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI7/MM10 N_XI0/XI61/XI7/NET35_XI0/XI61/XI7/MM10_d
+ N_XI0/XI61/XI7/NET36_XI0/XI61/XI7/MM10_g N_VDD_XI0/XI61/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI7/MM11 N_XI0/XI61/XI7/NET36_XI0/XI61/XI7/MM11_d
+ N_XI0/XI61/XI7/NET35_XI0/XI61/XI7/MM11_g N_VDD_XI0/XI61/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI8/MM2 N_XI0/XI61/XI8/NET34_XI0/XI61/XI8/MM2_d
+ N_XI0/XI61/XI8/NET33_XI0/XI61/XI8/MM2_g N_VSS_XI0/XI61/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM3 N_XI0/XI61/XI8/NET33_XI0/XI61/XI8/MM3_d
+ N_WL<118>_XI0/XI61/XI8/MM3_g N_BLN<7>_XI0/XI61/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM0 N_XI0/XI61/XI8/NET34_XI0/XI61/XI8/MM0_d
+ N_WL<118>_XI0/XI61/XI8/MM0_g N_BL<7>_XI0/XI61/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM1 N_XI0/XI61/XI8/NET33_XI0/XI61/XI8/MM1_d
+ N_XI0/XI61/XI8/NET34_XI0/XI61/XI8/MM1_g N_VSS_XI0/XI61/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM9 N_XI0/XI61/XI8/NET36_XI0/XI61/XI8/MM9_d
+ N_WL<119>_XI0/XI61/XI8/MM9_g N_BL<7>_XI0/XI61/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM6 N_XI0/XI61/XI8/NET35_XI0/XI61/XI8/MM6_d
+ N_XI0/XI61/XI8/NET36_XI0/XI61/XI8/MM6_g N_VSS_XI0/XI61/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM7 N_XI0/XI61/XI8/NET36_XI0/XI61/XI8/MM7_d
+ N_XI0/XI61/XI8/NET35_XI0/XI61/XI8/MM7_g N_VSS_XI0/XI61/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM8 N_XI0/XI61/XI8/NET35_XI0/XI61/XI8/MM8_d
+ N_WL<119>_XI0/XI61/XI8/MM8_g N_BLN<7>_XI0/XI61/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI8/MM5 N_XI0/XI61/XI8/NET34_XI0/XI61/XI8/MM5_d
+ N_XI0/XI61/XI8/NET33_XI0/XI61/XI8/MM5_g N_VDD_XI0/XI61/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI8/MM4 N_XI0/XI61/XI8/NET33_XI0/XI61/XI8/MM4_d
+ N_XI0/XI61/XI8/NET34_XI0/XI61/XI8/MM4_g N_VDD_XI0/XI61/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI8/MM10 N_XI0/XI61/XI8/NET35_XI0/XI61/XI8/MM10_d
+ N_XI0/XI61/XI8/NET36_XI0/XI61/XI8/MM10_g N_VDD_XI0/XI61/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI8/MM11 N_XI0/XI61/XI8/NET36_XI0/XI61/XI8/MM11_d
+ N_XI0/XI61/XI8/NET35_XI0/XI61/XI8/MM11_g N_VDD_XI0/XI61/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI9/MM2 N_XI0/XI61/XI9/NET34_XI0/XI61/XI9/MM2_d
+ N_XI0/XI61/XI9/NET33_XI0/XI61/XI9/MM2_g N_VSS_XI0/XI61/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM3 N_XI0/XI61/XI9/NET33_XI0/XI61/XI9/MM3_d
+ N_WL<118>_XI0/XI61/XI9/MM3_g N_BLN<6>_XI0/XI61/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM0 N_XI0/XI61/XI9/NET34_XI0/XI61/XI9/MM0_d
+ N_WL<118>_XI0/XI61/XI9/MM0_g N_BL<6>_XI0/XI61/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM1 N_XI0/XI61/XI9/NET33_XI0/XI61/XI9/MM1_d
+ N_XI0/XI61/XI9/NET34_XI0/XI61/XI9/MM1_g N_VSS_XI0/XI61/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM9 N_XI0/XI61/XI9/NET36_XI0/XI61/XI9/MM9_d
+ N_WL<119>_XI0/XI61/XI9/MM9_g N_BL<6>_XI0/XI61/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM6 N_XI0/XI61/XI9/NET35_XI0/XI61/XI9/MM6_d
+ N_XI0/XI61/XI9/NET36_XI0/XI61/XI9/MM6_g N_VSS_XI0/XI61/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM7 N_XI0/XI61/XI9/NET36_XI0/XI61/XI9/MM7_d
+ N_XI0/XI61/XI9/NET35_XI0/XI61/XI9/MM7_g N_VSS_XI0/XI61/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM8 N_XI0/XI61/XI9/NET35_XI0/XI61/XI9/MM8_d
+ N_WL<119>_XI0/XI61/XI9/MM8_g N_BLN<6>_XI0/XI61/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI9/MM5 N_XI0/XI61/XI9/NET34_XI0/XI61/XI9/MM5_d
+ N_XI0/XI61/XI9/NET33_XI0/XI61/XI9/MM5_g N_VDD_XI0/XI61/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI9/MM4 N_XI0/XI61/XI9/NET33_XI0/XI61/XI9/MM4_d
+ N_XI0/XI61/XI9/NET34_XI0/XI61/XI9/MM4_g N_VDD_XI0/XI61/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI9/MM10 N_XI0/XI61/XI9/NET35_XI0/XI61/XI9/MM10_d
+ N_XI0/XI61/XI9/NET36_XI0/XI61/XI9/MM10_g N_VDD_XI0/XI61/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI9/MM11 N_XI0/XI61/XI9/NET36_XI0/XI61/XI9/MM11_d
+ N_XI0/XI61/XI9/NET35_XI0/XI61/XI9/MM11_g N_VDD_XI0/XI61/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI10/MM2 N_XI0/XI61/XI10/NET34_XI0/XI61/XI10/MM2_d
+ N_XI0/XI61/XI10/NET33_XI0/XI61/XI10/MM2_g N_VSS_XI0/XI61/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM3 N_XI0/XI61/XI10/NET33_XI0/XI61/XI10/MM3_d
+ N_WL<118>_XI0/XI61/XI10/MM3_g N_BLN<5>_XI0/XI61/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM0 N_XI0/XI61/XI10/NET34_XI0/XI61/XI10/MM0_d
+ N_WL<118>_XI0/XI61/XI10/MM0_g N_BL<5>_XI0/XI61/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM1 N_XI0/XI61/XI10/NET33_XI0/XI61/XI10/MM1_d
+ N_XI0/XI61/XI10/NET34_XI0/XI61/XI10/MM1_g N_VSS_XI0/XI61/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM9 N_XI0/XI61/XI10/NET36_XI0/XI61/XI10/MM9_d
+ N_WL<119>_XI0/XI61/XI10/MM9_g N_BL<5>_XI0/XI61/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM6 N_XI0/XI61/XI10/NET35_XI0/XI61/XI10/MM6_d
+ N_XI0/XI61/XI10/NET36_XI0/XI61/XI10/MM6_g N_VSS_XI0/XI61/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM7 N_XI0/XI61/XI10/NET36_XI0/XI61/XI10/MM7_d
+ N_XI0/XI61/XI10/NET35_XI0/XI61/XI10/MM7_g N_VSS_XI0/XI61/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM8 N_XI0/XI61/XI10/NET35_XI0/XI61/XI10/MM8_d
+ N_WL<119>_XI0/XI61/XI10/MM8_g N_BLN<5>_XI0/XI61/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI10/MM5 N_XI0/XI61/XI10/NET34_XI0/XI61/XI10/MM5_d
+ N_XI0/XI61/XI10/NET33_XI0/XI61/XI10/MM5_g N_VDD_XI0/XI61/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI10/MM4 N_XI0/XI61/XI10/NET33_XI0/XI61/XI10/MM4_d
+ N_XI0/XI61/XI10/NET34_XI0/XI61/XI10/MM4_g N_VDD_XI0/XI61/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI10/MM10 N_XI0/XI61/XI10/NET35_XI0/XI61/XI10/MM10_d
+ N_XI0/XI61/XI10/NET36_XI0/XI61/XI10/MM10_g N_VDD_XI0/XI61/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI10/MM11 N_XI0/XI61/XI10/NET36_XI0/XI61/XI10/MM11_d
+ N_XI0/XI61/XI10/NET35_XI0/XI61/XI10/MM11_g N_VDD_XI0/XI61/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI11/MM2 N_XI0/XI61/XI11/NET34_XI0/XI61/XI11/MM2_d
+ N_XI0/XI61/XI11/NET33_XI0/XI61/XI11/MM2_g N_VSS_XI0/XI61/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM3 N_XI0/XI61/XI11/NET33_XI0/XI61/XI11/MM3_d
+ N_WL<118>_XI0/XI61/XI11/MM3_g N_BLN<4>_XI0/XI61/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM0 N_XI0/XI61/XI11/NET34_XI0/XI61/XI11/MM0_d
+ N_WL<118>_XI0/XI61/XI11/MM0_g N_BL<4>_XI0/XI61/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM1 N_XI0/XI61/XI11/NET33_XI0/XI61/XI11/MM1_d
+ N_XI0/XI61/XI11/NET34_XI0/XI61/XI11/MM1_g N_VSS_XI0/XI61/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM9 N_XI0/XI61/XI11/NET36_XI0/XI61/XI11/MM9_d
+ N_WL<119>_XI0/XI61/XI11/MM9_g N_BL<4>_XI0/XI61/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM6 N_XI0/XI61/XI11/NET35_XI0/XI61/XI11/MM6_d
+ N_XI0/XI61/XI11/NET36_XI0/XI61/XI11/MM6_g N_VSS_XI0/XI61/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM7 N_XI0/XI61/XI11/NET36_XI0/XI61/XI11/MM7_d
+ N_XI0/XI61/XI11/NET35_XI0/XI61/XI11/MM7_g N_VSS_XI0/XI61/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM8 N_XI0/XI61/XI11/NET35_XI0/XI61/XI11/MM8_d
+ N_WL<119>_XI0/XI61/XI11/MM8_g N_BLN<4>_XI0/XI61/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI11/MM5 N_XI0/XI61/XI11/NET34_XI0/XI61/XI11/MM5_d
+ N_XI0/XI61/XI11/NET33_XI0/XI61/XI11/MM5_g N_VDD_XI0/XI61/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI11/MM4 N_XI0/XI61/XI11/NET33_XI0/XI61/XI11/MM4_d
+ N_XI0/XI61/XI11/NET34_XI0/XI61/XI11/MM4_g N_VDD_XI0/XI61/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI11/MM10 N_XI0/XI61/XI11/NET35_XI0/XI61/XI11/MM10_d
+ N_XI0/XI61/XI11/NET36_XI0/XI61/XI11/MM10_g N_VDD_XI0/XI61/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI11/MM11 N_XI0/XI61/XI11/NET36_XI0/XI61/XI11/MM11_d
+ N_XI0/XI61/XI11/NET35_XI0/XI61/XI11/MM11_g N_VDD_XI0/XI61/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI12/MM2 N_XI0/XI61/XI12/NET34_XI0/XI61/XI12/MM2_d
+ N_XI0/XI61/XI12/NET33_XI0/XI61/XI12/MM2_g N_VSS_XI0/XI61/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM3 N_XI0/XI61/XI12/NET33_XI0/XI61/XI12/MM3_d
+ N_WL<118>_XI0/XI61/XI12/MM3_g N_BLN<3>_XI0/XI61/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM0 N_XI0/XI61/XI12/NET34_XI0/XI61/XI12/MM0_d
+ N_WL<118>_XI0/XI61/XI12/MM0_g N_BL<3>_XI0/XI61/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM1 N_XI0/XI61/XI12/NET33_XI0/XI61/XI12/MM1_d
+ N_XI0/XI61/XI12/NET34_XI0/XI61/XI12/MM1_g N_VSS_XI0/XI61/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM9 N_XI0/XI61/XI12/NET36_XI0/XI61/XI12/MM9_d
+ N_WL<119>_XI0/XI61/XI12/MM9_g N_BL<3>_XI0/XI61/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM6 N_XI0/XI61/XI12/NET35_XI0/XI61/XI12/MM6_d
+ N_XI0/XI61/XI12/NET36_XI0/XI61/XI12/MM6_g N_VSS_XI0/XI61/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM7 N_XI0/XI61/XI12/NET36_XI0/XI61/XI12/MM7_d
+ N_XI0/XI61/XI12/NET35_XI0/XI61/XI12/MM7_g N_VSS_XI0/XI61/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM8 N_XI0/XI61/XI12/NET35_XI0/XI61/XI12/MM8_d
+ N_WL<119>_XI0/XI61/XI12/MM8_g N_BLN<3>_XI0/XI61/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI12/MM5 N_XI0/XI61/XI12/NET34_XI0/XI61/XI12/MM5_d
+ N_XI0/XI61/XI12/NET33_XI0/XI61/XI12/MM5_g N_VDD_XI0/XI61/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI12/MM4 N_XI0/XI61/XI12/NET33_XI0/XI61/XI12/MM4_d
+ N_XI0/XI61/XI12/NET34_XI0/XI61/XI12/MM4_g N_VDD_XI0/XI61/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI12/MM10 N_XI0/XI61/XI12/NET35_XI0/XI61/XI12/MM10_d
+ N_XI0/XI61/XI12/NET36_XI0/XI61/XI12/MM10_g N_VDD_XI0/XI61/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI12/MM11 N_XI0/XI61/XI12/NET36_XI0/XI61/XI12/MM11_d
+ N_XI0/XI61/XI12/NET35_XI0/XI61/XI12/MM11_g N_VDD_XI0/XI61/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI13/MM2 N_XI0/XI61/XI13/NET34_XI0/XI61/XI13/MM2_d
+ N_XI0/XI61/XI13/NET33_XI0/XI61/XI13/MM2_g N_VSS_XI0/XI61/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM3 N_XI0/XI61/XI13/NET33_XI0/XI61/XI13/MM3_d
+ N_WL<118>_XI0/XI61/XI13/MM3_g N_BLN<2>_XI0/XI61/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM0 N_XI0/XI61/XI13/NET34_XI0/XI61/XI13/MM0_d
+ N_WL<118>_XI0/XI61/XI13/MM0_g N_BL<2>_XI0/XI61/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM1 N_XI0/XI61/XI13/NET33_XI0/XI61/XI13/MM1_d
+ N_XI0/XI61/XI13/NET34_XI0/XI61/XI13/MM1_g N_VSS_XI0/XI61/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM9 N_XI0/XI61/XI13/NET36_XI0/XI61/XI13/MM9_d
+ N_WL<119>_XI0/XI61/XI13/MM9_g N_BL<2>_XI0/XI61/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM6 N_XI0/XI61/XI13/NET35_XI0/XI61/XI13/MM6_d
+ N_XI0/XI61/XI13/NET36_XI0/XI61/XI13/MM6_g N_VSS_XI0/XI61/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM7 N_XI0/XI61/XI13/NET36_XI0/XI61/XI13/MM7_d
+ N_XI0/XI61/XI13/NET35_XI0/XI61/XI13/MM7_g N_VSS_XI0/XI61/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM8 N_XI0/XI61/XI13/NET35_XI0/XI61/XI13/MM8_d
+ N_WL<119>_XI0/XI61/XI13/MM8_g N_BLN<2>_XI0/XI61/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI13/MM5 N_XI0/XI61/XI13/NET34_XI0/XI61/XI13/MM5_d
+ N_XI0/XI61/XI13/NET33_XI0/XI61/XI13/MM5_g N_VDD_XI0/XI61/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI13/MM4 N_XI0/XI61/XI13/NET33_XI0/XI61/XI13/MM4_d
+ N_XI0/XI61/XI13/NET34_XI0/XI61/XI13/MM4_g N_VDD_XI0/XI61/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI13/MM10 N_XI0/XI61/XI13/NET35_XI0/XI61/XI13/MM10_d
+ N_XI0/XI61/XI13/NET36_XI0/XI61/XI13/MM10_g N_VDD_XI0/XI61/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI13/MM11 N_XI0/XI61/XI13/NET36_XI0/XI61/XI13/MM11_d
+ N_XI0/XI61/XI13/NET35_XI0/XI61/XI13/MM11_g N_VDD_XI0/XI61/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI14/MM2 N_XI0/XI61/XI14/NET34_XI0/XI61/XI14/MM2_d
+ N_XI0/XI61/XI14/NET33_XI0/XI61/XI14/MM2_g N_VSS_XI0/XI61/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM3 N_XI0/XI61/XI14/NET33_XI0/XI61/XI14/MM3_d
+ N_WL<118>_XI0/XI61/XI14/MM3_g N_BLN<1>_XI0/XI61/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM0 N_XI0/XI61/XI14/NET34_XI0/XI61/XI14/MM0_d
+ N_WL<118>_XI0/XI61/XI14/MM0_g N_BL<1>_XI0/XI61/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM1 N_XI0/XI61/XI14/NET33_XI0/XI61/XI14/MM1_d
+ N_XI0/XI61/XI14/NET34_XI0/XI61/XI14/MM1_g N_VSS_XI0/XI61/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM9 N_XI0/XI61/XI14/NET36_XI0/XI61/XI14/MM9_d
+ N_WL<119>_XI0/XI61/XI14/MM9_g N_BL<1>_XI0/XI61/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM6 N_XI0/XI61/XI14/NET35_XI0/XI61/XI14/MM6_d
+ N_XI0/XI61/XI14/NET36_XI0/XI61/XI14/MM6_g N_VSS_XI0/XI61/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM7 N_XI0/XI61/XI14/NET36_XI0/XI61/XI14/MM7_d
+ N_XI0/XI61/XI14/NET35_XI0/XI61/XI14/MM7_g N_VSS_XI0/XI61/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM8 N_XI0/XI61/XI14/NET35_XI0/XI61/XI14/MM8_d
+ N_WL<119>_XI0/XI61/XI14/MM8_g N_BLN<1>_XI0/XI61/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI14/MM5 N_XI0/XI61/XI14/NET34_XI0/XI61/XI14/MM5_d
+ N_XI0/XI61/XI14/NET33_XI0/XI61/XI14/MM5_g N_VDD_XI0/XI61/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI14/MM4 N_XI0/XI61/XI14/NET33_XI0/XI61/XI14/MM4_d
+ N_XI0/XI61/XI14/NET34_XI0/XI61/XI14/MM4_g N_VDD_XI0/XI61/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI14/MM10 N_XI0/XI61/XI14/NET35_XI0/XI61/XI14/MM10_d
+ N_XI0/XI61/XI14/NET36_XI0/XI61/XI14/MM10_g N_VDD_XI0/XI61/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI14/MM11 N_XI0/XI61/XI14/NET36_XI0/XI61/XI14/MM11_d
+ N_XI0/XI61/XI14/NET35_XI0/XI61/XI14/MM11_g N_VDD_XI0/XI61/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI15/MM2 N_XI0/XI61/XI15/NET34_XI0/XI61/XI15/MM2_d
+ N_XI0/XI61/XI15/NET33_XI0/XI61/XI15/MM2_g N_VSS_XI0/XI61/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM3 N_XI0/XI61/XI15/NET33_XI0/XI61/XI15/MM3_d
+ N_WL<118>_XI0/XI61/XI15/MM3_g N_BLN<0>_XI0/XI61/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM0 N_XI0/XI61/XI15/NET34_XI0/XI61/XI15/MM0_d
+ N_WL<118>_XI0/XI61/XI15/MM0_g N_BL<0>_XI0/XI61/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM1 N_XI0/XI61/XI15/NET33_XI0/XI61/XI15/MM1_d
+ N_XI0/XI61/XI15/NET34_XI0/XI61/XI15/MM1_g N_VSS_XI0/XI61/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM9 N_XI0/XI61/XI15/NET36_XI0/XI61/XI15/MM9_d
+ N_WL<119>_XI0/XI61/XI15/MM9_g N_BL<0>_XI0/XI61/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM6 N_XI0/XI61/XI15/NET35_XI0/XI61/XI15/MM6_d
+ N_XI0/XI61/XI15/NET36_XI0/XI61/XI15/MM6_g N_VSS_XI0/XI61/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM7 N_XI0/XI61/XI15/NET36_XI0/XI61/XI15/MM7_d
+ N_XI0/XI61/XI15/NET35_XI0/XI61/XI15/MM7_g N_VSS_XI0/XI61/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM8 N_XI0/XI61/XI15/NET35_XI0/XI61/XI15/MM8_d
+ N_WL<119>_XI0/XI61/XI15/MM8_g N_BLN<0>_XI0/XI61/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI61/XI15/MM5 N_XI0/XI61/XI15/NET34_XI0/XI61/XI15/MM5_d
+ N_XI0/XI61/XI15/NET33_XI0/XI61/XI15/MM5_g N_VDD_XI0/XI61/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI15/MM4 N_XI0/XI61/XI15/NET33_XI0/XI61/XI15/MM4_d
+ N_XI0/XI61/XI15/NET34_XI0/XI61/XI15/MM4_g N_VDD_XI0/XI61/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI15/MM10 N_XI0/XI61/XI15/NET35_XI0/XI61/XI15/MM10_d
+ N_XI0/XI61/XI15/NET36_XI0/XI61/XI15/MM10_g N_VDD_XI0/XI61/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI61/XI15/MM11 N_XI0/XI61/XI15/NET36_XI0/XI61/XI15/MM11_d
+ N_XI0/XI61/XI15/NET35_XI0/XI61/XI15/MM11_g N_VDD_XI0/XI61/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI0/MM2 N_XI0/XI62/XI0/NET34_XI0/XI62/XI0/MM2_d
+ N_XI0/XI62/XI0/NET33_XI0/XI62/XI0/MM2_g N_VSS_XI0/XI62/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM3 N_XI0/XI62/XI0/NET33_XI0/XI62/XI0/MM3_d
+ N_WL<120>_XI0/XI62/XI0/MM3_g N_BLN<15>_XI0/XI62/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM0 N_XI0/XI62/XI0/NET34_XI0/XI62/XI0/MM0_d
+ N_WL<120>_XI0/XI62/XI0/MM0_g N_BL<15>_XI0/XI62/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM1 N_XI0/XI62/XI0/NET33_XI0/XI62/XI0/MM1_d
+ N_XI0/XI62/XI0/NET34_XI0/XI62/XI0/MM1_g N_VSS_XI0/XI62/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM9 N_XI0/XI62/XI0/NET36_XI0/XI62/XI0/MM9_d
+ N_WL<121>_XI0/XI62/XI0/MM9_g N_BL<15>_XI0/XI62/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM6 N_XI0/XI62/XI0/NET35_XI0/XI62/XI0/MM6_d
+ N_XI0/XI62/XI0/NET36_XI0/XI62/XI0/MM6_g N_VSS_XI0/XI62/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM7 N_XI0/XI62/XI0/NET36_XI0/XI62/XI0/MM7_d
+ N_XI0/XI62/XI0/NET35_XI0/XI62/XI0/MM7_g N_VSS_XI0/XI62/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM8 N_XI0/XI62/XI0/NET35_XI0/XI62/XI0/MM8_d
+ N_WL<121>_XI0/XI62/XI0/MM8_g N_BLN<15>_XI0/XI62/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI0/MM5 N_XI0/XI62/XI0/NET34_XI0/XI62/XI0/MM5_d
+ N_XI0/XI62/XI0/NET33_XI0/XI62/XI0/MM5_g N_VDD_XI0/XI62/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI0/MM4 N_XI0/XI62/XI0/NET33_XI0/XI62/XI0/MM4_d
+ N_XI0/XI62/XI0/NET34_XI0/XI62/XI0/MM4_g N_VDD_XI0/XI62/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI0/MM10 N_XI0/XI62/XI0/NET35_XI0/XI62/XI0/MM10_d
+ N_XI0/XI62/XI0/NET36_XI0/XI62/XI0/MM10_g N_VDD_XI0/XI62/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI0/MM11 N_XI0/XI62/XI0/NET36_XI0/XI62/XI0/MM11_d
+ N_XI0/XI62/XI0/NET35_XI0/XI62/XI0/MM11_g N_VDD_XI0/XI62/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI1/MM2 N_XI0/XI62/XI1/NET34_XI0/XI62/XI1/MM2_d
+ N_XI0/XI62/XI1/NET33_XI0/XI62/XI1/MM2_g N_VSS_XI0/XI62/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM3 N_XI0/XI62/XI1/NET33_XI0/XI62/XI1/MM3_d
+ N_WL<120>_XI0/XI62/XI1/MM3_g N_BLN<14>_XI0/XI62/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM0 N_XI0/XI62/XI1/NET34_XI0/XI62/XI1/MM0_d
+ N_WL<120>_XI0/XI62/XI1/MM0_g N_BL<14>_XI0/XI62/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM1 N_XI0/XI62/XI1/NET33_XI0/XI62/XI1/MM1_d
+ N_XI0/XI62/XI1/NET34_XI0/XI62/XI1/MM1_g N_VSS_XI0/XI62/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM9 N_XI0/XI62/XI1/NET36_XI0/XI62/XI1/MM9_d
+ N_WL<121>_XI0/XI62/XI1/MM9_g N_BL<14>_XI0/XI62/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM6 N_XI0/XI62/XI1/NET35_XI0/XI62/XI1/MM6_d
+ N_XI0/XI62/XI1/NET36_XI0/XI62/XI1/MM6_g N_VSS_XI0/XI62/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM7 N_XI0/XI62/XI1/NET36_XI0/XI62/XI1/MM7_d
+ N_XI0/XI62/XI1/NET35_XI0/XI62/XI1/MM7_g N_VSS_XI0/XI62/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM8 N_XI0/XI62/XI1/NET35_XI0/XI62/XI1/MM8_d
+ N_WL<121>_XI0/XI62/XI1/MM8_g N_BLN<14>_XI0/XI62/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI1/MM5 N_XI0/XI62/XI1/NET34_XI0/XI62/XI1/MM5_d
+ N_XI0/XI62/XI1/NET33_XI0/XI62/XI1/MM5_g N_VDD_XI0/XI62/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI1/MM4 N_XI0/XI62/XI1/NET33_XI0/XI62/XI1/MM4_d
+ N_XI0/XI62/XI1/NET34_XI0/XI62/XI1/MM4_g N_VDD_XI0/XI62/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI1/MM10 N_XI0/XI62/XI1/NET35_XI0/XI62/XI1/MM10_d
+ N_XI0/XI62/XI1/NET36_XI0/XI62/XI1/MM10_g N_VDD_XI0/XI62/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI1/MM11 N_XI0/XI62/XI1/NET36_XI0/XI62/XI1/MM11_d
+ N_XI0/XI62/XI1/NET35_XI0/XI62/XI1/MM11_g N_VDD_XI0/XI62/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI2/MM2 N_XI0/XI62/XI2/NET34_XI0/XI62/XI2/MM2_d
+ N_XI0/XI62/XI2/NET33_XI0/XI62/XI2/MM2_g N_VSS_XI0/XI62/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM3 N_XI0/XI62/XI2/NET33_XI0/XI62/XI2/MM3_d
+ N_WL<120>_XI0/XI62/XI2/MM3_g N_BLN<13>_XI0/XI62/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM0 N_XI0/XI62/XI2/NET34_XI0/XI62/XI2/MM0_d
+ N_WL<120>_XI0/XI62/XI2/MM0_g N_BL<13>_XI0/XI62/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM1 N_XI0/XI62/XI2/NET33_XI0/XI62/XI2/MM1_d
+ N_XI0/XI62/XI2/NET34_XI0/XI62/XI2/MM1_g N_VSS_XI0/XI62/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM9 N_XI0/XI62/XI2/NET36_XI0/XI62/XI2/MM9_d
+ N_WL<121>_XI0/XI62/XI2/MM9_g N_BL<13>_XI0/XI62/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM6 N_XI0/XI62/XI2/NET35_XI0/XI62/XI2/MM6_d
+ N_XI0/XI62/XI2/NET36_XI0/XI62/XI2/MM6_g N_VSS_XI0/XI62/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM7 N_XI0/XI62/XI2/NET36_XI0/XI62/XI2/MM7_d
+ N_XI0/XI62/XI2/NET35_XI0/XI62/XI2/MM7_g N_VSS_XI0/XI62/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM8 N_XI0/XI62/XI2/NET35_XI0/XI62/XI2/MM8_d
+ N_WL<121>_XI0/XI62/XI2/MM8_g N_BLN<13>_XI0/XI62/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI2/MM5 N_XI0/XI62/XI2/NET34_XI0/XI62/XI2/MM5_d
+ N_XI0/XI62/XI2/NET33_XI0/XI62/XI2/MM5_g N_VDD_XI0/XI62/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI2/MM4 N_XI0/XI62/XI2/NET33_XI0/XI62/XI2/MM4_d
+ N_XI0/XI62/XI2/NET34_XI0/XI62/XI2/MM4_g N_VDD_XI0/XI62/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI2/MM10 N_XI0/XI62/XI2/NET35_XI0/XI62/XI2/MM10_d
+ N_XI0/XI62/XI2/NET36_XI0/XI62/XI2/MM10_g N_VDD_XI0/XI62/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI2/MM11 N_XI0/XI62/XI2/NET36_XI0/XI62/XI2/MM11_d
+ N_XI0/XI62/XI2/NET35_XI0/XI62/XI2/MM11_g N_VDD_XI0/XI62/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI3/MM2 N_XI0/XI62/XI3/NET34_XI0/XI62/XI3/MM2_d
+ N_XI0/XI62/XI3/NET33_XI0/XI62/XI3/MM2_g N_VSS_XI0/XI62/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM3 N_XI0/XI62/XI3/NET33_XI0/XI62/XI3/MM3_d
+ N_WL<120>_XI0/XI62/XI3/MM3_g N_BLN<12>_XI0/XI62/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM0 N_XI0/XI62/XI3/NET34_XI0/XI62/XI3/MM0_d
+ N_WL<120>_XI0/XI62/XI3/MM0_g N_BL<12>_XI0/XI62/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM1 N_XI0/XI62/XI3/NET33_XI0/XI62/XI3/MM1_d
+ N_XI0/XI62/XI3/NET34_XI0/XI62/XI3/MM1_g N_VSS_XI0/XI62/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM9 N_XI0/XI62/XI3/NET36_XI0/XI62/XI3/MM9_d
+ N_WL<121>_XI0/XI62/XI3/MM9_g N_BL<12>_XI0/XI62/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM6 N_XI0/XI62/XI3/NET35_XI0/XI62/XI3/MM6_d
+ N_XI0/XI62/XI3/NET36_XI0/XI62/XI3/MM6_g N_VSS_XI0/XI62/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM7 N_XI0/XI62/XI3/NET36_XI0/XI62/XI3/MM7_d
+ N_XI0/XI62/XI3/NET35_XI0/XI62/XI3/MM7_g N_VSS_XI0/XI62/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM8 N_XI0/XI62/XI3/NET35_XI0/XI62/XI3/MM8_d
+ N_WL<121>_XI0/XI62/XI3/MM8_g N_BLN<12>_XI0/XI62/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI3/MM5 N_XI0/XI62/XI3/NET34_XI0/XI62/XI3/MM5_d
+ N_XI0/XI62/XI3/NET33_XI0/XI62/XI3/MM5_g N_VDD_XI0/XI62/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI3/MM4 N_XI0/XI62/XI3/NET33_XI0/XI62/XI3/MM4_d
+ N_XI0/XI62/XI3/NET34_XI0/XI62/XI3/MM4_g N_VDD_XI0/XI62/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI3/MM10 N_XI0/XI62/XI3/NET35_XI0/XI62/XI3/MM10_d
+ N_XI0/XI62/XI3/NET36_XI0/XI62/XI3/MM10_g N_VDD_XI0/XI62/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI3/MM11 N_XI0/XI62/XI3/NET36_XI0/XI62/XI3/MM11_d
+ N_XI0/XI62/XI3/NET35_XI0/XI62/XI3/MM11_g N_VDD_XI0/XI62/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI4/MM2 N_XI0/XI62/XI4/NET34_XI0/XI62/XI4/MM2_d
+ N_XI0/XI62/XI4/NET33_XI0/XI62/XI4/MM2_g N_VSS_XI0/XI62/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM3 N_XI0/XI62/XI4/NET33_XI0/XI62/XI4/MM3_d
+ N_WL<120>_XI0/XI62/XI4/MM3_g N_BLN<11>_XI0/XI62/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM0 N_XI0/XI62/XI4/NET34_XI0/XI62/XI4/MM0_d
+ N_WL<120>_XI0/XI62/XI4/MM0_g N_BL<11>_XI0/XI62/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM1 N_XI0/XI62/XI4/NET33_XI0/XI62/XI4/MM1_d
+ N_XI0/XI62/XI4/NET34_XI0/XI62/XI4/MM1_g N_VSS_XI0/XI62/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM9 N_XI0/XI62/XI4/NET36_XI0/XI62/XI4/MM9_d
+ N_WL<121>_XI0/XI62/XI4/MM9_g N_BL<11>_XI0/XI62/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM6 N_XI0/XI62/XI4/NET35_XI0/XI62/XI4/MM6_d
+ N_XI0/XI62/XI4/NET36_XI0/XI62/XI4/MM6_g N_VSS_XI0/XI62/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM7 N_XI0/XI62/XI4/NET36_XI0/XI62/XI4/MM7_d
+ N_XI0/XI62/XI4/NET35_XI0/XI62/XI4/MM7_g N_VSS_XI0/XI62/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM8 N_XI0/XI62/XI4/NET35_XI0/XI62/XI4/MM8_d
+ N_WL<121>_XI0/XI62/XI4/MM8_g N_BLN<11>_XI0/XI62/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI4/MM5 N_XI0/XI62/XI4/NET34_XI0/XI62/XI4/MM5_d
+ N_XI0/XI62/XI4/NET33_XI0/XI62/XI4/MM5_g N_VDD_XI0/XI62/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI4/MM4 N_XI0/XI62/XI4/NET33_XI0/XI62/XI4/MM4_d
+ N_XI0/XI62/XI4/NET34_XI0/XI62/XI4/MM4_g N_VDD_XI0/XI62/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI4/MM10 N_XI0/XI62/XI4/NET35_XI0/XI62/XI4/MM10_d
+ N_XI0/XI62/XI4/NET36_XI0/XI62/XI4/MM10_g N_VDD_XI0/XI62/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI4/MM11 N_XI0/XI62/XI4/NET36_XI0/XI62/XI4/MM11_d
+ N_XI0/XI62/XI4/NET35_XI0/XI62/XI4/MM11_g N_VDD_XI0/XI62/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI5/MM2 N_XI0/XI62/XI5/NET34_XI0/XI62/XI5/MM2_d
+ N_XI0/XI62/XI5/NET33_XI0/XI62/XI5/MM2_g N_VSS_XI0/XI62/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM3 N_XI0/XI62/XI5/NET33_XI0/XI62/XI5/MM3_d
+ N_WL<120>_XI0/XI62/XI5/MM3_g N_BLN<10>_XI0/XI62/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM0 N_XI0/XI62/XI5/NET34_XI0/XI62/XI5/MM0_d
+ N_WL<120>_XI0/XI62/XI5/MM0_g N_BL<10>_XI0/XI62/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM1 N_XI0/XI62/XI5/NET33_XI0/XI62/XI5/MM1_d
+ N_XI0/XI62/XI5/NET34_XI0/XI62/XI5/MM1_g N_VSS_XI0/XI62/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM9 N_XI0/XI62/XI5/NET36_XI0/XI62/XI5/MM9_d
+ N_WL<121>_XI0/XI62/XI5/MM9_g N_BL<10>_XI0/XI62/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM6 N_XI0/XI62/XI5/NET35_XI0/XI62/XI5/MM6_d
+ N_XI0/XI62/XI5/NET36_XI0/XI62/XI5/MM6_g N_VSS_XI0/XI62/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM7 N_XI0/XI62/XI5/NET36_XI0/XI62/XI5/MM7_d
+ N_XI0/XI62/XI5/NET35_XI0/XI62/XI5/MM7_g N_VSS_XI0/XI62/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM8 N_XI0/XI62/XI5/NET35_XI0/XI62/XI5/MM8_d
+ N_WL<121>_XI0/XI62/XI5/MM8_g N_BLN<10>_XI0/XI62/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI5/MM5 N_XI0/XI62/XI5/NET34_XI0/XI62/XI5/MM5_d
+ N_XI0/XI62/XI5/NET33_XI0/XI62/XI5/MM5_g N_VDD_XI0/XI62/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI5/MM4 N_XI0/XI62/XI5/NET33_XI0/XI62/XI5/MM4_d
+ N_XI0/XI62/XI5/NET34_XI0/XI62/XI5/MM4_g N_VDD_XI0/XI62/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI5/MM10 N_XI0/XI62/XI5/NET35_XI0/XI62/XI5/MM10_d
+ N_XI0/XI62/XI5/NET36_XI0/XI62/XI5/MM10_g N_VDD_XI0/XI62/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI5/MM11 N_XI0/XI62/XI5/NET36_XI0/XI62/XI5/MM11_d
+ N_XI0/XI62/XI5/NET35_XI0/XI62/XI5/MM11_g N_VDD_XI0/XI62/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI6/MM2 N_XI0/XI62/XI6/NET34_XI0/XI62/XI6/MM2_d
+ N_XI0/XI62/XI6/NET33_XI0/XI62/XI6/MM2_g N_VSS_XI0/XI62/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM3 N_XI0/XI62/XI6/NET33_XI0/XI62/XI6/MM3_d
+ N_WL<120>_XI0/XI62/XI6/MM3_g N_BLN<9>_XI0/XI62/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM0 N_XI0/XI62/XI6/NET34_XI0/XI62/XI6/MM0_d
+ N_WL<120>_XI0/XI62/XI6/MM0_g N_BL<9>_XI0/XI62/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM1 N_XI0/XI62/XI6/NET33_XI0/XI62/XI6/MM1_d
+ N_XI0/XI62/XI6/NET34_XI0/XI62/XI6/MM1_g N_VSS_XI0/XI62/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM9 N_XI0/XI62/XI6/NET36_XI0/XI62/XI6/MM9_d
+ N_WL<121>_XI0/XI62/XI6/MM9_g N_BL<9>_XI0/XI62/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM6 N_XI0/XI62/XI6/NET35_XI0/XI62/XI6/MM6_d
+ N_XI0/XI62/XI6/NET36_XI0/XI62/XI6/MM6_g N_VSS_XI0/XI62/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM7 N_XI0/XI62/XI6/NET36_XI0/XI62/XI6/MM7_d
+ N_XI0/XI62/XI6/NET35_XI0/XI62/XI6/MM7_g N_VSS_XI0/XI62/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM8 N_XI0/XI62/XI6/NET35_XI0/XI62/XI6/MM8_d
+ N_WL<121>_XI0/XI62/XI6/MM8_g N_BLN<9>_XI0/XI62/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI6/MM5 N_XI0/XI62/XI6/NET34_XI0/XI62/XI6/MM5_d
+ N_XI0/XI62/XI6/NET33_XI0/XI62/XI6/MM5_g N_VDD_XI0/XI62/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI6/MM4 N_XI0/XI62/XI6/NET33_XI0/XI62/XI6/MM4_d
+ N_XI0/XI62/XI6/NET34_XI0/XI62/XI6/MM4_g N_VDD_XI0/XI62/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI6/MM10 N_XI0/XI62/XI6/NET35_XI0/XI62/XI6/MM10_d
+ N_XI0/XI62/XI6/NET36_XI0/XI62/XI6/MM10_g N_VDD_XI0/XI62/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI6/MM11 N_XI0/XI62/XI6/NET36_XI0/XI62/XI6/MM11_d
+ N_XI0/XI62/XI6/NET35_XI0/XI62/XI6/MM11_g N_VDD_XI0/XI62/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI7/MM2 N_XI0/XI62/XI7/NET34_XI0/XI62/XI7/MM2_d
+ N_XI0/XI62/XI7/NET33_XI0/XI62/XI7/MM2_g N_VSS_XI0/XI62/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM3 N_XI0/XI62/XI7/NET33_XI0/XI62/XI7/MM3_d
+ N_WL<120>_XI0/XI62/XI7/MM3_g N_BLN<8>_XI0/XI62/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM0 N_XI0/XI62/XI7/NET34_XI0/XI62/XI7/MM0_d
+ N_WL<120>_XI0/XI62/XI7/MM0_g N_BL<8>_XI0/XI62/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM1 N_XI0/XI62/XI7/NET33_XI0/XI62/XI7/MM1_d
+ N_XI0/XI62/XI7/NET34_XI0/XI62/XI7/MM1_g N_VSS_XI0/XI62/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM9 N_XI0/XI62/XI7/NET36_XI0/XI62/XI7/MM9_d
+ N_WL<121>_XI0/XI62/XI7/MM9_g N_BL<8>_XI0/XI62/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM6 N_XI0/XI62/XI7/NET35_XI0/XI62/XI7/MM6_d
+ N_XI0/XI62/XI7/NET36_XI0/XI62/XI7/MM6_g N_VSS_XI0/XI62/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM7 N_XI0/XI62/XI7/NET36_XI0/XI62/XI7/MM7_d
+ N_XI0/XI62/XI7/NET35_XI0/XI62/XI7/MM7_g N_VSS_XI0/XI62/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM8 N_XI0/XI62/XI7/NET35_XI0/XI62/XI7/MM8_d
+ N_WL<121>_XI0/XI62/XI7/MM8_g N_BLN<8>_XI0/XI62/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI7/MM5 N_XI0/XI62/XI7/NET34_XI0/XI62/XI7/MM5_d
+ N_XI0/XI62/XI7/NET33_XI0/XI62/XI7/MM5_g N_VDD_XI0/XI62/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI7/MM4 N_XI0/XI62/XI7/NET33_XI0/XI62/XI7/MM4_d
+ N_XI0/XI62/XI7/NET34_XI0/XI62/XI7/MM4_g N_VDD_XI0/XI62/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI7/MM10 N_XI0/XI62/XI7/NET35_XI0/XI62/XI7/MM10_d
+ N_XI0/XI62/XI7/NET36_XI0/XI62/XI7/MM10_g N_VDD_XI0/XI62/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI7/MM11 N_XI0/XI62/XI7/NET36_XI0/XI62/XI7/MM11_d
+ N_XI0/XI62/XI7/NET35_XI0/XI62/XI7/MM11_g N_VDD_XI0/XI62/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI8/MM2 N_XI0/XI62/XI8/NET34_XI0/XI62/XI8/MM2_d
+ N_XI0/XI62/XI8/NET33_XI0/XI62/XI8/MM2_g N_VSS_XI0/XI62/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM3 N_XI0/XI62/XI8/NET33_XI0/XI62/XI8/MM3_d
+ N_WL<120>_XI0/XI62/XI8/MM3_g N_BLN<7>_XI0/XI62/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM0 N_XI0/XI62/XI8/NET34_XI0/XI62/XI8/MM0_d
+ N_WL<120>_XI0/XI62/XI8/MM0_g N_BL<7>_XI0/XI62/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM1 N_XI0/XI62/XI8/NET33_XI0/XI62/XI8/MM1_d
+ N_XI0/XI62/XI8/NET34_XI0/XI62/XI8/MM1_g N_VSS_XI0/XI62/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM9 N_XI0/XI62/XI8/NET36_XI0/XI62/XI8/MM9_d
+ N_WL<121>_XI0/XI62/XI8/MM9_g N_BL<7>_XI0/XI62/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM6 N_XI0/XI62/XI8/NET35_XI0/XI62/XI8/MM6_d
+ N_XI0/XI62/XI8/NET36_XI0/XI62/XI8/MM6_g N_VSS_XI0/XI62/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM7 N_XI0/XI62/XI8/NET36_XI0/XI62/XI8/MM7_d
+ N_XI0/XI62/XI8/NET35_XI0/XI62/XI8/MM7_g N_VSS_XI0/XI62/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM8 N_XI0/XI62/XI8/NET35_XI0/XI62/XI8/MM8_d
+ N_WL<121>_XI0/XI62/XI8/MM8_g N_BLN<7>_XI0/XI62/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI8/MM5 N_XI0/XI62/XI8/NET34_XI0/XI62/XI8/MM5_d
+ N_XI0/XI62/XI8/NET33_XI0/XI62/XI8/MM5_g N_VDD_XI0/XI62/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI8/MM4 N_XI0/XI62/XI8/NET33_XI0/XI62/XI8/MM4_d
+ N_XI0/XI62/XI8/NET34_XI0/XI62/XI8/MM4_g N_VDD_XI0/XI62/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI8/MM10 N_XI0/XI62/XI8/NET35_XI0/XI62/XI8/MM10_d
+ N_XI0/XI62/XI8/NET36_XI0/XI62/XI8/MM10_g N_VDD_XI0/XI62/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI8/MM11 N_XI0/XI62/XI8/NET36_XI0/XI62/XI8/MM11_d
+ N_XI0/XI62/XI8/NET35_XI0/XI62/XI8/MM11_g N_VDD_XI0/XI62/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI9/MM2 N_XI0/XI62/XI9/NET34_XI0/XI62/XI9/MM2_d
+ N_XI0/XI62/XI9/NET33_XI0/XI62/XI9/MM2_g N_VSS_XI0/XI62/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM3 N_XI0/XI62/XI9/NET33_XI0/XI62/XI9/MM3_d
+ N_WL<120>_XI0/XI62/XI9/MM3_g N_BLN<6>_XI0/XI62/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM0 N_XI0/XI62/XI9/NET34_XI0/XI62/XI9/MM0_d
+ N_WL<120>_XI0/XI62/XI9/MM0_g N_BL<6>_XI0/XI62/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM1 N_XI0/XI62/XI9/NET33_XI0/XI62/XI9/MM1_d
+ N_XI0/XI62/XI9/NET34_XI0/XI62/XI9/MM1_g N_VSS_XI0/XI62/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM9 N_XI0/XI62/XI9/NET36_XI0/XI62/XI9/MM9_d
+ N_WL<121>_XI0/XI62/XI9/MM9_g N_BL<6>_XI0/XI62/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM6 N_XI0/XI62/XI9/NET35_XI0/XI62/XI9/MM6_d
+ N_XI0/XI62/XI9/NET36_XI0/XI62/XI9/MM6_g N_VSS_XI0/XI62/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM7 N_XI0/XI62/XI9/NET36_XI0/XI62/XI9/MM7_d
+ N_XI0/XI62/XI9/NET35_XI0/XI62/XI9/MM7_g N_VSS_XI0/XI62/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM8 N_XI0/XI62/XI9/NET35_XI0/XI62/XI9/MM8_d
+ N_WL<121>_XI0/XI62/XI9/MM8_g N_BLN<6>_XI0/XI62/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI9/MM5 N_XI0/XI62/XI9/NET34_XI0/XI62/XI9/MM5_d
+ N_XI0/XI62/XI9/NET33_XI0/XI62/XI9/MM5_g N_VDD_XI0/XI62/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI9/MM4 N_XI0/XI62/XI9/NET33_XI0/XI62/XI9/MM4_d
+ N_XI0/XI62/XI9/NET34_XI0/XI62/XI9/MM4_g N_VDD_XI0/XI62/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI9/MM10 N_XI0/XI62/XI9/NET35_XI0/XI62/XI9/MM10_d
+ N_XI0/XI62/XI9/NET36_XI0/XI62/XI9/MM10_g N_VDD_XI0/XI62/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI9/MM11 N_XI0/XI62/XI9/NET36_XI0/XI62/XI9/MM11_d
+ N_XI0/XI62/XI9/NET35_XI0/XI62/XI9/MM11_g N_VDD_XI0/XI62/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI10/MM2 N_XI0/XI62/XI10/NET34_XI0/XI62/XI10/MM2_d
+ N_XI0/XI62/XI10/NET33_XI0/XI62/XI10/MM2_g N_VSS_XI0/XI62/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM3 N_XI0/XI62/XI10/NET33_XI0/XI62/XI10/MM3_d
+ N_WL<120>_XI0/XI62/XI10/MM3_g N_BLN<5>_XI0/XI62/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM0 N_XI0/XI62/XI10/NET34_XI0/XI62/XI10/MM0_d
+ N_WL<120>_XI0/XI62/XI10/MM0_g N_BL<5>_XI0/XI62/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM1 N_XI0/XI62/XI10/NET33_XI0/XI62/XI10/MM1_d
+ N_XI0/XI62/XI10/NET34_XI0/XI62/XI10/MM1_g N_VSS_XI0/XI62/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM9 N_XI0/XI62/XI10/NET36_XI0/XI62/XI10/MM9_d
+ N_WL<121>_XI0/XI62/XI10/MM9_g N_BL<5>_XI0/XI62/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM6 N_XI0/XI62/XI10/NET35_XI0/XI62/XI10/MM6_d
+ N_XI0/XI62/XI10/NET36_XI0/XI62/XI10/MM6_g N_VSS_XI0/XI62/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM7 N_XI0/XI62/XI10/NET36_XI0/XI62/XI10/MM7_d
+ N_XI0/XI62/XI10/NET35_XI0/XI62/XI10/MM7_g N_VSS_XI0/XI62/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM8 N_XI0/XI62/XI10/NET35_XI0/XI62/XI10/MM8_d
+ N_WL<121>_XI0/XI62/XI10/MM8_g N_BLN<5>_XI0/XI62/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI10/MM5 N_XI0/XI62/XI10/NET34_XI0/XI62/XI10/MM5_d
+ N_XI0/XI62/XI10/NET33_XI0/XI62/XI10/MM5_g N_VDD_XI0/XI62/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI10/MM4 N_XI0/XI62/XI10/NET33_XI0/XI62/XI10/MM4_d
+ N_XI0/XI62/XI10/NET34_XI0/XI62/XI10/MM4_g N_VDD_XI0/XI62/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI10/MM10 N_XI0/XI62/XI10/NET35_XI0/XI62/XI10/MM10_d
+ N_XI0/XI62/XI10/NET36_XI0/XI62/XI10/MM10_g N_VDD_XI0/XI62/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI10/MM11 N_XI0/XI62/XI10/NET36_XI0/XI62/XI10/MM11_d
+ N_XI0/XI62/XI10/NET35_XI0/XI62/XI10/MM11_g N_VDD_XI0/XI62/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI11/MM2 N_XI0/XI62/XI11/NET34_XI0/XI62/XI11/MM2_d
+ N_XI0/XI62/XI11/NET33_XI0/XI62/XI11/MM2_g N_VSS_XI0/XI62/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM3 N_XI0/XI62/XI11/NET33_XI0/XI62/XI11/MM3_d
+ N_WL<120>_XI0/XI62/XI11/MM3_g N_BLN<4>_XI0/XI62/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM0 N_XI0/XI62/XI11/NET34_XI0/XI62/XI11/MM0_d
+ N_WL<120>_XI0/XI62/XI11/MM0_g N_BL<4>_XI0/XI62/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM1 N_XI0/XI62/XI11/NET33_XI0/XI62/XI11/MM1_d
+ N_XI0/XI62/XI11/NET34_XI0/XI62/XI11/MM1_g N_VSS_XI0/XI62/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM9 N_XI0/XI62/XI11/NET36_XI0/XI62/XI11/MM9_d
+ N_WL<121>_XI0/XI62/XI11/MM9_g N_BL<4>_XI0/XI62/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM6 N_XI0/XI62/XI11/NET35_XI0/XI62/XI11/MM6_d
+ N_XI0/XI62/XI11/NET36_XI0/XI62/XI11/MM6_g N_VSS_XI0/XI62/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM7 N_XI0/XI62/XI11/NET36_XI0/XI62/XI11/MM7_d
+ N_XI0/XI62/XI11/NET35_XI0/XI62/XI11/MM7_g N_VSS_XI0/XI62/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM8 N_XI0/XI62/XI11/NET35_XI0/XI62/XI11/MM8_d
+ N_WL<121>_XI0/XI62/XI11/MM8_g N_BLN<4>_XI0/XI62/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI11/MM5 N_XI0/XI62/XI11/NET34_XI0/XI62/XI11/MM5_d
+ N_XI0/XI62/XI11/NET33_XI0/XI62/XI11/MM5_g N_VDD_XI0/XI62/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI11/MM4 N_XI0/XI62/XI11/NET33_XI0/XI62/XI11/MM4_d
+ N_XI0/XI62/XI11/NET34_XI0/XI62/XI11/MM4_g N_VDD_XI0/XI62/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI11/MM10 N_XI0/XI62/XI11/NET35_XI0/XI62/XI11/MM10_d
+ N_XI0/XI62/XI11/NET36_XI0/XI62/XI11/MM10_g N_VDD_XI0/XI62/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI11/MM11 N_XI0/XI62/XI11/NET36_XI0/XI62/XI11/MM11_d
+ N_XI0/XI62/XI11/NET35_XI0/XI62/XI11/MM11_g N_VDD_XI0/XI62/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI12/MM2 N_XI0/XI62/XI12/NET34_XI0/XI62/XI12/MM2_d
+ N_XI0/XI62/XI12/NET33_XI0/XI62/XI12/MM2_g N_VSS_XI0/XI62/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM3 N_XI0/XI62/XI12/NET33_XI0/XI62/XI12/MM3_d
+ N_WL<120>_XI0/XI62/XI12/MM3_g N_BLN<3>_XI0/XI62/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM0 N_XI0/XI62/XI12/NET34_XI0/XI62/XI12/MM0_d
+ N_WL<120>_XI0/XI62/XI12/MM0_g N_BL<3>_XI0/XI62/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM1 N_XI0/XI62/XI12/NET33_XI0/XI62/XI12/MM1_d
+ N_XI0/XI62/XI12/NET34_XI0/XI62/XI12/MM1_g N_VSS_XI0/XI62/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM9 N_XI0/XI62/XI12/NET36_XI0/XI62/XI12/MM9_d
+ N_WL<121>_XI0/XI62/XI12/MM9_g N_BL<3>_XI0/XI62/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM6 N_XI0/XI62/XI12/NET35_XI0/XI62/XI12/MM6_d
+ N_XI0/XI62/XI12/NET36_XI0/XI62/XI12/MM6_g N_VSS_XI0/XI62/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM7 N_XI0/XI62/XI12/NET36_XI0/XI62/XI12/MM7_d
+ N_XI0/XI62/XI12/NET35_XI0/XI62/XI12/MM7_g N_VSS_XI0/XI62/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM8 N_XI0/XI62/XI12/NET35_XI0/XI62/XI12/MM8_d
+ N_WL<121>_XI0/XI62/XI12/MM8_g N_BLN<3>_XI0/XI62/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI12/MM5 N_XI0/XI62/XI12/NET34_XI0/XI62/XI12/MM5_d
+ N_XI0/XI62/XI12/NET33_XI0/XI62/XI12/MM5_g N_VDD_XI0/XI62/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI12/MM4 N_XI0/XI62/XI12/NET33_XI0/XI62/XI12/MM4_d
+ N_XI0/XI62/XI12/NET34_XI0/XI62/XI12/MM4_g N_VDD_XI0/XI62/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI12/MM10 N_XI0/XI62/XI12/NET35_XI0/XI62/XI12/MM10_d
+ N_XI0/XI62/XI12/NET36_XI0/XI62/XI12/MM10_g N_VDD_XI0/XI62/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI12/MM11 N_XI0/XI62/XI12/NET36_XI0/XI62/XI12/MM11_d
+ N_XI0/XI62/XI12/NET35_XI0/XI62/XI12/MM11_g N_VDD_XI0/XI62/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI13/MM2 N_XI0/XI62/XI13/NET34_XI0/XI62/XI13/MM2_d
+ N_XI0/XI62/XI13/NET33_XI0/XI62/XI13/MM2_g N_VSS_XI0/XI62/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM3 N_XI0/XI62/XI13/NET33_XI0/XI62/XI13/MM3_d
+ N_WL<120>_XI0/XI62/XI13/MM3_g N_BLN<2>_XI0/XI62/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM0 N_XI0/XI62/XI13/NET34_XI0/XI62/XI13/MM0_d
+ N_WL<120>_XI0/XI62/XI13/MM0_g N_BL<2>_XI0/XI62/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM1 N_XI0/XI62/XI13/NET33_XI0/XI62/XI13/MM1_d
+ N_XI0/XI62/XI13/NET34_XI0/XI62/XI13/MM1_g N_VSS_XI0/XI62/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM9 N_XI0/XI62/XI13/NET36_XI0/XI62/XI13/MM9_d
+ N_WL<121>_XI0/XI62/XI13/MM9_g N_BL<2>_XI0/XI62/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM6 N_XI0/XI62/XI13/NET35_XI0/XI62/XI13/MM6_d
+ N_XI0/XI62/XI13/NET36_XI0/XI62/XI13/MM6_g N_VSS_XI0/XI62/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM7 N_XI0/XI62/XI13/NET36_XI0/XI62/XI13/MM7_d
+ N_XI0/XI62/XI13/NET35_XI0/XI62/XI13/MM7_g N_VSS_XI0/XI62/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM8 N_XI0/XI62/XI13/NET35_XI0/XI62/XI13/MM8_d
+ N_WL<121>_XI0/XI62/XI13/MM8_g N_BLN<2>_XI0/XI62/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI13/MM5 N_XI0/XI62/XI13/NET34_XI0/XI62/XI13/MM5_d
+ N_XI0/XI62/XI13/NET33_XI0/XI62/XI13/MM5_g N_VDD_XI0/XI62/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI13/MM4 N_XI0/XI62/XI13/NET33_XI0/XI62/XI13/MM4_d
+ N_XI0/XI62/XI13/NET34_XI0/XI62/XI13/MM4_g N_VDD_XI0/XI62/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI13/MM10 N_XI0/XI62/XI13/NET35_XI0/XI62/XI13/MM10_d
+ N_XI0/XI62/XI13/NET36_XI0/XI62/XI13/MM10_g N_VDD_XI0/XI62/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI13/MM11 N_XI0/XI62/XI13/NET36_XI0/XI62/XI13/MM11_d
+ N_XI0/XI62/XI13/NET35_XI0/XI62/XI13/MM11_g N_VDD_XI0/XI62/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI14/MM2 N_XI0/XI62/XI14/NET34_XI0/XI62/XI14/MM2_d
+ N_XI0/XI62/XI14/NET33_XI0/XI62/XI14/MM2_g N_VSS_XI0/XI62/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM3 N_XI0/XI62/XI14/NET33_XI0/XI62/XI14/MM3_d
+ N_WL<120>_XI0/XI62/XI14/MM3_g N_BLN<1>_XI0/XI62/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM0 N_XI0/XI62/XI14/NET34_XI0/XI62/XI14/MM0_d
+ N_WL<120>_XI0/XI62/XI14/MM0_g N_BL<1>_XI0/XI62/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM1 N_XI0/XI62/XI14/NET33_XI0/XI62/XI14/MM1_d
+ N_XI0/XI62/XI14/NET34_XI0/XI62/XI14/MM1_g N_VSS_XI0/XI62/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM9 N_XI0/XI62/XI14/NET36_XI0/XI62/XI14/MM9_d
+ N_WL<121>_XI0/XI62/XI14/MM9_g N_BL<1>_XI0/XI62/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM6 N_XI0/XI62/XI14/NET35_XI0/XI62/XI14/MM6_d
+ N_XI0/XI62/XI14/NET36_XI0/XI62/XI14/MM6_g N_VSS_XI0/XI62/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM7 N_XI0/XI62/XI14/NET36_XI0/XI62/XI14/MM7_d
+ N_XI0/XI62/XI14/NET35_XI0/XI62/XI14/MM7_g N_VSS_XI0/XI62/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM8 N_XI0/XI62/XI14/NET35_XI0/XI62/XI14/MM8_d
+ N_WL<121>_XI0/XI62/XI14/MM8_g N_BLN<1>_XI0/XI62/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI14/MM5 N_XI0/XI62/XI14/NET34_XI0/XI62/XI14/MM5_d
+ N_XI0/XI62/XI14/NET33_XI0/XI62/XI14/MM5_g N_VDD_XI0/XI62/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI14/MM4 N_XI0/XI62/XI14/NET33_XI0/XI62/XI14/MM4_d
+ N_XI0/XI62/XI14/NET34_XI0/XI62/XI14/MM4_g N_VDD_XI0/XI62/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI14/MM10 N_XI0/XI62/XI14/NET35_XI0/XI62/XI14/MM10_d
+ N_XI0/XI62/XI14/NET36_XI0/XI62/XI14/MM10_g N_VDD_XI0/XI62/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI14/MM11 N_XI0/XI62/XI14/NET36_XI0/XI62/XI14/MM11_d
+ N_XI0/XI62/XI14/NET35_XI0/XI62/XI14/MM11_g N_VDD_XI0/XI62/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI15/MM2 N_XI0/XI62/XI15/NET34_XI0/XI62/XI15/MM2_d
+ N_XI0/XI62/XI15/NET33_XI0/XI62/XI15/MM2_g N_VSS_XI0/XI62/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM3 N_XI0/XI62/XI15/NET33_XI0/XI62/XI15/MM3_d
+ N_WL<120>_XI0/XI62/XI15/MM3_g N_BLN<0>_XI0/XI62/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM0 N_XI0/XI62/XI15/NET34_XI0/XI62/XI15/MM0_d
+ N_WL<120>_XI0/XI62/XI15/MM0_g N_BL<0>_XI0/XI62/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM1 N_XI0/XI62/XI15/NET33_XI0/XI62/XI15/MM1_d
+ N_XI0/XI62/XI15/NET34_XI0/XI62/XI15/MM1_g N_VSS_XI0/XI62/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM9 N_XI0/XI62/XI15/NET36_XI0/XI62/XI15/MM9_d
+ N_WL<121>_XI0/XI62/XI15/MM9_g N_BL<0>_XI0/XI62/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM6 N_XI0/XI62/XI15/NET35_XI0/XI62/XI15/MM6_d
+ N_XI0/XI62/XI15/NET36_XI0/XI62/XI15/MM6_g N_VSS_XI0/XI62/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM7 N_XI0/XI62/XI15/NET36_XI0/XI62/XI15/MM7_d
+ N_XI0/XI62/XI15/NET35_XI0/XI62/XI15/MM7_g N_VSS_XI0/XI62/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM8 N_XI0/XI62/XI15/NET35_XI0/XI62/XI15/MM8_d
+ N_WL<121>_XI0/XI62/XI15/MM8_g N_BLN<0>_XI0/XI62/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI62/XI15/MM5 N_XI0/XI62/XI15/NET34_XI0/XI62/XI15/MM5_d
+ N_XI0/XI62/XI15/NET33_XI0/XI62/XI15/MM5_g N_VDD_XI0/XI62/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI15/MM4 N_XI0/XI62/XI15/NET33_XI0/XI62/XI15/MM4_d
+ N_XI0/XI62/XI15/NET34_XI0/XI62/XI15/MM4_g N_VDD_XI0/XI62/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI15/MM10 N_XI0/XI62/XI15/NET35_XI0/XI62/XI15/MM10_d
+ N_XI0/XI62/XI15/NET36_XI0/XI62/XI15/MM10_g N_VDD_XI0/XI62/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI62/XI15/MM11 N_XI0/XI62/XI15/NET36_XI0/XI62/XI15/MM11_d
+ N_XI0/XI62/XI15/NET35_XI0/XI62/XI15/MM11_g N_VDD_XI0/XI62/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI0/MM2 N_XI0/XI63/XI0/NET34_XI0/XI63/XI0/MM2_d
+ N_XI0/XI63/XI0/NET33_XI0/XI63/XI0/MM2_g N_VSS_XI0/XI63/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM3 N_XI0/XI63/XI0/NET33_XI0/XI63/XI0/MM3_d
+ N_WL<122>_XI0/XI63/XI0/MM3_g N_BLN<15>_XI0/XI63/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM0 N_XI0/XI63/XI0/NET34_XI0/XI63/XI0/MM0_d
+ N_WL<122>_XI0/XI63/XI0/MM0_g N_BL<15>_XI0/XI63/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM1 N_XI0/XI63/XI0/NET33_XI0/XI63/XI0/MM1_d
+ N_XI0/XI63/XI0/NET34_XI0/XI63/XI0/MM1_g N_VSS_XI0/XI63/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM9 N_XI0/XI63/XI0/NET36_XI0/XI63/XI0/MM9_d
+ N_WL<123>_XI0/XI63/XI0/MM9_g N_BL<15>_XI0/XI63/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM6 N_XI0/XI63/XI0/NET35_XI0/XI63/XI0/MM6_d
+ N_XI0/XI63/XI0/NET36_XI0/XI63/XI0/MM6_g N_VSS_XI0/XI63/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM7 N_XI0/XI63/XI0/NET36_XI0/XI63/XI0/MM7_d
+ N_XI0/XI63/XI0/NET35_XI0/XI63/XI0/MM7_g N_VSS_XI0/XI63/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM8 N_XI0/XI63/XI0/NET35_XI0/XI63/XI0/MM8_d
+ N_WL<123>_XI0/XI63/XI0/MM8_g N_BLN<15>_XI0/XI63/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI0/MM5 N_XI0/XI63/XI0/NET34_XI0/XI63/XI0/MM5_d
+ N_XI0/XI63/XI0/NET33_XI0/XI63/XI0/MM5_g N_VDD_XI0/XI63/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI0/MM4 N_XI0/XI63/XI0/NET33_XI0/XI63/XI0/MM4_d
+ N_XI0/XI63/XI0/NET34_XI0/XI63/XI0/MM4_g N_VDD_XI0/XI63/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI0/MM10 N_XI0/XI63/XI0/NET35_XI0/XI63/XI0/MM10_d
+ N_XI0/XI63/XI0/NET36_XI0/XI63/XI0/MM10_g N_VDD_XI0/XI63/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI0/MM11 N_XI0/XI63/XI0/NET36_XI0/XI63/XI0/MM11_d
+ N_XI0/XI63/XI0/NET35_XI0/XI63/XI0/MM11_g N_VDD_XI0/XI63/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI1/MM2 N_XI0/XI63/XI1/NET34_XI0/XI63/XI1/MM2_d
+ N_XI0/XI63/XI1/NET33_XI0/XI63/XI1/MM2_g N_VSS_XI0/XI63/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM3 N_XI0/XI63/XI1/NET33_XI0/XI63/XI1/MM3_d
+ N_WL<122>_XI0/XI63/XI1/MM3_g N_BLN<14>_XI0/XI63/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM0 N_XI0/XI63/XI1/NET34_XI0/XI63/XI1/MM0_d
+ N_WL<122>_XI0/XI63/XI1/MM0_g N_BL<14>_XI0/XI63/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM1 N_XI0/XI63/XI1/NET33_XI0/XI63/XI1/MM1_d
+ N_XI0/XI63/XI1/NET34_XI0/XI63/XI1/MM1_g N_VSS_XI0/XI63/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM9 N_XI0/XI63/XI1/NET36_XI0/XI63/XI1/MM9_d
+ N_WL<123>_XI0/XI63/XI1/MM9_g N_BL<14>_XI0/XI63/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM6 N_XI0/XI63/XI1/NET35_XI0/XI63/XI1/MM6_d
+ N_XI0/XI63/XI1/NET36_XI0/XI63/XI1/MM6_g N_VSS_XI0/XI63/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM7 N_XI0/XI63/XI1/NET36_XI0/XI63/XI1/MM7_d
+ N_XI0/XI63/XI1/NET35_XI0/XI63/XI1/MM7_g N_VSS_XI0/XI63/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM8 N_XI0/XI63/XI1/NET35_XI0/XI63/XI1/MM8_d
+ N_WL<123>_XI0/XI63/XI1/MM8_g N_BLN<14>_XI0/XI63/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI1/MM5 N_XI0/XI63/XI1/NET34_XI0/XI63/XI1/MM5_d
+ N_XI0/XI63/XI1/NET33_XI0/XI63/XI1/MM5_g N_VDD_XI0/XI63/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI1/MM4 N_XI0/XI63/XI1/NET33_XI0/XI63/XI1/MM4_d
+ N_XI0/XI63/XI1/NET34_XI0/XI63/XI1/MM4_g N_VDD_XI0/XI63/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI1/MM10 N_XI0/XI63/XI1/NET35_XI0/XI63/XI1/MM10_d
+ N_XI0/XI63/XI1/NET36_XI0/XI63/XI1/MM10_g N_VDD_XI0/XI63/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI1/MM11 N_XI0/XI63/XI1/NET36_XI0/XI63/XI1/MM11_d
+ N_XI0/XI63/XI1/NET35_XI0/XI63/XI1/MM11_g N_VDD_XI0/XI63/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI2/MM2 N_XI0/XI63/XI2/NET34_XI0/XI63/XI2/MM2_d
+ N_XI0/XI63/XI2/NET33_XI0/XI63/XI2/MM2_g N_VSS_XI0/XI63/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM3 N_XI0/XI63/XI2/NET33_XI0/XI63/XI2/MM3_d
+ N_WL<122>_XI0/XI63/XI2/MM3_g N_BLN<13>_XI0/XI63/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM0 N_XI0/XI63/XI2/NET34_XI0/XI63/XI2/MM0_d
+ N_WL<122>_XI0/XI63/XI2/MM0_g N_BL<13>_XI0/XI63/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM1 N_XI0/XI63/XI2/NET33_XI0/XI63/XI2/MM1_d
+ N_XI0/XI63/XI2/NET34_XI0/XI63/XI2/MM1_g N_VSS_XI0/XI63/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM9 N_XI0/XI63/XI2/NET36_XI0/XI63/XI2/MM9_d
+ N_WL<123>_XI0/XI63/XI2/MM9_g N_BL<13>_XI0/XI63/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM6 N_XI0/XI63/XI2/NET35_XI0/XI63/XI2/MM6_d
+ N_XI0/XI63/XI2/NET36_XI0/XI63/XI2/MM6_g N_VSS_XI0/XI63/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM7 N_XI0/XI63/XI2/NET36_XI0/XI63/XI2/MM7_d
+ N_XI0/XI63/XI2/NET35_XI0/XI63/XI2/MM7_g N_VSS_XI0/XI63/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM8 N_XI0/XI63/XI2/NET35_XI0/XI63/XI2/MM8_d
+ N_WL<123>_XI0/XI63/XI2/MM8_g N_BLN<13>_XI0/XI63/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI2/MM5 N_XI0/XI63/XI2/NET34_XI0/XI63/XI2/MM5_d
+ N_XI0/XI63/XI2/NET33_XI0/XI63/XI2/MM5_g N_VDD_XI0/XI63/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI2/MM4 N_XI0/XI63/XI2/NET33_XI0/XI63/XI2/MM4_d
+ N_XI0/XI63/XI2/NET34_XI0/XI63/XI2/MM4_g N_VDD_XI0/XI63/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI2/MM10 N_XI0/XI63/XI2/NET35_XI0/XI63/XI2/MM10_d
+ N_XI0/XI63/XI2/NET36_XI0/XI63/XI2/MM10_g N_VDD_XI0/XI63/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI2/MM11 N_XI0/XI63/XI2/NET36_XI0/XI63/XI2/MM11_d
+ N_XI0/XI63/XI2/NET35_XI0/XI63/XI2/MM11_g N_VDD_XI0/XI63/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI3/MM2 N_XI0/XI63/XI3/NET34_XI0/XI63/XI3/MM2_d
+ N_XI0/XI63/XI3/NET33_XI0/XI63/XI3/MM2_g N_VSS_XI0/XI63/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM3 N_XI0/XI63/XI3/NET33_XI0/XI63/XI3/MM3_d
+ N_WL<122>_XI0/XI63/XI3/MM3_g N_BLN<12>_XI0/XI63/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM0 N_XI0/XI63/XI3/NET34_XI0/XI63/XI3/MM0_d
+ N_WL<122>_XI0/XI63/XI3/MM0_g N_BL<12>_XI0/XI63/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM1 N_XI0/XI63/XI3/NET33_XI0/XI63/XI3/MM1_d
+ N_XI0/XI63/XI3/NET34_XI0/XI63/XI3/MM1_g N_VSS_XI0/XI63/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM9 N_XI0/XI63/XI3/NET36_XI0/XI63/XI3/MM9_d
+ N_WL<123>_XI0/XI63/XI3/MM9_g N_BL<12>_XI0/XI63/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM6 N_XI0/XI63/XI3/NET35_XI0/XI63/XI3/MM6_d
+ N_XI0/XI63/XI3/NET36_XI0/XI63/XI3/MM6_g N_VSS_XI0/XI63/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM7 N_XI0/XI63/XI3/NET36_XI0/XI63/XI3/MM7_d
+ N_XI0/XI63/XI3/NET35_XI0/XI63/XI3/MM7_g N_VSS_XI0/XI63/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM8 N_XI0/XI63/XI3/NET35_XI0/XI63/XI3/MM8_d
+ N_WL<123>_XI0/XI63/XI3/MM8_g N_BLN<12>_XI0/XI63/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI3/MM5 N_XI0/XI63/XI3/NET34_XI0/XI63/XI3/MM5_d
+ N_XI0/XI63/XI3/NET33_XI0/XI63/XI3/MM5_g N_VDD_XI0/XI63/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI3/MM4 N_XI0/XI63/XI3/NET33_XI0/XI63/XI3/MM4_d
+ N_XI0/XI63/XI3/NET34_XI0/XI63/XI3/MM4_g N_VDD_XI0/XI63/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI3/MM10 N_XI0/XI63/XI3/NET35_XI0/XI63/XI3/MM10_d
+ N_XI0/XI63/XI3/NET36_XI0/XI63/XI3/MM10_g N_VDD_XI0/XI63/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI3/MM11 N_XI0/XI63/XI3/NET36_XI0/XI63/XI3/MM11_d
+ N_XI0/XI63/XI3/NET35_XI0/XI63/XI3/MM11_g N_VDD_XI0/XI63/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI4/MM2 N_XI0/XI63/XI4/NET34_XI0/XI63/XI4/MM2_d
+ N_XI0/XI63/XI4/NET33_XI0/XI63/XI4/MM2_g N_VSS_XI0/XI63/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM3 N_XI0/XI63/XI4/NET33_XI0/XI63/XI4/MM3_d
+ N_WL<122>_XI0/XI63/XI4/MM3_g N_BLN<11>_XI0/XI63/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM0 N_XI0/XI63/XI4/NET34_XI0/XI63/XI4/MM0_d
+ N_WL<122>_XI0/XI63/XI4/MM0_g N_BL<11>_XI0/XI63/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM1 N_XI0/XI63/XI4/NET33_XI0/XI63/XI4/MM1_d
+ N_XI0/XI63/XI4/NET34_XI0/XI63/XI4/MM1_g N_VSS_XI0/XI63/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM9 N_XI0/XI63/XI4/NET36_XI0/XI63/XI4/MM9_d
+ N_WL<123>_XI0/XI63/XI4/MM9_g N_BL<11>_XI0/XI63/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM6 N_XI0/XI63/XI4/NET35_XI0/XI63/XI4/MM6_d
+ N_XI0/XI63/XI4/NET36_XI0/XI63/XI4/MM6_g N_VSS_XI0/XI63/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM7 N_XI0/XI63/XI4/NET36_XI0/XI63/XI4/MM7_d
+ N_XI0/XI63/XI4/NET35_XI0/XI63/XI4/MM7_g N_VSS_XI0/XI63/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM8 N_XI0/XI63/XI4/NET35_XI0/XI63/XI4/MM8_d
+ N_WL<123>_XI0/XI63/XI4/MM8_g N_BLN<11>_XI0/XI63/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI4/MM5 N_XI0/XI63/XI4/NET34_XI0/XI63/XI4/MM5_d
+ N_XI0/XI63/XI4/NET33_XI0/XI63/XI4/MM5_g N_VDD_XI0/XI63/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI4/MM4 N_XI0/XI63/XI4/NET33_XI0/XI63/XI4/MM4_d
+ N_XI0/XI63/XI4/NET34_XI0/XI63/XI4/MM4_g N_VDD_XI0/XI63/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI4/MM10 N_XI0/XI63/XI4/NET35_XI0/XI63/XI4/MM10_d
+ N_XI0/XI63/XI4/NET36_XI0/XI63/XI4/MM10_g N_VDD_XI0/XI63/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI4/MM11 N_XI0/XI63/XI4/NET36_XI0/XI63/XI4/MM11_d
+ N_XI0/XI63/XI4/NET35_XI0/XI63/XI4/MM11_g N_VDD_XI0/XI63/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI5/MM2 N_XI0/XI63/XI5/NET34_XI0/XI63/XI5/MM2_d
+ N_XI0/XI63/XI5/NET33_XI0/XI63/XI5/MM2_g N_VSS_XI0/XI63/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM3 N_XI0/XI63/XI5/NET33_XI0/XI63/XI5/MM3_d
+ N_WL<122>_XI0/XI63/XI5/MM3_g N_BLN<10>_XI0/XI63/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM0 N_XI0/XI63/XI5/NET34_XI0/XI63/XI5/MM0_d
+ N_WL<122>_XI0/XI63/XI5/MM0_g N_BL<10>_XI0/XI63/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM1 N_XI0/XI63/XI5/NET33_XI0/XI63/XI5/MM1_d
+ N_XI0/XI63/XI5/NET34_XI0/XI63/XI5/MM1_g N_VSS_XI0/XI63/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM9 N_XI0/XI63/XI5/NET36_XI0/XI63/XI5/MM9_d
+ N_WL<123>_XI0/XI63/XI5/MM9_g N_BL<10>_XI0/XI63/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM6 N_XI0/XI63/XI5/NET35_XI0/XI63/XI5/MM6_d
+ N_XI0/XI63/XI5/NET36_XI0/XI63/XI5/MM6_g N_VSS_XI0/XI63/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM7 N_XI0/XI63/XI5/NET36_XI0/XI63/XI5/MM7_d
+ N_XI0/XI63/XI5/NET35_XI0/XI63/XI5/MM7_g N_VSS_XI0/XI63/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM8 N_XI0/XI63/XI5/NET35_XI0/XI63/XI5/MM8_d
+ N_WL<123>_XI0/XI63/XI5/MM8_g N_BLN<10>_XI0/XI63/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI5/MM5 N_XI0/XI63/XI5/NET34_XI0/XI63/XI5/MM5_d
+ N_XI0/XI63/XI5/NET33_XI0/XI63/XI5/MM5_g N_VDD_XI0/XI63/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI5/MM4 N_XI0/XI63/XI5/NET33_XI0/XI63/XI5/MM4_d
+ N_XI0/XI63/XI5/NET34_XI0/XI63/XI5/MM4_g N_VDD_XI0/XI63/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI5/MM10 N_XI0/XI63/XI5/NET35_XI0/XI63/XI5/MM10_d
+ N_XI0/XI63/XI5/NET36_XI0/XI63/XI5/MM10_g N_VDD_XI0/XI63/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI5/MM11 N_XI0/XI63/XI5/NET36_XI0/XI63/XI5/MM11_d
+ N_XI0/XI63/XI5/NET35_XI0/XI63/XI5/MM11_g N_VDD_XI0/XI63/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI6/MM2 N_XI0/XI63/XI6/NET34_XI0/XI63/XI6/MM2_d
+ N_XI0/XI63/XI6/NET33_XI0/XI63/XI6/MM2_g N_VSS_XI0/XI63/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM3 N_XI0/XI63/XI6/NET33_XI0/XI63/XI6/MM3_d
+ N_WL<122>_XI0/XI63/XI6/MM3_g N_BLN<9>_XI0/XI63/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM0 N_XI0/XI63/XI6/NET34_XI0/XI63/XI6/MM0_d
+ N_WL<122>_XI0/XI63/XI6/MM0_g N_BL<9>_XI0/XI63/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM1 N_XI0/XI63/XI6/NET33_XI0/XI63/XI6/MM1_d
+ N_XI0/XI63/XI6/NET34_XI0/XI63/XI6/MM1_g N_VSS_XI0/XI63/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM9 N_XI0/XI63/XI6/NET36_XI0/XI63/XI6/MM9_d
+ N_WL<123>_XI0/XI63/XI6/MM9_g N_BL<9>_XI0/XI63/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM6 N_XI0/XI63/XI6/NET35_XI0/XI63/XI6/MM6_d
+ N_XI0/XI63/XI6/NET36_XI0/XI63/XI6/MM6_g N_VSS_XI0/XI63/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM7 N_XI0/XI63/XI6/NET36_XI0/XI63/XI6/MM7_d
+ N_XI0/XI63/XI6/NET35_XI0/XI63/XI6/MM7_g N_VSS_XI0/XI63/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM8 N_XI0/XI63/XI6/NET35_XI0/XI63/XI6/MM8_d
+ N_WL<123>_XI0/XI63/XI6/MM8_g N_BLN<9>_XI0/XI63/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI6/MM5 N_XI0/XI63/XI6/NET34_XI0/XI63/XI6/MM5_d
+ N_XI0/XI63/XI6/NET33_XI0/XI63/XI6/MM5_g N_VDD_XI0/XI63/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI6/MM4 N_XI0/XI63/XI6/NET33_XI0/XI63/XI6/MM4_d
+ N_XI0/XI63/XI6/NET34_XI0/XI63/XI6/MM4_g N_VDD_XI0/XI63/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI6/MM10 N_XI0/XI63/XI6/NET35_XI0/XI63/XI6/MM10_d
+ N_XI0/XI63/XI6/NET36_XI0/XI63/XI6/MM10_g N_VDD_XI0/XI63/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI6/MM11 N_XI0/XI63/XI6/NET36_XI0/XI63/XI6/MM11_d
+ N_XI0/XI63/XI6/NET35_XI0/XI63/XI6/MM11_g N_VDD_XI0/XI63/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI7/MM2 N_XI0/XI63/XI7/NET34_XI0/XI63/XI7/MM2_d
+ N_XI0/XI63/XI7/NET33_XI0/XI63/XI7/MM2_g N_VSS_XI0/XI63/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM3 N_XI0/XI63/XI7/NET33_XI0/XI63/XI7/MM3_d
+ N_WL<122>_XI0/XI63/XI7/MM3_g N_BLN<8>_XI0/XI63/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM0 N_XI0/XI63/XI7/NET34_XI0/XI63/XI7/MM0_d
+ N_WL<122>_XI0/XI63/XI7/MM0_g N_BL<8>_XI0/XI63/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM1 N_XI0/XI63/XI7/NET33_XI0/XI63/XI7/MM1_d
+ N_XI0/XI63/XI7/NET34_XI0/XI63/XI7/MM1_g N_VSS_XI0/XI63/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM9 N_XI0/XI63/XI7/NET36_XI0/XI63/XI7/MM9_d
+ N_WL<123>_XI0/XI63/XI7/MM9_g N_BL<8>_XI0/XI63/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM6 N_XI0/XI63/XI7/NET35_XI0/XI63/XI7/MM6_d
+ N_XI0/XI63/XI7/NET36_XI0/XI63/XI7/MM6_g N_VSS_XI0/XI63/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM7 N_XI0/XI63/XI7/NET36_XI0/XI63/XI7/MM7_d
+ N_XI0/XI63/XI7/NET35_XI0/XI63/XI7/MM7_g N_VSS_XI0/XI63/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM8 N_XI0/XI63/XI7/NET35_XI0/XI63/XI7/MM8_d
+ N_WL<123>_XI0/XI63/XI7/MM8_g N_BLN<8>_XI0/XI63/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI7/MM5 N_XI0/XI63/XI7/NET34_XI0/XI63/XI7/MM5_d
+ N_XI0/XI63/XI7/NET33_XI0/XI63/XI7/MM5_g N_VDD_XI0/XI63/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI7/MM4 N_XI0/XI63/XI7/NET33_XI0/XI63/XI7/MM4_d
+ N_XI0/XI63/XI7/NET34_XI0/XI63/XI7/MM4_g N_VDD_XI0/XI63/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI7/MM10 N_XI0/XI63/XI7/NET35_XI0/XI63/XI7/MM10_d
+ N_XI0/XI63/XI7/NET36_XI0/XI63/XI7/MM10_g N_VDD_XI0/XI63/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI7/MM11 N_XI0/XI63/XI7/NET36_XI0/XI63/XI7/MM11_d
+ N_XI0/XI63/XI7/NET35_XI0/XI63/XI7/MM11_g N_VDD_XI0/XI63/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI8/MM2 N_XI0/XI63/XI8/NET34_XI0/XI63/XI8/MM2_d
+ N_XI0/XI63/XI8/NET33_XI0/XI63/XI8/MM2_g N_VSS_XI0/XI63/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM3 N_XI0/XI63/XI8/NET33_XI0/XI63/XI8/MM3_d
+ N_WL<122>_XI0/XI63/XI8/MM3_g N_BLN<7>_XI0/XI63/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM0 N_XI0/XI63/XI8/NET34_XI0/XI63/XI8/MM0_d
+ N_WL<122>_XI0/XI63/XI8/MM0_g N_BL<7>_XI0/XI63/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM1 N_XI0/XI63/XI8/NET33_XI0/XI63/XI8/MM1_d
+ N_XI0/XI63/XI8/NET34_XI0/XI63/XI8/MM1_g N_VSS_XI0/XI63/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM9 N_XI0/XI63/XI8/NET36_XI0/XI63/XI8/MM9_d
+ N_WL<123>_XI0/XI63/XI8/MM9_g N_BL<7>_XI0/XI63/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM6 N_XI0/XI63/XI8/NET35_XI0/XI63/XI8/MM6_d
+ N_XI0/XI63/XI8/NET36_XI0/XI63/XI8/MM6_g N_VSS_XI0/XI63/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM7 N_XI0/XI63/XI8/NET36_XI0/XI63/XI8/MM7_d
+ N_XI0/XI63/XI8/NET35_XI0/XI63/XI8/MM7_g N_VSS_XI0/XI63/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM8 N_XI0/XI63/XI8/NET35_XI0/XI63/XI8/MM8_d
+ N_WL<123>_XI0/XI63/XI8/MM8_g N_BLN<7>_XI0/XI63/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI8/MM5 N_XI0/XI63/XI8/NET34_XI0/XI63/XI8/MM5_d
+ N_XI0/XI63/XI8/NET33_XI0/XI63/XI8/MM5_g N_VDD_XI0/XI63/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI8/MM4 N_XI0/XI63/XI8/NET33_XI0/XI63/XI8/MM4_d
+ N_XI0/XI63/XI8/NET34_XI0/XI63/XI8/MM4_g N_VDD_XI0/XI63/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI8/MM10 N_XI0/XI63/XI8/NET35_XI0/XI63/XI8/MM10_d
+ N_XI0/XI63/XI8/NET36_XI0/XI63/XI8/MM10_g N_VDD_XI0/XI63/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI8/MM11 N_XI0/XI63/XI8/NET36_XI0/XI63/XI8/MM11_d
+ N_XI0/XI63/XI8/NET35_XI0/XI63/XI8/MM11_g N_VDD_XI0/XI63/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI9/MM2 N_XI0/XI63/XI9/NET34_XI0/XI63/XI9/MM2_d
+ N_XI0/XI63/XI9/NET33_XI0/XI63/XI9/MM2_g N_VSS_XI0/XI63/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM3 N_XI0/XI63/XI9/NET33_XI0/XI63/XI9/MM3_d
+ N_WL<122>_XI0/XI63/XI9/MM3_g N_BLN<6>_XI0/XI63/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM0 N_XI0/XI63/XI9/NET34_XI0/XI63/XI9/MM0_d
+ N_WL<122>_XI0/XI63/XI9/MM0_g N_BL<6>_XI0/XI63/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM1 N_XI0/XI63/XI9/NET33_XI0/XI63/XI9/MM1_d
+ N_XI0/XI63/XI9/NET34_XI0/XI63/XI9/MM1_g N_VSS_XI0/XI63/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM9 N_XI0/XI63/XI9/NET36_XI0/XI63/XI9/MM9_d
+ N_WL<123>_XI0/XI63/XI9/MM9_g N_BL<6>_XI0/XI63/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM6 N_XI0/XI63/XI9/NET35_XI0/XI63/XI9/MM6_d
+ N_XI0/XI63/XI9/NET36_XI0/XI63/XI9/MM6_g N_VSS_XI0/XI63/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM7 N_XI0/XI63/XI9/NET36_XI0/XI63/XI9/MM7_d
+ N_XI0/XI63/XI9/NET35_XI0/XI63/XI9/MM7_g N_VSS_XI0/XI63/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM8 N_XI0/XI63/XI9/NET35_XI0/XI63/XI9/MM8_d
+ N_WL<123>_XI0/XI63/XI9/MM8_g N_BLN<6>_XI0/XI63/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI9/MM5 N_XI0/XI63/XI9/NET34_XI0/XI63/XI9/MM5_d
+ N_XI0/XI63/XI9/NET33_XI0/XI63/XI9/MM5_g N_VDD_XI0/XI63/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI9/MM4 N_XI0/XI63/XI9/NET33_XI0/XI63/XI9/MM4_d
+ N_XI0/XI63/XI9/NET34_XI0/XI63/XI9/MM4_g N_VDD_XI0/XI63/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI9/MM10 N_XI0/XI63/XI9/NET35_XI0/XI63/XI9/MM10_d
+ N_XI0/XI63/XI9/NET36_XI0/XI63/XI9/MM10_g N_VDD_XI0/XI63/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI9/MM11 N_XI0/XI63/XI9/NET36_XI0/XI63/XI9/MM11_d
+ N_XI0/XI63/XI9/NET35_XI0/XI63/XI9/MM11_g N_VDD_XI0/XI63/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI10/MM2 N_XI0/XI63/XI10/NET34_XI0/XI63/XI10/MM2_d
+ N_XI0/XI63/XI10/NET33_XI0/XI63/XI10/MM2_g N_VSS_XI0/XI63/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM3 N_XI0/XI63/XI10/NET33_XI0/XI63/XI10/MM3_d
+ N_WL<122>_XI0/XI63/XI10/MM3_g N_BLN<5>_XI0/XI63/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM0 N_XI0/XI63/XI10/NET34_XI0/XI63/XI10/MM0_d
+ N_WL<122>_XI0/XI63/XI10/MM0_g N_BL<5>_XI0/XI63/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM1 N_XI0/XI63/XI10/NET33_XI0/XI63/XI10/MM1_d
+ N_XI0/XI63/XI10/NET34_XI0/XI63/XI10/MM1_g N_VSS_XI0/XI63/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM9 N_XI0/XI63/XI10/NET36_XI0/XI63/XI10/MM9_d
+ N_WL<123>_XI0/XI63/XI10/MM9_g N_BL<5>_XI0/XI63/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM6 N_XI0/XI63/XI10/NET35_XI0/XI63/XI10/MM6_d
+ N_XI0/XI63/XI10/NET36_XI0/XI63/XI10/MM6_g N_VSS_XI0/XI63/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM7 N_XI0/XI63/XI10/NET36_XI0/XI63/XI10/MM7_d
+ N_XI0/XI63/XI10/NET35_XI0/XI63/XI10/MM7_g N_VSS_XI0/XI63/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM8 N_XI0/XI63/XI10/NET35_XI0/XI63/XI10/MM8_d
+ N_WL<123>_XI0/XI63/XI10/MM8_g N_BLN<5>_XI0/XI63/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI10/MM5 N_XI0/XI63/XI10/NET34_XI0/XI63/XI10/MM5_d
+ N_XI0/XI63/XI10/NET33_XI0/XI63/XI10/MM5_g N_VDD_XI0/XI63/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI10/MM4 N_XI0/XI63/XI10/NET33_XI0/XI63/XI10/MM4_d
+ N_XI0/XI63/XI10/NET34_XI0/XI63/XI10/MM4_g N_VDD_XI0/XI63/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI10/MM10 N_XI0/XI63/XI10/NET35_XI0/XI63/XI10/MM10_d
+ N_XI0/XI63/XI10/NET36_XI0/XI63/XI10/MM10_g N_VDD_XI0/XI63/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI10/MM11 N_XI0/XI63/XI10/NET36_XI0/XI63/XI10/MM11_d
+ N_XI0/XI63/XI10/NET35_XI0/XI63/XI10/MM11_g N_VDD_XI0/XI63/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI11/MM2 N_XI0/XI63/XI11/NET34_XI0/XI63/XI11/MM2_d
+ N_XI0/XI63/XI11/NET33_XI0/XI63/XI11/MM2_g N_VSS_XI0/XI63/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM3 N_XI0/XI63/XI11/NET33_XI0/XI63/XI11/MM3_d
+ N_WL<122>_XI0/XI63/XI11/MM3_g N_BLN<4>_XI0/XI63/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM0 N_XI0/XI63/XI11/NET34_XI0/XI63/XI11/MM0_d
+ N_WL<122>_XI0/XI63/XI11/MM0_g N_BL<4>_XI0/XI63/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM1 N_XI0/XI63/XI11/NET33_XI0/XI63/XI11/MM1_d
+ N_XI0/XI63/XI11/NET34_XI0/XI63/XI11/MM1_g N_VSS_XI0/XI63/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM9 N_XI0/XI63/XI11/NET36_XI0/XI63/XI11/MM9_d
+ N_WL<123>_XI0/XI63/XI11/MM9_g N_BL<4>_XI0/XI63/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM6 N_XI0/XI63/XI11/NET35_XI0/XI63/XI11/MM6_d
+ N_XI0/XI63/XI11/NET36_XI0/XI63/XI11/MM6_g N_VSS_XI0/XI63/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM7 N_XI0/XI63/XI11/NET36_XI0/XI63/XI11/MM7_d
+ N_XI0/XI63/XI11/NET35_XI0/XI63/XI11/MM7_g N_VSS_XI0/XI63/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM8 N_XI0/XI63/XI11/NET35_XI0/XI63/XI11/MM8_d
+ N_WL<123>_XI0/XI63/XI11/MM8_g N_BLN<4>_XI0/XI63/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI11/MM5 N_XI0/XI63/XI11/NET34_XI0/XI63/XI11/MM5_d
+ N_XI0/XI63/XI11/NET33_XI0/XI63/XI11/MM5_g N_VDD_XI0/XI63/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI11/MM4 N_XI0/XI63/XI11/NET33_XI0/XI63/XI11/MM4_d
+ N_XI0/XI63/XI11/NET34_XI0/XI63/XI11/MM4_g N_VDD_XI0/XI63/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI11/MM10 N_XI0/XI63/XI11/NET35_XI0/XI63/XI11/MM10_d
+ N_XI0/XI63/XI11/NET36_XI0/XI63/XI11/MM10_g N_VDD_XI0/XI63/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI11/MM11 N_XI0/XI63/XI11/NET36_XI0/XI63/XI11/MM11_d
+ N_XI0/XI63/XI11/NET35_XI0/XI63/XI11/MM11_g N_VDD_XI0/XI63/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI12/MM2 N_XI0/XI63/XI12/NET34_XI0/XI63/XI12/MM2_d
+ N_XI0/XI63/XI12/NET33_XI0/XI63/XI12/MM2_g N_VSS_XI0/XI63/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM3 N_XI0/XI63/XI12/NET33_XI0/XI63/XI12/MM3_d
+ N_WL<122>_XI0/XI63/XI12/MM3_g N_BLN<3>_XI0/XI63/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM0 N_XI0/XI63/XI12/NET34_XI0/XI63/XI12/MM0_d
+ N_WL<122>_XI0/XI63/XI12/MM0_g N_BL<3>_XI0/XI63/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM1 N_XI0/XI63/XI12/NET33_XI0/XI63/XI12/MM1_d
+ N_XI0/XI63/XI12/NET34_XI0/XI63/XI12/MM1_g N_VSS_XI0/XI63/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM9 N_XI0/XI63/XI12/NET36_XI0/XI63/XI12/MM9_d
+ N_WL<123>_XI0/XI63/XI12/MM9_g N_BL<3>_XI0/XI63/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM6 N_XI0/XI63/XI12/NET35_XI0/XI63/XI12/MM6_d
+ N_XI0/XI63/XI12/NET36_XI0/XI63/XI12/MM6_g N_VSS_XI0/XI63/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM7 N_XI0/XI63/XI12/NET36_XI0/XI63/XI12/MM7_d
+ N_XI0/XI63/XI12/NET35_XI0/XI63/XI12/MM7_g N_VSS_XI0/XI63/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM8 N_XI0/XI63/XI12/NET35_XI0/XI63/XI12/MM8_d
+ N_WL<123>_XI0/XI63/XI12/MM8_g N_BLN<3>_XI0/XI63/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI12/MM5 N_XI0/XI63/XI12/NET34_XI0/XI63/XI12/MM5_d
+ N_XI0/XI63/XI12/NET33_XI0/XI63/XI12/MM5_g N_VDD_XI0/XI63/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI12/MM4 N_XI0/XI63/XI12/NET33_XI0/XI63/XI12/MM4_d
+ N_XI0/XI63/XI12/NET34_XI0/XI63/XI12/MM4_g N_VDD_XI0/XI63/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI12/MM10 N_XI0/XI63/XI12/NET35_XI0/XI63/XI12/MM10_d
+ N_XI0/XI63/XI12/NET36_XI0/XI63/XI12/MM10_g N_VDD_XI0/XI63/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI12/MM11 N_XI0/XI63/XI12/NET36_XI0/XI63/XI12/MM11_d
+ N_XI0/XI63/XI12/NET35_XI0/XI63/XI12/MM11_g N_VDD_XI0/XI63/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI13/MM2 N_XI0/XI63/XI13/NET34_XI0/XI63/XI13/MM2_d
+ N_XI0/XI63/XI13/NET33_XI0/XI63/XI13/MM2_g N_VSS_XI0/XI63/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM3 N_XI0/XI63/XI13/NET33_XI0/XI63/XI13/MM3_d
+ N_WL<122>_XI0/XI63/XI13/MM3_g N_BLN<2>_XI0/XI63/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM0 N_XI0/XI63/XI13/NET34_XI0/XI63/XI13/MM0_d
+ N_WL<122>_XI0/XI63/XI13/MM0_g N_BL<2>_XI0/XI63/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM1 N_XI0/XI63/XI13/NET33_XI0/XI63/XI13/MM1_d
+ N_XI0/XI63/XI13/NET34_XI0/XI63/XI13/MM1_g N_VSS_XI0/XI63/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM9 N_XI0/XI63/XI13/NET36_XI0/XI63/XI13/MM9_d
+ N_WL<123>_XI0/XI63/XI13/MM9_g N_BL<2>_XI0/XI63/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM6 N_XI0/XI63/XI13/NET35_XI0/XI63/XI13/MM6_d
+ N_XI0/XI63/XI13/NET36_XI0/XI63/XI13/MM6_g N_VSS_XI0/XI63/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM7 N_XI0/XI63/XI13/NET36_XI0/XI63/XI13/MM7_d
+ N_XI0/XI63/XI13/NET35_XI0/XI63/XI13/MM7_g N_VSS_XI0/XI63/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM8 N_XI0/XI63/XI13/NET35_XI0/XI63/XI13/MM8_d
+ N_WL<123>_XI0/XI63/XI13/MM8_g N_BLN<2>_XI0/XI63/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI13/MM5 N_XI0/XI63/XI13/NET34_XI0/XI63/XI13/MM5_d
+ N_XI0/XI63/XI13/NET33_XI0/XI63/XI13/MM5_g N_VDD_XI0/XI63/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI13/MM4 N_XI0/XI63/XI13/NET33_XI0/XI63/XI13/MM4_d
+ N_XI0/XI63/XI13/NET34_XI0/XI63/XI13/MM4_g N_VDD_XI0/XI63/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI13/MM10 N_XI0/XI63/XI13/NET35_XI0/XI63/XI13/MM10_d
+ N_XI0/XI63/XI13/NET36_XI0/XI63/XI13/MM10_g N_VDD_XI0/XI63/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI13/MM11 N_XI0/XI63/XI13/NET36_XI0/XI63/XI13/MM11_d
+ N_XI0/XI63/XI13/NET35_XI0/XI63/XI13/MM11_g N_VDD_XI0/XI63/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI14/MM2 N_XI0/XI63/XI14/NET34_XI0/XI63/XI14/MM2_d
+ N_XI0/XI63/XI14/NET33_XI0/XI63/XI14/MM2_g N_VSS_XI0/XI63/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM3 N_XI0/XI63/XI14/NET33_XI0/XI63/XI14/MM3_d
+ N_WL<122>_XI0/XI63/XI14/MM3_g N_BLN<1>_XI0/XI63/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM0 N_XI0/XI63/XI14/NET34_XI0/XI63/XI14/MM0_d
+ N_WL<122>_XI0/XI63/XI14/MM0_g N_BL<1>_XI0/XI63/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM1 N_XI0/XI63/XI14/NET33_XI0/XI63/XI14/MM1_d
+ N_XI0/XI63/XI14/NET34_XI0/XI63/XI14/MM1_g N_VSS_XI0/XI63/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM9 N_XI0/XI63/XI14/NET36_XI0/XI63/XI14/MM9_d
+ N_WL<123>_XI0/XI63/XI14/MM9_g N_BL<1>_XI0/XI63/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM6 N_XI0/XI63/XI14/NET35_XI0/XI63/XI14/MM6_d
+ N_XI0/XI63/XI14/NET36_XI0/XI63/XI14/MM6_g N_VSS_XI0/XI63/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM7 N_XI0/XI63/XI14/NET36_XI0/XI63/XI14/MM7_d
+ N_XI0/XI63/XI14/NET35_XI0/XI63/XI14/MM7_g N_VSS_XI0/XI63/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM8 N_XI0/XI63/XI14/NET35_XI0/XI63/XI14/MM8_d
+ N_WL<123>_XI0/XI63/XI14/MM8_g N_BLN<1>_XI0/XI63/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI14/MM5 N_XI0/XI63/XI14/NET34_XI0/XI63/XI14/MM5_d
+ N_XI0/XI63/XI14/NET33_XI0/XI63/XI14/MM5_g N_VDD_XI0/XI63/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI14/MM4 N_XI0/XI63/XI14/NET33_XI0/XI63/XI14/MM4_d
+ N_XI0/XI63/XI14/NET34_XI0/XI63/XI14/MM4_g N_VDD_XI0/XI63/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI14/MM10 N_XI0/XI63/XI14/NET35_XI0/XI63/XI14/MM10_d
+ N_XI0/XI63/XI14/NET36_XI0/XI63/XI14/MM10_g N_VDD_XI0/XI63/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI14/MM11 N_XI0/XI63/XI14/NET36_XI0/XI63/XI14/MM11_d
+ N_XI0/XI63/XI14/NET35_XI0/XI63/XI14/MM11_g N_VDD_XI0/XI63/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI15/MM2 N_XI0/XI63/XI15/NET34_XI0/XI63/XI15/MM2_d
+ N_XI0/XI63/XI15/NET33_XI0/XI63/XI15/MM2_g N_VSS_XI0/XI63/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM3 N_XI0/XI63/XI15/NET33_XI0/XI63/XI15/MM3_d
+ N_WL<122>_XI0/XI63/XI15/MM3_g N_BLN<0>_XI0/XI63/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM0 N_XI0/XI63/XI15/NET34_XI0/XI63/XI15/MM0_d
+ N_WL<122>_XI0/XI63/XI15/MM0_g N_BL<0>_XI0/XI63/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM1 N_XI0/XI63/XI15/NET33_XI0/XI63/XI15/MM1_d
+ N_XI0/XI63/XI15/NET34_XI0/XI63/XI15/MM1_g N_VSS_XI0/XI63/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM9 N_XI0/XI63/XI15/NET36_XI0/XI63/XI15/MM9_d
+ N_WL<123>_XI0/XI63/XI15/MM9_g N_BL<0>_XI0/XI63/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM6 N_XI0/XI63/XI15/NET35_XI0/XI63/XI15/MM6_d
+ N_XI0/XI63/XI15/NET36_XI0/XI63/XI15/MM6_g N_VSS_XI0/XI63/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM7 N_XI0/XI63/XI15/NET36_XI0/XI63/XI15/MM7_d
+ N_XI0/XI63/XI15/NET35_XI0/XI63/XI15/MM7_g N_VSS_XI0/XI63/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM8 N_XI0/XI63/XI15/NET35_XI0/XI63/XI15/MM8_d
+ N_WL<123>_XI0/XI63/XI15/MM8_g N_BLN<0>_XI0/XI63/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI63/XI15/MM5 N_XI0/XI63/XI15/NET34_XI0/XI63/XI15/MM5_d
+ N_XI0/XI63/XI15/NET33_XI0/XI63/XI15/MM5_g N_VDD_XI0/XI63/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI15/MM4 N_XI0/XI63/XI15/NET33_XI0/XI63/XI15/MM4_d
+ N_XI0/XI63/XI15/NET34_XI0/XI63/XI15/MM4_g N_VDD_XI0/XI63/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI15/MM10 N_XI0/XI63/XI15/NET35_XI0/XI63/XI15/MM10_d
+ N_XI0/XI63/XI15/NET36_XI0/XI63/XI15/MM10_g N_VDD_XI0/XI63/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI63/XI15/MM11 N_XI0/XI63/XI15/NET36_XI0/XI63/XI15/MM11_d
+ N_XI0/XI63/XI15/NET35_XI0/XI63/XI15/MM11_g N_VDD_XI0/XI63/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI0/MM2 N_XI0/XI64/XI0/NET34_XI0/XI64/XI0/MM2_d
+ N_XI0/XI64/XI0/NET33_XI0/XI64/XI0/MM2_g N_VSS_XI0/XI64/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM3 N_XI0/XI64/XI0/NET33_XI0/XI64/XI0/MM3_d
+ N_WL<124>_XI0/XI64/XI0/MM3_g N_BLN<15>_XI0/XI64/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM0 N_XI0/XI64/XI0/NET34_XI0/XI64/XI0/MM0_d
+ N_WL<124>_XI0/XI64/XI0/MM0_g N_BL<15>_XI0/XI64/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM1 N_XI0/XI64/XI0/NET33_XI0/XI64/XI0/MM1_d
+ N_XI0/XI64/XI0/NET34_XI0/XI64/XI0/MM1_g N_VSS_XI0/XI64/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM9 N_XI0/XI64/XI0/NET36_XI0/XI64/XI0/MM9_d
+ N_WL<125>_XI0/XI64/XI0/MM9_g N_BL<15>_XI0/XI64/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM6 N_XI0/XI64/XI0/NET35_XI0/XI64/XI0/MM6_d
+ N_XI0/XI64/XI0/NET36_XI0/XI64/XI0/MM6_g N_VSS_XI0/XI64/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM7 N_XI0/XI64/XI0/NET36_XI0/XI64/XI0/MM7_d
+ N_XI0/XI64/XI0/NET35_XI0/XI64/XI0/MM7_g N_VSS_XI0/XI64/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM8 N_XI0/XI64/XI0/NET35_XI0/XI64/XI0/MM8_d
+ N_WL<125>_XI0/XI64/XI0/MM8_g N_BLN<15>_XI0/XI64/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI0/MM5 N_XI0/XI64/XI0/NET34_XI0/XI64/XI0/MM5_d
+ N_XI0/XI64/XI0/NET33_XI0/XI64/XI0/MM5_g N_VDD_XI0/XI64/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI0/MM4 N_XI0/XI64/XI0/NET33_XI0/XI64/XI0/MM4_d
+ N_XI0/XI64/XI0/NET34_XI0/XI64/XI0/MM4_g N_VDD_XI0/XI64/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI0/MM10 N_XI0/XI64/XI0/NET35_XI0/XI64/XI0/MM10_d
+ N_XI0/XI64/XI0/NET36_XI0/XI64/XI0/MM10_g N_VDD_XI0/XI64/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI0/MM11 N_XI0/XI64/XI0/NET36_XI0/XI64/XI0/MM11_d
+ N_XI0/XI64/XI0/NET35_XI0/XI64/XI0/MM11_g N_VDD_XI0/XI64/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI1/MM2 N_XI0/XI64/XI1/NET34_XI0/XI64/XI1/MM2_d
+ N_XI0/XI64/XI1/NET33_XI0/XI64/XI1/MM2_g N_VSS_XI0/XI64/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM3 N_XI0/XI64/XI1/NET33_XI0/XI64/XI1/MM3_d
+ N_WL<124>_XI0/XI64/XI1/MM3_g N_BLN<14>_XI0/XI64/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM0 N_XI0/XI64/XI1/NET34_XI0/XI64/XI1/MM0_d
+ N_WL<124>_XI0/XI64/XI1/MM0_g N_BL<14>_XI0/XI64/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM1 N_XI0/XI64/XI1/NET33_XI0/XI64/XI1/MM1_d
+ N_XI0/XI64/XI1/NET34_XI0/XI64/XI1/MM1_g N_VSS_XI0/XI64/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM9 N_XI0/XI64/XI1/NET36_XI0/XI64/XI1/MM9_d
+ N_WL<125>_XI0/XI64/XI1/MM9_g N_BL<14>_XI0/XI64/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM6 N_XI0/XI64/XI1/NET35_XI0/XI64/XI1/MM6_d
+ N_XI0/XI64/XI1/NET36_XI0/XI64/XI1/MM6_g N_VSS_XI0/XI64/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM7 N_XI0/XI64/XI1/NET36_XI0/XI64/XI1/MM7_d
+ N_XI0/XI64/XI1/NET35_XI0/XI64/XI1/MM7_g N_VSS_XI0/XI64/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM8 N_XI0/XI64/XI1/NET35_XI0/XI64/XI1/MM8_d
+ N_WL<125>_XI0/XI64/XI1/MM8_g N_BLN<14>_XI0/XI64/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI1/MM5 N_XI0/XI64/XI1/NET34_XI0/XI64/XI1/MM5_d
+ N_XI0/XI64/XI1/NET33_XI0/XI64/XI1/MM5_g N_VDD_XI0/XI64/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI1/MM4 N_XI0/XI64/XI1/NET33_XI0/XI64/XI1/MM4_d
+ N_XI0/XI64/XI1/NET34_XI0/XI64/XI1/MM4_g N_VDD_XI0/XI64/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI1/MM10 N_XI0/XI64/XI1/NET35_XI0/XI64/XI1/MM10_d
+ N_XI0/XI64/XI1/NET36_XI0/XI64/XI1/MM10_g N_VDD_XI0/XI64/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI1/MM11 N_XI0/XI64/XI1/NET36_XI0/XI64/XI1/MM11_d
+ N_XI0/XI64/XI1/NET35_XI0/XI64/XI1/MM11_g N_VDD_XI0/XI64/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI2/MM2 N_XI0/XI64/XI2/NET34_XI0/XI64/XI2/MM2_d
+ N_XI0/XI64/XI2/NET33_XI0/XI64/XI2/MM2_g N_VSS_XI0/XI64/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM3 N_XI0/XI64/XI2/NET33_XI0/XI64/XI2/MM3_d
+ N_WL<124>_XI0/XI64/XI2/MM3_g N_BLN<13>_XI0/XI64/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM0 N_XI0/XI64/XI2/NET34_XI0/XI64/XI2/MM0_d
+ N_WL<124>_XI0/XI64/XI2/MM0_g N_BL<13>_XI0/XI64/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM1 N_XI0/XI64/XI2/NET33_XI0/XI64/XI2/MM1_d
+ N_XI0/XI64/XI2/NET34_XI0/XI64/XI2/MM1_g N_VSS_XI0/XI64/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM9 N_XI0/XI64/XI2/NET36_XI0/XI64/XI2/MM9_d
+ N_WL<125>_XI0/XI64/XI2/MM9_g N_BL<13>_XI0/XI64/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM6 N_XI0/XI64/XI2/NET35_XI0/XI64/XI2/MM6_d
+ N_XI0/XI64/XI2/NET36_XI0/XI64/XI2/MM6_g N_VSS_XI0/XI64/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM7 N_XI0/XI64/XI2/NET36_XI0/XI64/XI2/MM7_d
+ N_XI0/XI64/XI2/NET35_XI0/XI64/XI2/MM7_g N_VSS_XI0/XI64/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM8 N_XI0/XI64/XI2/NET35_XI0/XI64/XI2/MM8_d
+ N_WL<125>_XI0/XI64/XI2/MM8_g N_BLN<13>_XI0/XI64/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI2/MM5 N_XI0/XI64/XI2/NET34_XI0/XI64/XI2/MM5_d
+ N_XI0/XI64/XI2/NET33_XI0/XI64/XI2/MM5_g N_VDD_XI0/XI64/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI2/MM4 N_XI0/XI64/XI2/NET33_XI0/XI64/XI2/MM4_d
+ N_XI0/XI64/XI2/NET34_XI0/XI64/XI2/MM4_g N_VDD_XI0/XI64/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI2/MM10 N_XI0/XI64/XI2/NET35_XI0/XI64/XI2/MM10_d
+ N_XI0/XI64/XI2/NET36_XI0/XI64/XI2/MM10_g N_VDD_XI0/XI64/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI2/MM11 N_XI0/XI64/XI2/NET36_XI0/XI64/XI2/MM11_d
+ N_XI0/XI64/XI2/NET35_XI0/XI64/XI2/MM11_g N_VDD_XI0/XI64/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI3/MM2 N_XI0/XI64/XI3/NET34_XI0/XI64/XI3/MM2_d
+ N_XI0/XI64/XI3/NET33_XI0/XI64/XI3/MM2_g N_VSS_XI0/XI64/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM3 N_XI0/XI64/XI3/NET33_XI0/XI64/XI3/MM3_d
+ N_WL<124>_XI0/XI64/XI3/MM3_g N_BLN<12>_XI0/XI64/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM0 N_XI0/XI64/XI3/NET34_XI0/XI64/XI3/MM0_d
+ N_WL<124>_XI0/XI64/XI3/MM0_g N_BL<12>_XI0/XI64/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM1 N_XI0/XI64/XI3/NET33_XI0/XI64/XI3/MM1_d
+ N_XI0/XI64/XI3/NET34_XI0/XI64/XI3/MM1_g N_VSS_XI0/XI64/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM9 N_XI0/XI64/XI3/NET36_XI0/XI64/XI3/MM9_d
+ N_WL<125>_XI0/XI64/XI3/MM9_g N_BL<12>_XI0/XI64/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM6 N_XI0/XI64/XI3/NET35_XI0/XI64/XI3/MM6_d
+ N_XI0/XI64/XI3/NET36_XI0/XI64/XI3/MM6_g N_VSS_XI0/XI64/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM7 N_XI0/XI64/XI3/NET36_XI0/XI64/XI3/MM7_d
+ N_XI0/XI64/XI3/NET35_XI0/XI64/XI3/MM7_g N_VSS_XI0/XI64/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM8 N_XI0/XI64/XI3/NET35_XI0/XI64/XI3/MM8_d
+ N_WL<125>_XI0/XI64/XI3/MM8_g N_BLN<12>_XI0/XI64/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI3/MM5 N_XI0/XI64/XI3/NET34_XI0/XI64/XI3/MM5_d
+ N_XI0/XI64/XI3/NET33_XI0/XI64/XI3/MM5_g N_VDD_XI0/XI64/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI3/MM4 N_XI0/XI64/XI3/NET33_XI0/XI64/XI3/MM4_d
+ N_XI0/XI64/XI3/NET34_XI0/XI64/XI3/MM4_g N_VDD_XI0/XI64/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI3/MM10 N_XI0/XI64/XI3/NET35_XI0/XI64/XI3/MM10_d
+ N_XI0/XI64/XI3/NET36_XI0/XI64/XI3/MM10_g N_VDD_XI0/XI64/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI3/MM11 N_XI0/XI64/XI3/NET36_XI0/XI64/XI3/MM11_d
+ N_XI0/XI64/XI3/NET35_XI0/XI64/XI3/MM11_g N_VDD_XI0/XI64/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI4/MM2 N_XI0/XI64/XI4/NET34_XI0/XI64/XI4/MM2_d
+ N_XI0/XI64/XI4/NET33_XI0/XI64/XI4/MM2_g N_VSS_XI0/XI64/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM3 N_XI0/XI64/XI4/NET33_XI0/XI64/XI4/MM3_d
+ N_WL<124>_XI0/XI64/XI4/MM3_g N_BLN<11>_XI0/XI64/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM0 N_XI0/XI64/XI4/NET34_XI0/XI64/XI4/MM0_d
+ N_WL<124>_XI0/XI64/XI4/MM0_g N_BL<11>_XI0/XI64/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM1 N_XI0/XI64/XI4/NET33_XI0/XI64/XI4/MM1_d
+ N_XI0/XI64/XI4/NET34_XI0/XI64/XI4/MM1_g N_VSS_XI0/XI64/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM9 N_XI0/XI64/XI4/NET36_XI0/XI64/XI4/MM9_d
+ N_WL<125>_XI0/XI64/XI4/MM9_g N_BL<11>_XI0/XI64/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM6 N_XI0/XI64/XI4/NET35_XI0/XI64/XI4/MM6_d
+ N_XI0/XI64/XI4/NET36_XI0/XI64/XI4/MM6_g N_VSS_XI0/XI64/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM7 N_XI0/XI64/XI4/NET36_XI0/XI64/XI4/MM7_d
+ N_XI0/XI64/XI4/NET35_XI0/XI64/XI4/MM7_g N_VSS_XI0/XI64/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM8 N_XI0/XI64/XI4/NET35_XI0/XI64/XI4/MM8_d
+ N_WL<125>_XI0/XI64/XI4/MM8_g N_BLN<11>_XI0/XI64/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI4/MM5 N_XI0/XI64/XI4/NET34_XI0/XI64/XI4/MM5_d
+ N_XI0/XI64/XI4/NET33_XI0/XI64/XI4/MM5_g N_VDD_XI0/XI64/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI4/MM4 N_XI0/XI64/XI4/NET33_XI0/XI64/XI4/MM4_d
+ N_XI0/XI64/XI4/NET34_XI0/XI64/XI4/MM4_g N_VDD_XI0/XI64/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI4/MM10 N_XI0/XI64/XI4/NET35_XI0/XI64/XI4/MM10_d
+ N_XI0/XI64/XI4/NET36_XI0/XI64/XI4/MM10_g N_VDD_XI0/XI64/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI4/MM11 N_XI0/XI64/XI4/NET36_XI0/XI64/XI4/MM11_d
+ N_XI0/XI64/XI4/NET35_XI0/XI64/XI4/MM11_g N_VDD_XI0/XI64/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI5/MM2 N_XI0/XI64/XI5/NET34_XI0/XI64/XI5/MM2_d
+ N_XI0/XI64/XI5/NET33_XI0/XI64/XI5/MM2_g N_VSS_XI0/XI64/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM3 N_XI0/XI64/XI5/NET33_XI0/XI64/XI5/MM3_d
+ N_WL<124>_XI0/XI64/XI5/MM3_g N_BLN<10>_XI0/XI64/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM0 N_XI0/XI64/XI5/NET34_XI0/XI64/XI5/MM0_d
+ N_WL<124>_XI0/XI64/XI5/MM0_g N_BL<10>_XI0/XI64/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM1 N_XI0/XI64/XI5/NET33_XI0/XI64/XI5/MM1_d
+ N_XI0/XI64/XI5/NET34_XI0/XI64/XI5/MM1_g N_VSS_XI0/XI64/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM9 N_XI0/XI64/XI5/NET36_XI0/XI64/XI5/MM9_d
+ N_WL<125>_XI0/XI64/XI5/MM9_g N_BL<10>_XI0/XI64/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM6 N_XI0/XI64/XI5/NET35_XI0/XI64/XI5/MM6_d
+ N_XI0/XI64/XI5/NET36_XI0/XI64/XI5/MM6_g N_VSS_XI0/XI64/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM7 N_XI0/XI64/XI5/NET36_XI0/XI64/XI5/MM7_d
+ N_XI0/XI64/XI5/NET35_XI0/XI64/XI5/MM7_g N_VSS_XI0/XI64/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM8 N_XI0/XI64/XI5/NET35_XI0/XI64/XI5/MM8_d
+ N_WL<125>_XI0/XI64/XI5/MM8_g N_BLN<10>_XI0/XI64/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI5/MM5 N_XI0/XI64/XI5/NET34_XI0/XI64/XI5/MM5_d
+ N_XI0/XI64/XI5/NET33_XI0/XI64/XI5/MM5_g N_VDD_XI0/XI64/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI5/MM4 N_XI0/XI64/XI5/NET33_XI0/XI64/XI5/MM4_d
+ N_XI0/XI64/XI5/NET34_XI0/XI64/XI5/MM4_g N_VDD_XI0/XI64/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI5/MM10 N_XI0/XI64/XI5/NET35_XI0/XI64/XI5/MM10_d
+ N_XI0/XI64/XI5/NET36_XI0/XI64/XI5/MM10_g N_VDD_XI0/XI64/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI5/MM11 N_XI0/XI64/XI5/NET36_XI0/XI64/XI5/MM11_d
+ N_XI0/XI64/XI5/NET35_XI0/XI64/XI5/MM11_g N_VDD_XI0/XI64/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI6/MM2 N_XI0/XI64/XI6/NET34_XI0/XI64/XI6/MM2_d
+ N_XI0/XI64/XI6/NET33_XI0/XI64/XI6/MM2_g N_VSS_XI0/XI64/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM3 N_XI0/XI64/XI6/NET33_XI0/XI64/XI6/MM3_d
+ N_WL<124>_XI0/XI64/XI6/MM3_g N_BLN<9>_XI0/XI64/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM0 N_XI0/XI64/XI6/NET34_XI0/XI64/XI6/MM0_d
+ N_WL<124>_XI0/XI64/XI6/MM0_g N_BL<9>_XI0/XI64/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM1 N_XI0/XI64/XI6/NET33_XI0/XI64/XI6/MM1_d
+ N_XI0/XI64/XI6/NET34_XI0/XI64/XI6/MM1_g N_VSS_XI0/XI64/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM9 N_XI0/XI64/XI6/NET36_XI0/XI64/XI6/MM9_d
+ N_WL<125>_XI0/XI64/XI6/MM9_g N_BL<9>_XI0/XI64/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM6 N_XI0/XI64/XI6/NET35_XI0/XI64/XI6/MM6_d
+ N_XI0/XI64/XI6/NET36_XI0/XI64/XI6/MM6_g N_VSS_XI0/XI64/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM7 N_XI0/XI64/XI6/NET36_XI0/XI64/XI6/MM7_d
+ N_XI0/XI64/XI6/NET35_XI0/XI64/XI6/MM7_g N_VSS_XI0/XI64/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM8 N_XI0/XI64/XI6/NET35_XI0/XI64/XI6/MM8_d
+ N_WL<125>_XI0/XI64/XI6/MM8_g N_BLN<9>_XI0/XI64/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI6/MM5 N_XI0/XI64/XI6/NET34_XI0/XI64/XI6/MM5_d
+ N_XI0/XI64/XI6/NET33_XI0/XI64/XI6/MM5_g N_VDD_XI0/XI64/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI6/MM4 N_XI0/XI64/XI6/NET33_XI0/XI64/XI6/MM4_d
+ N_XI0/XI64/XI6/NET34_XI0/XI64/XI6/MM4_g N_VDD_XI0/XI64/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI6/MM10 N_XI0/XI64/XI6/NET35_XI0/XI64/XI6/MM10_d
+ N_XI0/XI64/XI6/NET36_XI0/XI64/XI6/MM10_g N_VDD_XI0/XI64/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI6/MM11 N_XI0/XI64/XI6/NET36_XI0/XI64/XI6/MM11_d
+ N_XI0/XI64/XI6/NET35_XI0/XI64/XI6/MM11_g N_VDD_XI0/XI64/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI7/MM2 N_XI0/XI64/XI7/NET34_XI0/XI64/XI7/MM2_d
+ N_XI0/XI64/XI7/NET33_XI0/XI64/XI7/MM2_g N_VSS_XI0/XI64/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM3 N_XI0/XI64/XI7/NET33_XI0/XI64/XI7/MM3_d
+ N_WL<124>_XI0/XI64/XI7/MM3_g N_BLN<8>_XI0/XI64/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM0 N_XI0/XI64/XI7/NET34_XI0/XI64/XI7/MM0_d
+ N_WL<124>_XI0/XI64/XI7/MM0_g N_BL<8>_XI0/XI64/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM1 N_XI0/XI64/XI7/NET33_XI0/XI64/XI7/MM1_d
+ N_XI0/XI64/XI7/NET34_XI0/XI64/XI7/MM1_g N_VSS_XI0/XI64/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM9 N_XI0/XI64/XI7/NET36_XI0/XI64/XI7/MM9_d
+ N_WL<125>_XI0/XI64/XI7/MM9_g N_BL<8>_XI0/XI64/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM6 N_XI0/XI64/XI7/NET35_XI0/XI64/XI7/MM6_d
+ N_XI0/XI64/XI7/NET36_XI0/XI64/XI7/MM6_g N_VSS_XI0/XI64/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM7 N_XI0/XI64/XI7/NET36_XI0/XI64/XI7/MM7_d
+ N_XI0/XI64/XI7/NET35_XI0/XI64/XI7/MM7_g N_VSS_XI0/XI64/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM8 N_XI0/XI64/XI7/NET35_XI0/XI64/XI7/MM8_d
+ N_WL<125>_XI0/XI64/XI7/MM8_g N_BLN<8>_XI0/XI64/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI7/MM5 N_XI0/XI64/XI7/NET34_XI0/XI64/XI7/MM5_d
+ N_XI0/XI64/XI7/NET33_XI0/XI64/XI7/MM5_g N_VDD_XI0/XI64/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI7/MM4 N_XI0/XI64/XI7/NET33_XI0/XI64/XI7/MM4_d
+ N_XI0/XI64/XI7/NET34_XI0/XI64/XI7/MM4_g N_VDD_XI0/XI64/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI7/MM10 N_XI0/XI64/XI7/NET35_XI0/XI64/XI7/MM10_d
+ N_XI0/XI64/XI7/NET36_XI0/XI64/XI7/MM10_g N_VDD_XI0/XI64/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI7/MM11 N_XI0/XI64/XI7/NET36_XI0/XI64/XI7/MM11_d
+ N_XI0/XI64/XI7/NET35_XI0/XI64/XI7/MM11_g N_VDD_XI0/XI64/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI8/MM2 N_XI0/XI64/XI8/NET34_XI0/XI64/XI8/MM2_d
+ N_XI0/XI64/XI8/NET33_XI0/XI64/XI8/MM2_g N_VSS_XI0/XI64/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM3 N_XI0/XI64/XI8/NET33_XI0/XI64/XI8/MM3_d
+ N_WL<124>_XI0/XI64/XI8/MM3_g N_BLN<7>_XI0/XI64/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM0 N_XI0/XI64/XI8/NET34_XI0/XI64/XI8/MM0_d
+ N_WL<124>_XI0/XI64/XI8/MM0_g N_BL<7>_XI0/XI64/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM1 N_XI0/XI64/XI8/NET33_XI0/XI64/XI8/MM1_d
+ N_XI0/XI64/XI8/NET34_XI0/XI64/XI8/MM1_g N_VSS_XI0/XI64/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM9 N_XI0/XI64/XI8/NET36_XI0/XI64/XI8/MM9_d
+ N_WL<125>_XI0/XI64/XI8/MM9_g N_BL<7>_XI0/XI64/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM6 N_XI0/XI64/XI8/NET35_XI0/XI64/XI8/MM6_d
+ N_XI0/XI64/XI8/NET36_XI0/XI64/XI8/MM6_g N_VSS_XI0/XI64/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM7 N_XI0/XI64/XI8/NET36_XI0/XI64/XI8/MM7_d
+ N_XI0/XI64/XI8/NET35_XI0/XI64/XI8/MM7_g N_VSS_XI0/XI64/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM8 N_XI0/XI64/XI8/NET35_XI0/XI64/XI8/MM8_d
+ N_WL<125>_XI0/XI64/XI8/MM8_g N_BLN<7>_XI0/XI64/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI8/MM5 N_XI0/XI64/XI8/NET34_XI0/XI64/XI8/MM5_d
+ N_XI0/XI64/XI8/NET33_XI0/XI64/XI8/MM5_g N_VDD_XI0/XI64/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI8/MM4 N_XI0/XI64/XI8/NET33_XI0/XI64/XI8/MM4_d
+ N_XI0/XI64/XI8/NET34_XI0/XI64/XI8/MM4_g N_VDD_XI0/XI64/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI8/MM10 N_XI0/XI64/XI8/NET35_XI0/XI64/XI8/MM10_d
+ N_XI0/XI64/XI8/NET36_XI0/XI64/XI8/MM10_g N_VDD_XI0/XI64/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI8/MM11 N_XI0/XI64/XI8/NET36_XI0/XI64/XI8/MM11_d
+ N_XI0/XI64/XI8/NET35_XI0/XI64/XI8/MM11_g N_VDD_XI0/XI64/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI9/MM2 N_XI0/XI64/XI9/NET34_XI0/XI64/XI9/MM2_d
+ N_XI0/XI64/XI9/NET33_XI0/XI64/XI9/MM2_g N_VSS_XI0/XI64/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM3 N_XI0/XI64/XI9/NET33_XI0/XI64/XI9/MM3_d
+ N_WL<124>_XI0/XI64/XI9/MM3_g N_BLN<6>_XI0/XI64/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM0 N_XI0/XI64/XI9/NET34_XI0/XI64/XI9/MM0_d
+ N_WL<124>_XI0/XI64/XI9/MM0_g N_BL<6>_XI0/XI64/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM1 N_XI0/XI64/XI9/NET33_XI0/XI64/XI9/MM1_d
+ N_XI0/XI64/XI9/NET34_XI0/XI64/XI9/MM1_g N_VSS_XI0/XI64/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM9 N_XI0/XI64/XI9/NET36_XI0/XI64/XI9/MM9_d
+ N_WL<125>_XI0/XI64/XI9/MM9_g N_BL<6>_XI0/XI64/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM6 N_XI0/XI64/XI9/NET35_XI0/XI64/XI9/MM6_d
+ N_XI0/XI64/XI9/NET36_XI0/XI64/XI9/MM6_g N_VSS_XI0/XI64/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM7 N_XI0/XI64/XI9/NET36_XI0/XI64/XI9/MM7_d
+ N_XI0/XI64/XI9/NET35_XI0/XI64/XI9/MM7_g N_VSS_XI0/XI64/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM8 N_XI0/XI64/XI9/NET35_XI0/XI64/XI9/MM8_d
+ N_WL<125>_XI0/XI64/XI9/MM8_g N_BLN<6>_XI0/XI64/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI9/MM5 N_XI0/XI64/XI9/NET34_XI0/XI64/XI9/MM5_d
+ N_XI0/XI64/XI9/NET33_XI0/XI64/XI9/MM5_g N_VDD_XI0/XI64/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI9/MM4 N_XI0/XI64/XI9/NET33_XI0/XI64/XI9/MM4_d
+ N_XI0/XI64/XI9/NET34_XI0/XI64/XI9/MM4_g N_VDD_XI0/XI64/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI9/MM10 N_XI0/XI64/XI9/NET35_XI0/XI64/XI9/MM10_d
+ N_XI0/XI64/XI9/NET36_XI0/XI64/XI9/MM10_g N_VDD_XI0/XI64/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI9/MM11 N_XI0/XI64/XI9/NET36_XI0/XI64/XI9/MM11_d
+ N_XI0/XI64/XI9/NET35_XI0/XI64/XI9/MM11_g N_VDD_XI0/XI64/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI10/MM2 N_XI0/XI64/XI10/NET34_XI0/XI64/XI10/MM2_d
+ N_XI0/XI64/XI10/NET33_XI0/XI64/XI10/MM2_g N_VSS_XI0/XI64/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM3 N_XI0/XI64/XI10/NET33_XI0/XI64/XI10/MM3_d
+ N_WL<124>_XI0/XI64/XI10/MM3_g N_BLN<5>_XI0/XI64/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM0 N_XI0/XI64/XI10/NET34_XI0/XI64/XI10/MM0_d
+ N_WL<124>_XI0/XI64/XI10/MM0_g N_BL<5>_XI0/XI64/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM1 N_XI0/XI64/XI10/NET33_XI0/XI64/XI10/MM1_d
+ N_XI0/XI64/XI10/NET34_XI0/XI64/XI10/MM1_g N_VSS_XI0/XI64/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM9 N_XI0/XI64/XI10/NET36_XI0/XI64/XI10/MM9_d
+ N_WL<125>_XI0/XI64/XI10/MM9_g N_BL<5>_XI0/XI64/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM6 N_XI0/XI64/XI10/NET35_XI0/XI64/XI10/MM6_d
+ N_XI0/XI64/XI10/NET36_XI0/XI64/XI10/MM6_g N_VSS_XI0/XI64/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM7 N_XI0/XI64/XI10/NET36_XI0/XI64/XI10/MM7_d
+ N_XI0/XI64/XI10/NET35_XI0/XI64/XI10/MM7_g N_VSS_XI0/XI64/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM8 N_XI0/XI64/XI10/NET35_XI0/XI64/XI10/MM8_d
+ N_WL<125>_XI0/XI64/XI10/MM8_g N_BLN<5>_XI0/XI64/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI10/MM5 N_XI0/XI64/XI10/NET34_XI0/XI64/XI10/MM5_d
+ N_XI0/XI64/XI10/NET33_XI0/XI64/XI10/MM5_g N_VDD_XI0/XI64/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI10/MM4 N_XI0/XI64/XI10/NET33_XI0/XI64/XI10/MM4_d
+ N_XI0/XI64/XI10/NET34_XI0/XI64/XI10/MM4_g N_VDD_XI0/XI64/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI10/MM10 N_XI0/XI64/XI10/NET35_XI0/XI64/XI10/MM10_d
+ N_XI0/XI64/XI10/NET36_XI0/XI64/XI10/MM10_g N_VDD_XI0/XI64/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI10/MM11 N_XI0/XI64/XI10/NET36_XI0/XI64/XI10/MM11_d
+ N_XI0/XI64/XI10/NET35_XI0/XI64/XI10/MM11_g N_VDD_XI0/XI64/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI11/MM2 N_XI0/XI64/XI11/NET34_XI0/XI64/XI11/MM2_d
+ N_XI0/XI64/XI11/NET33_XI0/XI64/XI11/MM2_g N_VSS_XI0/XI64/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM3 N_XI0/XI64/XI11/NET33_XI0/XI64/XI11/MM3_d
+ N_WL<124>_XI0/XI64/XI11/MM3_g N_BLN<4>_XI0/XI64/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM0 N_XI0/XI64/XI11/NET34_XI0/XI64/XI11/MM0_d
+ N_WL<124>_XI0/XI64/XI11/MM0_g N_BL<4>_XI0/XI64/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM1 N_XI0/XI64/XI11/NET33_XI0/XI64/XI11/MM1_d
+ N_XI0/XI64/XI11/NET34_XI0/XI64/XI11/MM1_g N_VSS_XI0/XI64/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM9 N_XI0/XI64/XI11/NET36_XI0/XI64/XI11/MM9_d
+ N_WL<125>_XI0/XI64/XI11/MM9_g N_BL<4>_XI0/XI64/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM6 N_XI0/XI64/XI11/NET35_XI0/XI64/XI11/MM6_d
+ N_XI0/XI64/XI11/NET36_XI0/XI64/XI11/MM6_g N_VSS_XI0/XI64/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM7 N_XI0/XI64/XI11/NET36_XI0/XI64/XI11/MM7_d
+ N_XI0/XI64/XI11/NET35_XI0/XI64/XI11/MM7_g N_VSS_XI0/XI64/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM8 N_XI0/XI64/XI11/NET35_XI0/XI64/XI11/MM8_d
+ N_WL<125>_XI0/XI64/XI11/MM8_g N_BLN<4>_XI0/XI64/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI11/MM5 N_XI0/XI64/XI11/NET34_XI0/XI64/XI11/MM5_d
+ N_XI0/XI64/XI11/NET33_XI0/XI64/XI11/MM5_g N_VDD_XI0/XI64/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI11/MM4 N_XI0/XI64/XI11/NET33_XI0/XI64/XI11/MM4_d
+ N_XI0/XI64/XI11/NET34_XI0/XI64/XI11/MM4_g N_VDD_XI0/XI64/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI11/MM10 N_XI0/XI64/XI11/NET35_XI0/XI64/XI11/MM10_d
+ N_XI0/XI64/XI11/NET36_XI0/XI64/XI11/MM10_g N_VDD_XI0/XI64/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI11/MM11 N_XI0/XI64/XI11/NET36_XI0/XI64/XI11/MM11_d
+ N_XI0/XI64/XI11/NET35_XI0/XI64/XI11/MM11_g N_VDD_XI0/XI64/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI12/MM2 N_XI0/XI64/XI12/NET34_XI0/XI64/XI12/MM2_d
+ N_XI0/XI64/XI12/NET33_XI0/XI64/XI12/MM2_g N_VSS_XI0/XI64/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM3 N_XI0/XI64/XI12/NET33_XI0/XI64/XI12/MM3_d
+ N_WL<124>_XI0/XI64/XI12/MM3_g N_BLN<3>_XI0/XI64/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM0 N_XI0/XI64/XI12/NET34_XI0/XI64/XI12/MM0_d
+ N_WL<124>_XI0/XI64/XI12/MM0_g N_BL<3>_XI0/XI64/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM1 N_XI0/XI64/XI12/NET33_XI0/XI64/XI12/MM1_d
+ N_XI0/XI64/XI12/NET34_XI0/XI64/XI12/MM1_g N_VSS_XI0/XI64/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM9 N_XI0/XI64/XI12/NET36_XI0/XI64/XI12/MM9_d
+ N_WL<125>_XI0/XI64/XI12/MM9_g N_BL<3>_XI0/XI64/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM6 N_XI0/XI64/XI12/NET35_XI0/XI64/XI12/MM6_d
+ N_XI0/XI64/XI12/NET36_XI0/XI64/XI12/MM6_g N_VSS_XI0/XI64/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM7 N_XI0/XI64/XI12/NET36_XI0/XI64/XI12/MM7_d
+ N_XI0/XI64/XI12/NET35_XI0/XI64/XI12/MM7_g N_VSS_XI0/XI64/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM8 N_XI0/XI64/XI12/NET35_XI0/XI64/XI12/MM8_d
+ N_WL<125>_XI0/XI64/XI12/MM8_g N_BLN<3>_XI0/XI64/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI12/MM5 N_XI0/XI64/XI12/NET34_XI0/XI64/XI12/MM5_d
+ N_XI0/XI64/XI12/NET33_XI0/XI64/XI12/MM5_g N_VDD_XI0/XI64/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI12/MM4 N_XI0/XI64/XI12/NET33_XI0/XI64/XI12/MM4_d
+ N_XI0/XI64/XI12/NET34_XI0/XI64/XI12/MM4_g N_VDD_XI0/XI64/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI12/MM10 N_XI0/XI64/XI12/NET35_XI0/XI64/XI12/MM10_d
+ N_XI0/XI64/XI12/NET36_XI0/XI64/XI12/MM10_g N_VDD_XI0/XI64/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI12/MM11 N_XI0/XI64/XI12/NET36_XI0/XI64/XI12/MM11_d
+ N_XI0/XI64/XI12/NET35_XI0/XI64/XI12/MM11_g N_VDD_XI0/XI64/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI13/MM2 N_XI0/XI64/XI13/NET34_XI0/XI64/XI13/MM2_d
+ N_XI0/XI64/XI13/NET33_XI0/XI64/XI13/MM2_g N_VSS_XI0/XI64/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM3 N_XI0/XI64/XI13/NET33_XI0/XI64/XI13/MM3_d
+ N_WL<124>_XI0/XI64/XI13/MM3_g N_BLN<2>_XI0/XI64/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM0 N_XI0/XI64/XI13/NET34_XI0/XI64/XI13/MM0_d
+ N_WL<124>_XI0/XI64/XI13/MM0_g N_BL<2>_XI0/XI64/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM1 N_XI0/XI64/XI13/NET33_XI0/XI64/XI13/MM1_d
+ N_XI0/XI64/XI13/NET34_XI0/XI64/XI13/MM1_g N_VSS_XI0/XI64/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM9 N_XI0/XI64/XI13/NET36_XI0/XI64/XI13/MM9_d
+ N_WL<125>_XI0/XI64/XI13/MM9_g N_BL<2>_XI0/XI64/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM6 N_XI0/XI64/XI13/NET35_XI0/XI64/XI13/MM6_d
+ N_XI0/XI64/XI13/NET36_XI0/XI64/XI13/MM6_g N_VSS_XI0/XI64/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM7 N_XI0/XI64/XI13/NET36_XI0/XI64/XI13/MM7_d
+ N_XI0/XI64/XI13/NET35_XI0/XI64/XI13/MM7_g N_VSS_XI0/XI64/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM8 N_XI0/XI64/XI13/NET35_XI0/XI64/XI13/MM8_d
+ N_WL<125>_XI0/XI64/XI13/MM8_g N_BLN<2>_XI0/XI64/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI13/MM5 N_XI0/XI64/XI13/NET34_XI0/XI64/XI13/MM5_d
+ N_XI0/XI64/XI13/NET33_XI0/XI64/XI13/MM5_g N_VDD_XI0/XI64/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI13/MM4 N_XI0/XI64/XI13/NET33_XI0/XI64/XI13/MM4_d
+ N_XI0/XI64/XI13/NET34_XI0/XI64/XI13/MM4_g N_VDD_XI0/XI64/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI13/MM10 N_XI0/XI64/XI13/NET35_XI0/XI64/XI13/MM10_d
+ N_XI0/XI64/XI13/NET36_XI0/XI64/XI13/MM10_g N_VDD_XI0/XI64/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI13/MM11 N_XI0/XI64/XI13/NET36_XI0/XI64/XI13/MM11_d
+ N_XI0/XI64/XI13/NET35_XI0/XI64/XI13/MM11_g N_VDD_XI0/XI64/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI14/MM2 N_XI0/XI64/XI14/NET34_XI0/XI64/XI14/MM2_d
+ N_XI0/XI64/XI14/NET33_XI0/XI64/XI14/MM2_g N_VSS_XI0/XI64/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM3 N_XI0/XI64/XI14/NET33_XI0/XI64/XI14/MM3_d
+ N_WL<124>_XI0/XI64/XI14/MM3_g N_BLN<1>_XI0/XI64/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM0 N_XI0/XI64/XI14/NET34_XI0/XI64/XI14/MM0_d
+ N_WL<124>_XI0/XI64/XI14/MM0_g N_BL<1>_XI0/XI64/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM1 N_XI0/XI64/XI14/NET33_XI0/XI64/XI14/MM1_d
+ N_XI0/XI64/XI14/NET34_XI0/XI64/XI14/MM1_g N_VSS_XI0/XI64/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM9 N_XI0/XI64/XI14/NET36_XI0/XI64/XI14/MM9_d
+ N_WL<125>_XI0/XI64/XI14/MM9_g N_BL<1>_XI0/XI64/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM6 N_XI0/XI64/XI14/NET35_XI0/XI64/XI14/MM6_d
+ N_XI0/XI64/XI14/NET36_XI0/XI64/XI14/MM6_g N_VSS_XI0/XI64/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM7 N_XI0/XI64/XI14/NET36_XI0/XI64/XI14/MM7_d
+ N_XI0/XI64/XI14/NET35_XI0/XI64/XI14/MM7_g N_VSS_XI0/XI64/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM8 N_XI0/XI64/XI14/NET35_XI0/XI64/XI14/MM8_d
+ N_WL<125>_XI0/XI64/XI14/MM8_g N_BLN<1>_XI0/XI64/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI14/MM5 N_XI0/XI64/XI14/NET34_XI0/XI64/XI14/MM5_d
+ N_XI0/XI64/XI14/NET33_XI0/XI64/XI14/MM5_g N_VDD_XI0/XI64/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI14/MM4 N_XI0/XI64/XI14/NET33_XI0/XI64/XI14/MM4_d
+ N_XI0/XI64/XI14/NET34_XI0/XI64/XI14/MM4_g N_VDD_XI0/XI64/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI14/MM10 N_XI0/XI64/XI14/NET35_XI0/XI64/XI14/MM10_d
+ N_XI0/XI64/XI14/NET36_XI0/XI64/XI14/MM10_g N_VDD_XI0/XI64/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI14/MM11 N_XI0/XI64/XI14/NET36_XI0/XI64/XI14/MM11_d
+ N_XI0/XI64/XI14/NET35_XI0/XI64/XI14/MM11_g N_VDD_XI0/XI64/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI15/MM2 N_XI0/XI64/XI15/NET34_XI0/XI64/XI15/MM2_d
+ N_XI0/XI64/XI15/NET33_XI0/XI64/XI15/MM2_g N_VSS_XI0/XI64/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM3 N_XI0/XI64/XI15/NET33_XI0/XI64/XI15/MM3_d
+ N_WL<124>_XI0/XI64/XI15/MM3_g N_BLN<0>_XI0/XI64/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM0 N_XI0/XI64/XI15/NET34_XI0/XI64/XI15/MM0_d
+ N_WL<124>_XI0/XI64/XI15/MM0_g N_BL<0>_XI0/XI64/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM1 N_XI0/XI64/XI15/NET33_XI0/XI64/XI15/MM1_d
+ N_XI0/XI64/XI15/NET34_XI0/XI64/XI15/MM1_g N_VSS_XI0/XI64/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM9 N_XI0/XI64/XI15/NET36_XI0/XI64/XI15/MM9_d
+ N_WL<125>_XI0/XI64/XI15/MM9_g N_BL<0>_XI0/XI64/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM6 N_XI0/XI64/XI15/NET35_XI0/XI64/XI15/MM6_d
+ N_XI0/XI64/XI15/NET36_XI0/XI64/XI15/MM6_g N_VSS_XI0/XI64/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM7 N_XI0/XI64/XI15/NET36_XI0/XI64/XI15/MM7_d
+ N_XI0/XI64/XI15/NET35_XI0/XI64/XI15/MM7_g N_VSS_XI0/XI64/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM8 N_XI0/XI64/XI15/NET35_XI0/XI64/XI15/MM8_d
+ N_WL<125>_XI0/XI64/XI15/MM8_g N_BLN<0>_XI0/XI64/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI64/XI15/MM5 N_XI0/XI64/XI15/NET34_XI0/XI64/XI15/MM5_d
+ N_XI0/XI64/XI15/NET33_XI0/XI64/XI15/MM5_g N_VDD_XI0/XI64/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI15/MM4 N_XI0/XI64/XI15/NET33_XI0/XI64/XI15/MM4_d
+ N_XI0/XI64/XI15/NET34_XI0/XI64/XI15/MM4_g N_VDD_XI0/XI64/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI15/MM10 N_XI0/XI64/XI15/NET35_XI0/XI64/XI15/MM10_d
+ N_XI0/XI64/XI15/NET36_XI0/XI64/XI15/MM10_g N_VDD_XI0/XI64/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI64/XI15/MM11 N_XI0/XI64/XI15/NET36_XI0/XI64/XI15/MM11_d
+ N_XI0/XI64/XI15/NET35_XI0/XI64/XI15/MM11_g N_VDD_XI0/XI64/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI0/MM2 N_XI0/XI65/XI0/NET34_XI0/XI65/XI0/MM2_d
+ N_XI0/XI65/XI0/NET33_XI0/XI65/XI0/MM2_g N_VSS_XI0/XI65/XI0/MM2_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM3 N_XI0/XI65/XI0/NET33_XI0/XI65/XI0/MM3_d
+ N_WL<126>_XI0/XI65/XI0/MM3_g N_BLN<15>_XI0/XI65/XI0/MM3_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM0 N_XI0/XI65/XI0/NET34_XI0/XI65/XI0/MM0_d
+ N_WL<126>_XI0/XI65/XI0/MM0_g N_BL<15>_XI0/XI65/XI0/MM0_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM1 N_XI0/XI65/XI0/NET33_XI0/XI65/XI0/MM1_d
+ N_XI0/XI65/XI0/NET34_XI0/XI65/XI0/MM1_g N_VSS_XI0/XI65/XI0/MM1_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM9 N_XI0/XI65/XI0/NET36_XI0/XI65/XI0/MM9_d
+ N_WL<127>_XI0/XI65/XI0/MM9_g N_BL<15>_XI0/XI65/XI0/MM9_s N_VSS_XI1/XI0/MM0_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM6 N_XI0/XI65/XI0/NET35_XI0/XI65/XI0/MM6_d
+ N_XI0/XI65/XI0/NET36_XI0/XI65/XI0/MM6_g N_VSS_XI0/XI65/XI0/MM6_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM7 N_XI0/XI65/XI0/NET36_XI0/XI65/XI0/MM7_d
+ N_XI0/XI65/XI0/NET35_XI0/XI65/XI0/MM7_g N_VSS_XI0/XI65/XI0/MM7_s
+ N_VSS_XI1/XI0/MM0_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM8 N_XI0/XI65/XI0/NET35_XI0/XI65/XI0/MM8_d
+ N_WL<127>_XI0/XI65/XI0/MM8_g N_BLN<15>_XI0/XI65/XI0/MM8_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI0/MM5 N_XI0/XI65/XI0/NET34_XI0/XI65/XI0/MM5_d
+ N_XI0/XI65/XI0/NET33_XI0/XI65/XI0/MM5_g N_VDD_XI0/XI65/XI0/MM5_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI0/MM4 N_XI0/XI65/XI0/NET33_XI0/XI65/XI0/MM4_d
+ N_XI0/XI65/XI0/NET34_XI0/XI65/XI0/MM4_g N_VDD_XI0/XI65/XI0/MM4_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI0/MM10 N_XI0/XI65/XI0/NET35_XI0/XI65/XI0/MM10_d
+ N_XI0/XI65/XI0/NET36_XI0/XI65/XI0/MM10_g N_VDD_XI0/XI65/XI0/MM10_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI0/MM11 N_XI0/XI65/XI0/NET36_XI0/XI65/XI0/MM11_d
+ N_XI0/XI65/XI0/NET35_XI0/XI65/XI0/MM11_g N_VDD_XI0/XI65/XI0/MM11_s
+ N_VDD_XI1/XI0/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI1/MM2 N_XI0/XI65/XI1/NET34_XI0/XI65/XI1/MM2_d
+ N_XI0/XI65/XI1/NET33_XI0/XI65/XI1/MM2_g N_VSS_XI0/XI65/XI1/MM2_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM3 N_XI0/XI65/XI1/NET33_XI0/XI65/XI1/MM3_d
+ N_WL<126>_XI0/XI65/XI1/MM3_g N_BLN<14>_XI0/XI65/XI1/MM3_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM0 N_XI0/XI65/XI1/NET34_XI0/XI65/XI1/MM0_d
+ N_WL<126>_XI0/XI65/XI1/MM0_g N_BL<14>_XI0/XI65/XI1/MM0_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM1 N_XI0/XI65/XI1/NET33_XI0/XI65/XI1/MM1_d
+ N_XI0/XI65/XI1/NET34_XI0/XI65/XI1/MM1_g N_VSS_XI0/XI65/XI1/MM1_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM9 N_XI0/XI65/XI1/NET36_XI0/XI65/XI1/MM9_d
+ N_WL<127>_XI0/XI65/XI1/MM9_g N_BL<14>_XI0/XI65/XI1/MM9_s N_VSS_XI1/XI0/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM6 N_XI0/XI65/XI1/NET35_XI0/XI65/XI1/MM6_d
+ N_XI0/XI65/XI1/NET36_XI0/XI65/XI1/MM6_g N_VSS_XI0/XI65/XI1/MM6_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM7 N_XI0/XI65/XI1/NET36_XI0/XI65/XI1/MM7_d
+ N_XI0/XI65/XI1/NET35_XI0/XI65/XI1/MM7_g N_VSS_XI0/XI65/XI1/MM7_s
+ N_VSS_XI1/XI0/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM8 N_XI0/XI65/XI1/NET35_XI0/XI65/XI1/MM8_d
+ N_WL<127>_XI0/XI65/XI1/MM8_g N_BLN<14>_XI0/XI65/XI1/MM8_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI1/MM5 N_XI0/XI65/XI1/NET34_XI0/XI65/XI1/MM5_d
+ N_XI0/XI65/XI1/NET33_XI0/XI65/XI1/MM5_g N_VDD_XI0/XI65/XI1/MM5_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI1/MM4 N_XI0/XI65/XI1/NET33_XI0/XI65/XI1/MM4_d
+ N_XI0/XI65/XI1/NET34_XI0/XI65/XI1/MM4_g N_VDD_XI0/XI65/XI1/MM4_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI1/MM10 N_XI0/XI65/XI1/NET35_XI0/XI65/XI1/MM10_d
+ N_XI0/XI65/XI1/NET36_XI0/XI65/XI1/MM10_g N_VDD_XI0/XI65/XI1/MM10_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI1/MM11 N_XI0/XI65/XI1/NET36_XI0/XI65/XI1/MM11_d
+ N_XI0/XI65/XI1/NET35_XI0/XI65/XI1/MM11_g N_VDD_XI0/XI65/XI1/MM11_s
+ N_VDD_XI1/XI4/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI2/MM2 N_XI0/XI65/XI2/NET34_XI0/XI65/XI2/MM2_d
+ N_XI0/XI65/XI2/NET33_XI0/XI65/XI2/MM2_g N_VSS_XI0/XI65/XI2/MM2_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM3 N_XI0/XI65/XI2/NET33_XI0/XI65/XI2/MM3_d
+ N_WL<126>_XI0/XI65/XI2/MM3_g N_BLN<13>_XI0/XI65/XI2/MM3_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM0 N_XI0/XI65/XI2/NET34_XI0/XI65/XI2/MM0_d
+ N_WL<126>_XI0/XI65/XI2/MM0_g N_BL<13>_XI0/XI65/XI2/MM0_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM1 N_XI0/XI65/XI2/NET33_XI0/XI65/XI2/MM1_d
+ N_XI0/XI65/XI2/NET34_XI0/XI65/XI2/MM1_g N_VSS_XI0/XI65/XI2/MM1_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM9 N_XI0/XI65/XI2/NET36_XI0/XI65/XI2/MM9_d
+ N_WL<127>_XI0/XI65/XI2/MM9_g N_BL<13>_XI0/XI65/XI2/MM9_s N_VSS_XI1/XI4/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM6 N_XI0/XI65/XI2/NET35_XI0/XI65/XI2/MM6_d
+ N_XI0/XI65/XI2/NET36_XI0/XI65/XI2/MM6_g N_VSS_XI0/XI65/XI2/MM6_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM7 N_XI0/XI65/XI2/NET36_XI0/XI65/XI2/MM7_d
+ N_XI0/XI65/XI2/NET35_XI0/XI65/XI2/MM7_g N_VSS_XI0/XI65/XI2/MM7_s
+ N_VSS_XI1/XI4/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM8 N_XI0/XI65/XI2/NET35_XI0/XI65/XI2/MM8_d
+ N_WL<127>_XI0/XI65/XI2/MM8_g N_BLN<13>_XI0/XI65/XI2/MM8_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI2/MM5 N_XI0/XI65/XI2/NET34_XI0/XI65/XI2/MM5_d
+ N_XI0/XI65/XI2/NET33_XI0/XI65/XI2/MM5_g N_VDD_XI0/XI65/XI2/MM5_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI2/MM4 N_XI0/XI65/XI2/NET33_XI0/XI65/XI2/MM4_d
+ N_XI0/XI65/XI2/NET34_XI0/XI65/XI2/MM4_g N_VDD_XI0/XI65/XI2/MM4_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI2/MM10 N_XI0/XI65/XI2/NET35_XI0/XI65/XI2/MM10_d
+ N_XI0/XI65/XI2/NET36_XI0/XI65/XI2/MM10_g N_VDD_XI0/XI65/XI2/MM10_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI2/MM11 N_XI0/XI65/XI2/NET36_XI0/XI65/XI2/MM11_d
+ N_XI0/XI65/XI2/NET35_XI0/XI65/XI2/MM11_g N_VDD_XI0/XI65/XI2/MM11_s
+ N_VDD_XI1/XI8/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI3/MM2 N_XI0/XI65/XI3/NET34_XI0/XI65/XI3/MM2_d
+ N_XI0/XI65/XI3/NET33_XI0/XI65/XI3/MM2_g N_VSS_XI0/XI65/XI3/MM2_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM3 N_XI0/XI65/XI3/NET33_XI0/XI65/XI3/MM3_d
+ N_WL<126>_XI0/XI65/XI3/MM3_g N_BLN<12>_XI0/XI65/XI3/MM3_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM0 N_XI0/XI65/XI3/NET34_XI0/XI65/XI3/MM0_d
+ N_WL<126>_XI0/XI65/XI3/MM0_g N_BL<12>_XI0/XI65/XI3/MM0_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM1 N_XI0/XI65/XI3/NET33_XI0/XI65/XI3/MM1_d
+ N_XI0/XI65/XI3/NET34_XI0/XI65/XI3/MM1_g N_VSS_XI0/XI65/XI3/MM1_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM9 N_XI0/XI65/XI3/NET36_XI0/XI65/XI3/MM9_d
+ N_WL<127>_XI0/XI65/XI3/MM9_g N_BL<12>_XI0/XI65/XI3/MM9_s N_VSS_XI1/XI8/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM6 N_XI0/XI65/XI3/NET35_XI0/XI65/XI3/MM6_d
+ N_XI0/XI65/XI3/NET36_XI0/XI65/XI3/MM6_g N_VSS_XI0/XI65/XI3/MM6_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM7 N_XI0/XI65/XI3/NET36_XI0/XI65/XI3/MM7_d
+ N_XI0/XI65/XI3/NET35_XI0/XI65/XI3/MM7_g N_VSS_XI0/XI65/XI3/MM7_s
+ N_VSS_XI1/XI8/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM8 N_XI0/XI65/XI3/NET35_XI0/XI65/XI3/MM8_d
+ N_WL<127>_XI0/XI65/XI3/MM8_g N_BLN<12>_XI0/XI65/XI3/MM8_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI3/MM5 N_XI0/XI65/XI3/NET34_XI0/XI65/XI3/MM5_d
+ N_XI0/XI65/XI3/NET33_XI0/XI65/XI3/MM5_g N_VDD_XI0/XI65/XI3/MM5_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI3/MM4 N_XI0/XI65/XI3/NET33_XI0/XI65/XI3/MM4_d
+ N_XI0/XI65/XI3/NET34_XI0/XI65/XI3/MM4_g N_VDD_XI0/XI65/XI3/MM4_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI3/MM10 N_XI0/XI65/XI3/NET35_XI0/XI65/XI3/MM10_d
+ N_XI0/XI65/XI3/NET36_XI0/XI65/XI3/MM10_g N_VDD_XI0/XI65/XI3/MM10_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI3/MM11 N_XI0/XI65/XI3/NET36_XI0/XI65/XI3/MM11_d
+ N_XI0/XI65/XI3/NET35_XI0/XI65/XI3/MM11_g N_VDD_XI0/XI65/XI3/MM11_s
+ N_VDD_XI1/XI12/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI4/MM2 N_XI0/XI65/XI4/NET34_XI0/XI65/XI4/MM2_d
+ N_XI0/XI65/XI4/NET33_XI0/XI65/XI4/MM2_g N_VSS_XI0/XI65/XI4/MM2_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM3 N_XI0/XI65/XI4/NET33_XI0/XI65/XI4/MM3_d
+ N_WL<126>_XI0/XI65/XI4/MM3_g N_BLN<11>_XI0/XI65/XI4/MM3_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM0 N_XI0/XI65/XI4/NET34_XI0/XI65/XI4/MM0_d
+ N_WL<126>_XI0/XI65/XI4/MM0_g N_BL<11>_XI0/XI65/XI4/MM0_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM1 N_XI0/XI65/XI4/NET33_XI0/XI65/XI4/MM1_d
+ N_XI0/XI65/XI4/NET34_XI0/XI65/XI4/MM1_g N_VSS_XI0/XI65/XI4/MM1_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM9 N_XI0/XI65/XI4/NET36_XI0/XI65/XI4/MM9_d
+ N_WL<127>_XI0/XI65/XI4/MM9_g N_BL<11>_XI0/XI65/XI4/MM9_s N_VSS_XI1/XI12/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM6 N_XI0/XI65/XI4/NET35_XI0/XI65/XI4/MM6_d
+ N_XI0/XI65/XI4/NET36_XI0/XI65/XI4/MM6_g N_VSS_XI0/XI65/XI4/MM6_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM7 N_XI0/XI65/XI4/NET36_XI0/XI65/XI4/MM7_d
+ N_XI0/XI65/XI4/NET35_XI0/XI65/XI4/MM7_g N_VSS_XI0/XI65/XI4/MM7_s
+ N_VSS_XI1/XI12/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM8 N_XI0/XI65/XI4/NET35_XI0/XI65/XI4/MM8_d
+ N_WL<127>_XI0/XI65/XI4/MM8_g N_BLN<11>_XI0/XI65/XI4/MM8_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI4/MM5 N_XI0/XI65/XI4/NET34_XI0/XI65/XI4/MM5_d
+ N_XI0/XI65/XI4/NET33_XI0/XI65/XI4/MM5_g N_VDD_XI0/XI65/XI4/MM5_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI4/MM4 N_XI0/XI65/XI4/NET33_XI0/XI65/XI4/MM4_d
+ N_XI0/XI65/XI4/NET34_XI0/XI65/XI4/MM4_g N_VDD_XI0/XI65/XI4/MM4_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI4/MM10 N_XI0/XI65/XI4/NET35_XI0/XI65/XI4/MM10_d
+ N_XI0/XI65/XI4/NET36_XI0/XI65/XI4/MM10_g N_VDD_XI0/XI65/XI4/MM10_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI4/MM11 N_XI0/XI65/XI4/NET36_XI0/XI65/XI4/MM11_d
+ N_XI0/XI65/XI4/NET35_XI0/XI65/XI4/MM11_g N_VDD_XI0/XI65/XI4/MM11_s
+ N_VDD_XI1/XI1/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI5/MM2 N_XI0/XI65/XI5/NET34_XI0/XI65/XI5/MM2_d
+ N_XI0/XI65/XI5/NET33_XI0/XI65/XI5/MM2_g N_VSS_XI0/XI65/XI5/MM2_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM3 N_XI0/XI65/XI5/NET33_XI0/XI65/XI5/MM3_d
+ N_WL<126>_XI0/XI65/XI5/MM3_g N_BLN<10>_XI0/XI65/XI5/MM3_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM0 N_XI0/XI65/XI5/NET34_XI0/XI65/XI5/MM0_d
+ N_WL<126>_XI0/XI65/XI5/MM0_g N_BL<10>_XI0/XI65/XI5/MM0_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM1 N_XI0/XI65/XI5/NET33_XI0/XI65/XI5/MM1_d
+ N_XI0/XI65/XI5/NET34_XI0/XI65/XI5/MM1_g N_VSS_XI0/XI65/XI5/MM1_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM9 N_XI0/XI65/XI5/NET36_XI0/XI65/XI5/MM9_d
+ N_WL<127>_XI0/XI65/XI5/MM9_g N_BL<10>_XI0/XI65/XI5/MM9_s N_VSS_XI1/XI1/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM6 N_XI0/XI65/XI5/NET35_XI0/XI65/XI5/MM6_d
+ N_XI0/XI65/XI5/NET36_XI0/XI65/XI5/MM6_g N_VSS_XI0/XI65/XI5/MM6_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM7 N_XI0/XI65/XI5/NET36_XI0/XI65/XI5/MM7_d
+ N_XI0/XI65/XI5/NET35_XI0/XI65/XI5/MM7_g N_VSS_XI0/XI65/XI5/MM7_s
+ N_VSS_XI1/XI1/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM8 N_XI0/XI65/XI5/NET35_XI0/XI65/XI5/MM8_d
+ N_WL<127>_XI0/XI65/XI5/MM8_g N_BLN<10>_XI0/XI65/XI5/MM8_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI5/MM5 N_XI0/XI65/XI5/NET34_XI0/XI65/XI5/MM5_d
+ N_XI0/XI65/XI5/NET33_XI0/XI65/XI5/MM5_g N_VDD_XI0/XI65/XI5/MM5_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI5/MM4 N_XI0/XI65/XI5/NET33_XI0/XI65/XI5/MM4_d
+ N_XI0/XI65/XI5/NET34_XI0/XI65/XI5/MM4_g N_VDD_XI0/XI65/XI5/MM4_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI5/MM10 N_XI0/XI65/XI5/NET35_XI0/XI65/XI5/MM10_d
+ N_XI0/XI65/XI5/NET36_XI0/XI65/XI5/MM10_g N_VDD_XI0/XI65/XI5/MM10_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI5/MM11 N_XI0/XI65/XI5/NET36_XI0/XI65/XI5/MM11_d
+ N_XI0/XI65/XI5/NET35_XI0/XI65/XI5/MM11_g N_VDD_XI0/XI65/XI5/MM11_s
+ N_VDD_XI1/XI5/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI6/MM2 N_XI0/XI65/XI6/NET34_XI0/XI65/XI6/MM2_d
+ N_XI0/XI65/XI6/NET33_XI0/XI65/XI6/MM2_g N_VSS_XI0/XI65/XI6/MM2_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM3 N_XI0/XI65/XI6/NET33_XI0/XI65/XI6/MM3_d
+ N_WL<126>_XI0/XI65/XI6/MM3_g N_BLN<9>_XI0/XI65/XI6/MM3_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM0 N_XI0/XI65/XI6/NET34_XI0/XI65/XI6/MM0_d
+ N_WL<126>_XI0/XI65/XI6/MM0_g N_BL<9>_XI0/XI65/XI6/MM0_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM1 N_XI0/XI65/XI6/NET33_XI0/XI65/XI6/MM1_d
+ N_XI0/XI65/XI6/NET34_XI0/XI65/XI6/MM1_g N_VSS_XI0/XI65/XI6/MM1_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM9 N_XI0/XI65/XI6/NET36_XI0/XI65/XI6/MM9_d
+ N_WL<127>_XI0/XI65/XI6/MM9_g N_BL<9>_XI0/XI65/XI6/MM9_s N_VSS_XI1/XI5/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM6 N_XI0/XI65/XI6/NET35_XI0/XI65/XI6/MM6_d
+ N_XI0/XI65/XI6/NET36_XI0/XI65/XI6/MM6_g N_VSS_XI0/XI65/XI6/MM6_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM7 N_XI0/XI65/XI6/NET36_XI0/XI65/XI6/MM7_d
+ N_XI0/XI65/XI6/NET35_XI0/XI65/XI6/MM7_g N_VSS_XI0/XI65/XI6/MM7_s
+ N_VSS_XI1/XI5/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM8 N_XI0/XI65/XI6/NET35_XI0/XI65/XI6/MM8_d
+ N_WL<127>_XI0/XI65/XI6/MM8_g N_BLN<9>_XI0/XI65/XI6/MM8_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI6/MM5 N_XI0/XI65/XI6/NET34_XI0/XI65/XI6/MM5_d
+ N_XI0/XI65/XI6/NET33_XI0/XI65/XI6/MM5_g N_VDD_XI0/XI65/XI6/MM5_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI6/MM4 N_XI0/XI65/XI6/NET33_XI0/XI65/XI6/MM4_d
+ N_XI0/XI65/XI6/NET34_XI0/XI65/XI6/MM4_g N_VDD_XI0/XI65/XI6/MM4_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI6/MM10 N_XI0/XI65/XI6/NET35_XI0/XI65/XI6/MM10_d
+ N_XI0/XI65/XI6/NET36_XI0/XI65/XI6/MM10_g N_VDD_XI0/XI65/XI6/MM10_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI6/MM11 N_XI0/XI65/XI6/NET36_XI0/XI65/XI6/MM11_d
+ N_XI0/XI65/XI6/NET35_XI0/XI65/XI6/MM11_g N_VDD_XI0/XI65/XI6/MM11_s
+ N_VDD_XI1/XI9/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI7/MM2 N_XI0/XI65/XI7/NET34_XI0/XI65/XI7/MM2_d
+ N_XI0/XI65/XI7/NET33_XI0/XI65/XI7/MM2_g N_VSS_XI0/XI65/XI7/MM2_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM3 N_XI0/XI65/XI7/NET33_XI0/XI65/XI7/MM3_d
+ N_WL<126>_XI0/XI65/XI7/MM3_g N_BLN<8>_XI0/XI65/XI7/MM3_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM0 N_XI0/XI65/XI7/NET34_XI0/XI65/XI7/MM0_d
+ N_WL<126>_XI0/XI65/XI7/MM0_g N_BL<8>_XI0/XI65/XI7/MM0_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM1 N_XI0/XI65/XI7/NET33_XI0/XI65/XI7/MM1_d
+ N_XI0/XI65/XI7/NET34_XI0/XI65/XI7/MM1_g N_VSS_XI0/XI65/XI7/MM1_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM9 N_XI0/XI65/XI7/NET36_XI0/XI65/XI7/MM9_d
+ N_WL<127>_XI0/XI65/XI7/MM9_g N_BL<8>_XI0/XI65/XI7/MM9_s N_VSS_XI1/XI9/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM6 N_XI0/XI65/XI7/NET35_XI0/XI65/XI7/MM6_d
+ N_XI0/XI65/XI7/NET36_XI0/XI65/XI7/MM6_g N_VSS_XI0/XI65/XI7/MM6_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM7 N_XI0/XI65/XI7/NET36_XI0/XI65/XI7/MM7_d
+ N_XI0/XI65/XI7/NET35_XI0/XI65/XI7/MM7_g N_VSS_XI0/XI65/XI7/MM7_s
+ N_VSS_XI1/XI9/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM8 N_XI0/XI65/XI7/NET35_XI0/XI65/XI7/MM8_d
+ N_WL<127>_XI0/XI65/XI7/MM8_g N_BLN<8>_XI0/XI65/XI7/MM8_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI7/MM5 N_XI0/XI65/XI7/NET34_XI0/XI65/XI7/MM5_d
+ N_XI0/XI65/XI7/NET33_XI0/XI65/XI7/MM5_g N_VDD_XI0/XI65/XI7/MM5_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI7/MM4 N_XI0/XI65/XI7/NET33_XI0/XI65/XI7/MM4_d
+ N_XI0/XI65/XI7/NET34_XI0/XI65/XI7/MM4_g N_VDD_XI0/XI65/XI7/MM4_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI7/MM10 N_XI0/XI65/XI7/NET35_XI0/XI65/XI7/MM10_d
+ N_XI0/XI65/XI7/NET36_XI0/XI65/XI7/MM10_g N_VDD_XI0/XI65/XI7/MM10_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI7/MM11 N_XI0/XI65/XI7/NET36_XI0/XI65/XI7/MM11_d
+ N_XI0/XI65/XI7/NET35_XI0/XI65/XI7/MM11_g N_VDD_XI0/XI65/XI7/MM11_s
+ N_VDD_XI1/XI13/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI8/MM2 N_XI0/XI65/XI8/NET34_XI0/XI65/XI8/MM2_d
+ N_XI0/XI65/XI8/NET33_XI0/XI65/XI8/MM2_g N_VSS_XI0/XI65/XI8/MM2_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM3 N_XI0/XI65/XI8/NET33_XI0/XI65/XI8/MM3_d
+ N_WL<126>_XI0/XI65/XI8/MM3_g N_BLN<7>_XI0/XI65/XI8/MM3_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM0 N_XI0/XI65/XI8/NET34_XI0/XI65/XI8/MM0_d
+ N_WL<126>_XI0/XI65/XI8/MM0_g N_BL<7>_XI0/XI65/XI8/MM0_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM1 N_XI0/XI65/XI8/NET33_XI0/XI65/XI8/MM1_d
+ N_XI0/XI65/XI8/NET34_XI0/XI65/XI8/MM1_g N_VSS_XI0/XI65/XI8/MM1_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM9 N_XI0/XI65/XI8/NET36_XI0/XI65/XI8/MM9_d
+ N_WL<127>_XI0/XI65/XI8/MM9_g N_BL<7>_XI0/XI65/XI8/MM9_s N_VSS_XI1/XI13/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM6 N_XI0/XI65/XI8/NET35_XI0/XI65/XI8/MM6_d
+ N_XI0/XI65/XI8/NET36_XI0/XI65/XI8/MM6_g N_VSS_XI0/XI65/XI8/MM6_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM7 N_XI0/XI65/XI8/NET36_XI0/XI65/XI8/MM7_d
+ N_XI0/XI65/XI8/NET35_XI0/XI65/XI8/MM7_g N_VSS_XI0/XI65/XI8/MM7_s
+ N_VSS_XI1/XI13/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM8 N_XI0/XI65/XI8/NET35_XI0/XI65/XI8/MM8_d
+ N_WL<127>_XI0/XI65/XI8/MM8_g N_BLN<7>_XI0/XI65/XI8/MM8_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI8/MM5 N_XI0/XI65/XI8/NET34_XI0/XI65/XI8/MM5_d
+ N_XI0/XI65/XI8/NET33_XI0/XI65/XI8/MM5_g N_VDD_XI0/XI65/XI8/MM5_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI8/MM4 N_XI0/XI65/XI8/NET33_XI0/XI65/XI8/MM4_d
+ N_XI0/XI65/XI8/NET34_XI0/XI65/XI8/MM4_g N_VDD_XI0/XI65/XI8/MM4_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI8/MM10 N_XI0/XI65/XI8/NET35_XI0/XI65/XI8/MM10_d
+ N_XI0/XI65/XI8/NET36_XI0/XI65/XI8/MM10_g N_VDD_XI0/XI65/XI8/MM10_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI8/MM11 N_XI0/XI65/XI8/NET36_XI0/XI65/XI8/MM11_d
+ N_XI0/XI65/XI8/NET35_XI0/XI65/XI8/MM11_g N_VDD_XI0/XI65/XI8/MM11_s
+ N_VDD_XI1/XI2/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI9/MM2 N_XI0/XI65/XI9/NET34_XI0/XI65/XI9/MM2_d
+ N_XI0/XI65/XI9/NET33_XI0/XI65/XI9/MM2_g N_VSS_XI0/XI65/XI9/MM2_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM3 N_XI0/XI65/XI9/NET33_XI0/XI65/XI9/MM3_d
+ N_WL<126>_XI0/XI65/XI9/MM3_g N_BLN<6>_XI0/XI65/XI9/MM3_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM0 N_XI0/XI65/XI9/NET34_XI0/XI65/XI9/MM0_d
+ N_WL<126>_XI0/XI65/XI9/MM0_g N_BL<6>_XI0/XI65/XI9/MM0_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM1 N_XI0/XI65/XI9/NET33_XI0/XI65/XI9/MM1_d
+ N_XI0/XI65/XI9/NET34_XI0/XI65/XI9/MM1_g N_VSS_XI0/XI65/XI9/MM1_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM9 N_XI0/XI65/XI9/NET36_XI0/XI65/XI9/MM9_d
+ N_WL<127>_XI0/XI65/XI9/MM9_g N_BL<6>_XI0/XI65/XI9/MM9_s N_VSS_XI1/XI2/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM6 N_XI0/XI65/XI9/NET35_XI0/XI65/XI9/MM6_d
+ N_XI0/XI65/XI9/NET36_XI0/XI65/XI9/MM6_g N_VSS_XI0/XI65/XI9/MM6_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM7 N_XI0/XI65/XI9/NET36_XI0/XI65/XI9/MM7_d
+ N_XI0/XI65/XI9/NET35_XI0/XI65/XI9/MM7_g N_VSS_XI0/XI65/XI9/MM7_s
+ N_VSS_XI1/XI2/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM8 N_XI0/XI65/XI9/NET35_XI0/XI65/XI9/MM8_d
+ N_WL<127>_XI0/XI65/XI9/MM8_g N_BLN<6>_XI0/XI65/XI9/MM8_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI9/MM5 N_XI0/XI65/XI9/NET34_XI0/XI65/XI9/MM5_d
+ N_XI0/XI65/XI9/NET33_XI0/XI65/XI9/MM5_g N_VDD_XI0/XI65/XI9/MM5_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI9/MM4 N_XI0/XI65/XI9/NET33_XI0/XI65/XI9/MM4_d
+ N_XI0/XI65/XI9/NET34_XI0/XI65/XI9/MM4_g N_VDD_XI0/XI65/XI9/MM4_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI9/MM10 N_XI0/XI65/XI9/NET35_XI0/XI65/XI9/MM10_d
+ N_XI0/XI65/XI9/NET36_XI0/XI65/XI9/MM10_g N_VDD_XI0/XI65/XI9/MM10_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI9/MM11 N_XI0/XI65/XI9/NET36_XI0/XI65/XI9/MM11_d
+ N_XI0/XI65/XI9/NET35_XI0/XI65/XI9/MM11_g N_VDD_XI0/XI65/XI9/MM11_s
+ N_VDD_XI1/XI6/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI10/MM2 N_XI0/XI65/XI10/NET34_XI0/XI65/XI10/MM2_d
+ N_XI0/XI65/XI10/NET33_XI0/XI65/XI10/MM2_g N_VSS_XI0/XI65/XI10/MM2_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM3 N_XI0/XI65/XI10/NET33_XI0/XI65/XI10/MM3_d
+ N_WL<126>_XI0/XI65/XI10/MM3_g N_BLN<5>_XI0/XI65/XI10/MM3_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM0 N_XI0/XI65/XI10/NET34_XI0/XI65/XI10/MM0_d
+ N_WL<126>_XI0/XI65/XI10/MM0_g N_BL<5>_XI0/XI65/XI10/MM0_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM1 N_XI0/XI65/XI10/NET33_XI0/XI65/XI10/MM1_d
+ N_XI0/XI65/XI10/NET34_XI0/XI65/XI10/MM1_g N_VSS_XI0/XI65/XI10/MM1_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM9 N_XI0/XI65/XI10/NET36_XI0/XI65/XI10/MM9_d
+ N_WL<127>_XI0/XI65/XI10/MM9_g N_BL<5>_XI0/XI65/XI10/MM9_s N_VSS_XI1/XI6/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM6 N_XI0/XI65/XI10/NET35_XI0/XI65/XI10/MM6_d
+ N_XI0/XI65/XI10/NET36_XI0/XI65/XI10/MM6_g N_VSS_XI0/XI65/XI10/MM6_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM7 N_XI0/XI65/XI10/NET36_XI0/XI65/XI10/MM7_d
+ N_XI0/XI65/XI10/NET35_XI0/XI65/XI10/MM7_g N_VSS_XI0/XI65/XI10/MM7_s
+ N_VSS_XI1/XI6/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM8 N_XI0/XI65/XI10/NET35_XI0/XI65/XI10/MM8_d
+ N_WL<127>_XI0/XI65/XI10/MM8_g N_BLN<5>_XI0/XI65/XI10/MM8_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI10/MM5 N_XI0/XI65/XI10/NET34_XI0/XI65/XI10/MM5_d
+ N_XI0/XI65/XI10/NET33_XI0/XI65/XI10/MM5_g N_VDD_XI0/XI65/XI10/MM5_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI10/MM4 N_XI0/XI65/XI10/NET33_XI0/XI65/XI10/MM4_d
+ N_XI0/XI65/XI10/NET34_XI0/XI65/XI10/MM4_g N_VDD_XI0/XI65/XI10/MM4_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI10/MM10 N_XI0/XI65/XI10/NET35_XI0/XI65/XI10/MM10_d
+ N_XI0/XI65/XI10/NET36_XI0/XI65/XI10/MM10_g N_VDD_XI0/XI65/XI10/MM10_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI10/MM11 N_XI0/XI65/XI10/NET36_XI0/XI65/XI10/MM11_d
+ N_XI0/XI65/XI10/NET35_XI0/XI65/XI10/MM11_g N_VDD_XI0/XI65/XI10/MM11_s
+ N_VDD_XI1/XI10/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI11/MM2 N_XI0/XI65/XI11/NET34_XI0/XI65/XI11/MM2_d
+ N_XI0/XI65/XI11/NET33_XI0/XI65/XI11/MM2_g N_VSS_XI0/XI65/XI11/MM2_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM3 N_XI0/XI65/XI11/NET33_XI0/XI65/XI11/MM3_d
+ N_WL<126>_XI0/XI65/XI11/MM3_g N_BLN<4>_XI0/XI65/XI11/MM3_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM0 N_XI0/XI65/XI11/NET34_XI0/XI65/XI11/MM0_d
+ N_WL<126>_XI0/XI65/XI11/MM0_g N_BL<4>_XI0/XI65/XI11/MM0_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM1 N_XI0/XI65/XI11/NET33_XI0/XI65/XI11/MM1_d
+ N_XI0/XI65/XI11/NET34_XI0/XI65/XI11/MM1_g N_VSS_XI0/XI65/XI11/MM1_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM9 N_XI0/XI65/XI11/NET36_XI0/XI65/XI11/MM9_d
+ N_WL<127>_XI0/XI65/XI11/MM9_g N_BL<4>_XI0/XI65/XI11/MM9_s N_VSS_XI1/XI10/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM6 N_XI0/XI65/XI11/NET35_XI0/XI65/XI11/MM6_d
+ N_XI0/XI65/XI11/NET36_XI0/XI65/XI11/MM6_g N_VSS_XI0/XI65/XI11/MM6_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM7 N_XI0/XI65/XI11/NET36_XI0/XI65/XI11/MM7_d
+ N_XI0/XI65/XI11/NET35_XI0/XI65/XI11/MM7_g N_VSS_XI0/XI65/XI11/MM7_s
+ N_VSS_XI1/XI10/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM8 N_XI0/XI65/XI11/NET35_XI0/XI65/XI11/MM8_d
+ N_WL<127>_XI0/XI65/XI11/MM8_g N_BLN<4>_XI0/XI65/XI11/MM8_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI11/MM5 N_XI0/XI65/XI11/NET34_XI0/XI65/XI11/MM5_d
+ N_XI0/XI65/XI11/NET33_XI0/XI65/XI11/MM5_g N_VDD_XI0/XI65/XI11/MM5_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI11/MM4 N_XI0/XI65/XI11/NET33_XI0/XI65/XI11/MM4_d
+ N_XI0/XI65/XI11/NET34_XI0/XI65/XI11/MM4_g N_VDD_XI0/XI65/XI11/MM4_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI11/MM10 N_XI0/XI65/XI11/NET35_XI0/XI65/XI11/MM10_d
+ N_XI0/XI65/XI11/NET36_XI0/XI65/XI11/MM10_g N_VDD_XI0/XI65/XI11/MM10_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI11/MM11 N_XI0/XI65/XI11/NET36_XI0/XI65/XI11/MM11_d
+ N_XI0/XI65/XI11/NET35_XI0/XI65/XI11/MM11_g N_VDD_XI0/XI65/XI11/MM11_s
+ N_VDD_XI1/XI14/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI12/MM2 N_XI0/XI65/XI12/NET34_XI0/XI65/XI12/MM2_d
+ N_XI0/XI65/XI12/NET33_XI0/XI65/XI12/MM2_g N_VSS_XI0/XI65/XI12/MM2_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM3 N_XI0/XI65/XI12/NET33_XI0/XI65/XI12/MM3_d
+ N_WL<126>_XI0/XI65/XI12/MM3_g N_BLN<3>_XI0/XI65/XI12/MM3_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM0 N_XI0/XI65/XI12/NET34_XI0/XI65/XI12/MM0_d
+ N_WL<126>_XI0/XI65/XI12/MM0_g N_BL<3>_XI0/XI65/XI12/MM0_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM1 N_XI0/XI65/XI12/NET33_XI0/XI65/XI12/MM1_d
+ N_XI0/XI65/XI12/NET34_XI0/XI65/XI12/MM1_g N_VSS_XI0/XI65/XI12/MM1_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM9 N_XI0/XI65/XI12/NET36_XI0/XI65/XI12/MM9_d
+ N_WL<127>_XI0/XI65/XI12/MM9_g N_BL<3>_XI0/XI65/XI12/MM9_s N_VSS_XI1/XI14/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM6 N_XI0/XI65/XI12/NET35_XI0/XI65/XI12/MM6_d
+ N_XI0/XI65/XI12/NET36_XI0/XI65/XI12/MM6_g N_VSS_XI0/XI65/XI12/MM6_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM7 N_XI0/XI65/XI12/NET36_XI0/XI65/XI12/MM7_d
+ N_XI0/XI65/XI12/NET35_XI0/XI65/XI12/MM7_g N_VSS_XI0/XI65/XI12/MM7_s
+ N_VSS_XI1/XI14/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM8 N_XI0/XI65/XI12/NET35_XI0/XI65/XI12/MM8_d
+ N_WL<127>_XI0/XI65/XI12/MM8_g N_BLN<3>_XI0/XI65/XI12/MM8_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI12/MM5 N_XI0/XI65/XI12/NET34_XI0/XI65/XI12/MM5_d
+ N_XI0/XI65/XI12/NET33_XI0/XI65/XI12/MM5_g N_VDD_XI0/XI65/XI12/MM5_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI12/MM4 N_XI0/XI65/XI12/NET33_XI0/XI65/XI12/MM4_d
+ N_XI0/XI65/XI12/NET34_XI0/XI65/XI12/MM4_g N_VDD_XI0/XI65/XI12/MM4_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI12/MM10 N_XI0/XI65/XI12/NET35_XI0/XI65/XI12/MM10_d
+ N_XI0/XI65/XI12/NET36_XI0/XI65/XI12/MM10_g N_VDD_XI0/XI65/XI12/MM10_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI12/MM11 N_XI0/XI65/XI12/NET36_XI0/XI65/XI12/MM11_d
+ N_XI0/XI65/XI12/NET35_XI0/XI65/XI12/MM11_g N_VDD_XI0/XI65/XI12/MM11_s
+ N_VDD_XI1/XI3/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI13/MM2 N_XI0/XI65/XI13/NET34_XI0/XI65/XI13/MM2_d
+ N_XI0/XI65/XI13/NET33_XI0/XI65/XI13/MM2_g N_VSS_XI0/XI65/XI13/MM2_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM3 N_XI0/XI65/XI13/NET33_XI0/XI65/XI13/MM3_d
+ N_WL<126>_XI0/XI65/XI13/MM3_g N_BLN<2>_XI0/XI65/XI13/MM3_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM0 N_XI0/XI65/XI13/NET34_XI0/XI65/XI13/MM0_d
+ N_WL<126>_XI0/XI65/XI13/MM0_g N_BL<2>_XI0/XI65/XI13/MM0_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM1 N_XI0/XI65/XI13/NET33_XI0/XI65/XI13/MM1_d
+ N_XI0/XI65/XI13/NET34_XI0/XI65/XI13/MM1_g N_VSS_XI0/XI65/XI13/MM1_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM9 N_XI0/XI65/XI13/NET36_XI0/XI65/XI13/MM9_d
+ N_WL<127>_XI0/XI65/XI13/MM9_g N_BL<2>_XI0/XI65/XI13/MM9_s N_VSS_XI1/XI3/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM6 N_XI0/XI65/XI13/NET35_XI0/XI65/XI13/MM6_d
+ N_XI0/XI65/XI13/NET36_XI0/XI65/XI13/MM6_g N_VSS_XI0/XI65/XI13/MM6_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM7 N_XI0/XI65/XI13/NET36_XI0/XI65/XI13/MM7_d
+ N_XI0/XI65/XI13/NET35_XI0/XI65/XI13/MM7_g N_VSS_XI0/XI65/XI13/MM7_s
+ N_VSS_XI1/XI3/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM8 N_XI0/XI65/XI13/NET35_XI0/XI65/XI13/MM8_d
+ N_WL<127>_XI0/XI65/XI13/MM8_g N_BLN<2>_XI0/XI65/XI13/MM8_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI13/MM5 N_XI0/XI65/XI13/NET34_XI0/XI65/XI13/MM5_d
+ N_XI0/XI65/XI13/NET33_XI0/XI65/XI13/MM5_g N_VDD_XI0/XI65/XI13/MM5_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI13/MM4 N_XI0/XI65/XI13/NET33_XI0/XI65/XI13/MM4_d
+ N_XI0/XI65/XI13/NET34_XI0/XI65/XI13/MM4_g N_VDD_XI0/XI65/XI13/MM4_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI13/MM10 N_XI0/XI65/XI13/NET35_XI0/XI65/XI13/MM10_d
+ N_XI0/XI65/XI13/NET36_XI0/XI65/XI13/MM10_g N_VDD_XI0/XI65/XI13/MM10_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI13/MM11 N_XI0/XI65/XI13/NET36_XI0/XI65/XI13/MM11_d
+ N_XI0/XI65/XI13/NET35_XI0/XI65/XI13/MM11_g N_VDD_XI0/XI65/XI13/MM11_s
+ N_VDD_XI1/XI7/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI14/MM2 N_XI0/XI65/XI14/NET34_XI0/XI65/XI14/MM2_d
+ N_XI0/XI65/XI14/NET33_XI0/XI65/XI14/MM2_g N_VSS_XI0/XI65/XI14/MM2_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM3 N_XI0/XI65/XI14/NET33_XI0/XI65/XI14/MM3_d
+ N_WL<126>_XI0/XI65/XI14/MM3_g N_BLN<1>_XI0/XI65/XI14/MM3_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM0 N_XI0/XI65/XI14/NET34_XI0/XI65/XI14/MM0_d
+ N_WL<126>_XI0/XI65/XI14/MM0_g N_BL<1>_XI0/XI65/XI14/MM0_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM1 N_XI0/XI65/XI14/NET33_XI0/XI65/XI14/MM1_d
+ N_XI0/XI65/XI14/NET34_XI0/XI65/XI14/MM1_g N_VSS_XI0/XI65/XI14/MM1_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM9 N_XI0/XI65/XI14/NET36_XI0/XI65/XI14/MM9_d
+ N_WL<127>_XI0/XI65/XI14/MM9_g N_BL<1>_XI0/XI65/XI14/MM9_s N_VSS_XI1/XI7/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM6 N_XI0/XI65/XI14/NET35_XI0/XI65/XI14/MM6_d
+ N_XI0/XI65/XI14/NET36_XI0/XI65/XI14/MM6_g N_VSS_XI0/XI65/XI14/MM6_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM7 N_XI0/XI65/XI14/NET36_XI0/XI65/XI14/MM7_d
+ N_XI0/XI65/XI14/NET35_XI0/XI65/XI14/MM7_g N_VSS_XI0/XI65/XI14/MM7_s
+ N_VSS_XI1/XI7/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM8 N_XI0/XI65/XI14/NET35_XI0/XI65/XI14/MM8_d
+ N_WL<127>_XI0/XI65/XI14/MM8_g N_BLN<1>_XI0/XI65/XI14/MM8_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI14/MM5 N_XI0/XI65/XI14/NET34_XI0/XI65/XI14/MM5_d
+ N_XI0/XI65/XI14/NET33_XI0/XI65/XI14/MM5_g N_VDD_XI0/XI65/XI14/MM5_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI14/MM4 N_XI0/XI65/XI14/NET33_XI0/XI65/XI14/MM4_d
+ N_XI0/XI65/XI14/NET34_XI0/XI65/XI14/MM4_g N_VDD_XI0/XI65/XI14/MM4_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI14/MM10 N_XI0/XI65/XI14/NET35_XI0/XI65/XI14/MM10_d
+ N_XI0/XI65/XI14/NET36_XI0/XI65/XI14/MM10_g N_VDD_XI0/XI65/XI14/MM10_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI14/MM11 N_XI0/XI65/XI14/NET36_XI0/XI65/XI14/MM11_d
+ N_XI0/XI65/XI14/NET35_XI0/XI65/XI14/MM11_g N_VDD_XI0/XI65/XI14/MM11_s
+ N_VDD_XI1/XI11/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI15/MM2 N_XI0/XI65/XI15/NET34_XI0/XI65/XI15/MM2_d
+ N_XI0/XI65/XI15/NET33_XI0/XI65/XI15/MM2_g N_VSS_XI0/XI65/XI15/MM2_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM3 N_XI0/XI65/XI15/NET33_XI0/XI65/XI15/MM3_d
+ N_WL<126>_XI0/XI65/XI15/MM3_g N_BLN<0>_XI0/XI65/XI15/MM3_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM0 N_XI0/XI65/XI15/NET34_XI0/XI65/XI15/MM0_d
+ N_WL<126>_XI0/XI65/XI15/MM0_g N_BL<0>_XI0/XI65/XI15/MM0_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM1 N_XI0/XI65/XI15/NET33_XI0/XI65/XI15/MM1_d
+ N_XI0/XI65/XI15/NET34_XI0/XI65/XI15/MM1_g N_VSS_XI0/XI65/XI15/MM1_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM9 N_XI0/XI65/XI15/NET36_XI0/XI65/XI15/MM9_d
+ N_WL<127>_XI0/XI65/XI15/MM9_g N_BL<0>_XI0/XI65/XI15/MM9_s N_VSS_XI1/XI11/MM1_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM6 N_XI0/XI65/XI15/NET35_XI0/XI65/XI15/MM6_d
+ N_XI0/XI65/XI15/NET36_XI0/XI65/XI15/MM6_g N_VSS_XI0/XI65/XI15/MM6_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM7 N_XI0/XI65/XI15/NET36_XI0/XI65/XI15/MM7_d
+ N_XI0/XI65/XI15/NET35_XI0/XI65/XI15/MM7_g N_VSS_XI0/XI65/XI15/MM7_s
+ N_VSS_XI1/XI11/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM8 N_XI0/XI65/XI15/NET35_XI0/XI65/XI15/MM8_d
+ N_WL<127>_XI0/XI65/XI15/MM8_g N_BLN<0>_XI0/XI65/XI15/MM8_s
+ N_VSS_XI1/XI15/MM1_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI65/XI15/MM5 N_XI0/XI65/XI15/NET34_XI0/XI65/XI15/MM5_d
+ N_XI0/XI65/XI15/NET33_XI0/XI65/XI15/MM5_g N_VDD_XI0/XI65/XI15/MM5_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI15/MM4 N_XI0/XI65/XI15/NET33_XI0/XI65/XI15/MM4_d
+ N_XI0/XI65/XI15/NET34_XI0/XI65/XI15/MM4_g N_VDD_XI0/XI65/XI15/MM4_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI15/MM10 N_XI0/XI65/XI15/NET35_XI0/XI65/XI15/MM10_d
+ N_XI0/XI65/XI15/NET36_XI0/XI65/XI15/MM10_g N_VDD_XI0/XI65/XI15/MM10_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI65/XI15/MM11 N_XI0/XI65/XI15/NET36_XI0/XI65/XI15/MM11_d
+ N_XI0/XI65/XI15/NET35_XI0/XI65/XI15/MM11_g N_VDD_XI0/XI65/XI15/MM11_s
+ N_VDD_XI1/XI15/MM6_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
*
.include "netlist.sp.SRAMNSA_1.pxi"
*
.ends
*
*
