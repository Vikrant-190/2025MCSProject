* File: netlist.sp
* Created: Fri Jun 13 14:32:41 2025
* Program "Calibre xRC"
* Version "v2019.2_26.18"
* 
.include "netlist.sp.pex"
.subckt sram_array_1  VSS BL<15> VDD BLN<15> BL<14> BLN<14> BL<13> BLN<13>
+ BL<12> BLN<12> BL<11> BLN<11> BL<10> BLN<10> BL<9> BLN<9> BL<8> BLN<8> BL<7>
+ BLN<7> BL<6> BLN<6> BL<5> BLN<5> BL<4> BLN<4> BL<3> BLN<3> BL<2> BLN<2> BL<1>
+ BLN<1> BL<0> BLN<0> WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> WL<6> WL<7> WL<8>
+ WL<9> WL<10> WL<11> WL<12> WL<13> WL<14> WL<15> WL<16> WL<17> WL<18> WL<19>
+ WL<20> WL<21> WL<22> WL<23> WL<24> WL<25> WL<26> WL<27> WL<28> WL<29> WL<30>
+ WL<31> WL<32> WL<33> WL<34> WL<35> WL<36> WL<37> WL<38> WL<39> WL<40> WL<41>
+ WL<42> WL<43> WL<44> WL<45> WL<46> WL<47> WL<48> WL<49> WL<50> WL<51> WL<52>
+ WL<53> WL<54> WL<55> WL<56> WL<57> WL<58> WL<59> WL<60> WL<61> WL<62> WL<63>
+ WL<64> WL<65> WL<66> WL<67> WL<68> WL<69> WL<70> WL<71> WL<72> WL<73> WL<74>
+ WL<75> WL<76> WL<77> WL<78> WL<79> WL<80> WL<81> WL<82> WL<83> WL<84> WL<85>
+ WL<86> WL<87> WL<88> WL<89> WL<90> WL<91> WL<92> WL<93> WL<94> WL<95> WL<96>
+ WL<97> WL<98> WL<99> WL<100> WL<101> WL<102> WL<103> WL<104> WL<105> WL<106>
+ WL<107> WL<108> WL<109> WL<110> WL<111> WL<112> WL<113> WL<114> WL<115>
+ WL<116> WL<117> WL<118> WL<119> WL<120> WL<121> WL<122> WL<123> WL<124>
+ WL<125> WL<126> WL<127>
* 
* WL<127>	WL<127>
* WL<126>	WL<126>
* WL<125>	WL<125>
* WL<124>	WL<124>
* WL<123>	WL<123>
* WL<122>	WL<122>
* WL<121>	WL<121>
* WL<120>	WL<120>
* WL<119>	WL<119>
* WL<118>	WL<118>
* WL<117>	WL<117>
* WL<116>	WL<116>
* WL<115>	WL<115>
* WL<114>	WL<114>
* WL<113>	WL<113>
* WL<112>	WL<112>
* WL<111>	WL<111>
* WL<110>	WL<110>
* WL<109>	WL<109>
* WL<108>	WL<108>
* WL<107>	WL<107>
* WL<106>	WL<106>
* WL<105>	WL<105>
* WL<104>	WL<104>
* WL<103>	WL<103>
* WL<102>	WL<102>
* WL<101>	WL<101>
* WL<100>	WL<100>
* WL<99>	WL<99>
* WL<98>	WL<98>
* WL<97>	WL<97>
* WL<96>	WL<96>
* WL<95>	WL<95>
* WL<94>	WL<94>
* WL<93>	WL<93>
* WL<92>	WL<92>
* WL<91>	WL<91>
* WL<90>	WL<90>
* WL<89>	WL<89>
* WL<88>	WL<88>
* WL<87>	WL<87>
* WL<86>	WL<86>
* WL<85>	WL<85>
* WL<84>	WL<84>
* WL<83>	WL<83>
* WL<82>	WL<82>
* WL<81>	WL<81>
* WL<80>	WL<80>
* WL<79>	WL<79>
* WL<78>	WL<78>
* WL<77>	WL<77>
* WL<76>	WL<76>
* WL<75>	WL<75>
* WL<74>	WL<74>
* WL<73>	WL<73>
* WL<72>	WL<72>
* WL<71>	WL<71>
* WL<70>	WL<70>
* WL<69>	WL<69>
* WL<68>	WL<68>
* WL<67>	WL<67>
* WL<66>	WL<66>
* WL<65>	WL<65>
* WL<64>	WL<64>
* WL<63>	WL<63>
* WL<62>	WL<62>
* WL<61>	WL<61>
* WL<60>	WL<60>
* WL<59>	WL<59>
* WL<58>	WL<58>
* WL<57>	WL<57>
* WL<56>	WL<56>
* WL<55>	WL<55>
* WL<54>	WL<54>
* WL<53>	WL<53>
* WL<52>	WL<52>
* WL<51>	WL<51>
* WL<50>	WL<50>
* WL<49>	WL<49>
* WL<48>	WL<48>
* WL<47>	WL<47>
* WL<46>	WL<46>
* WL<45>	WL<45>
* WL<44>	WL<44>
* WL<43>	WL<43>
* WL<42>	WL<42>
* WL<41>	WL<41>
* WL<40>	WL<40>
* WL<39>	WL<39>
* WL<38>	WL<38>
* WL<37>	WL<37>
* WL<36>	WL<36>
* WL<35>	WL<35>
* WL<34>	WL<34>
* WL<33>	WL<33>
* WL<32>	WL<32>
* WL<31>	WL<31>
* WL<30>	WL<30>
* WL<29>	WL<29>
* WL<28>	WL<28>
* WL<27>	WL<27>
* WL<26>	WL<26>
* WL<25>	WL<25>
* WL<24>	WL<24>
* WL<23>	WL<23>
* WL<22>	WL<22>
* WL<21>	WL<21>
* WL<20>	WL<20>
* WL<19>	WL<19>
* WL<18>	WL<18>
* WL<17>	WL<17>
* WL<16>	WL<16>
* WL<15>	WL<15>
* WL<14>	WL<14>
* WL<13>	WL<13>
* WL<12>	WL<12>
* WL<11>	WL<11>
* WL<10>	WL<10>
* WL<9>	WL<9>
* WL<8>	WL<8>
* WL<7>	WL<7>
* WL<6>	WL<6>
* WL<5>	WL<5>
* WL<4>	WL<4>
* WL<3>	WL<3>
* WL<2>	WL<2>
* WL<1>	WL<1>
* WL<0>	WL<0>
* BLN<0>	BLN<0>
* BL<0>	BL<0>
* BLN<1>	BLN<1>
* BL<1>	BL<1>
* BLN<2>	BLN<2>
* BL<2>	BL<2>
* BLN<3>	BLN<3>
* BL<3>	BL<3>
* BLN<4>	BLN<4>
* BL<4>	BL<4>
* BLN<5>	BLN<5>
* BL<5>	BL<5>
* BLN<6>	BLN<6>
* BL<6>	BL<6>
* BLN<7>	BLN<7>
* BL<7>	BL<7>
* BLN<8>	BLN<8>
* BL<8>	BL<8>
* BLN<9>	BLN<9>
* BL<9>	BL<9>
* BLN<10>	BLN<10>
* BL<10>	BL<10>
* BLN<11>	BLN<11>
* BL<11>	BL<11>
* BLN<12>	BLN<12>
* BL<12>	BL<12>
* BLN<13>	BLN<13>
* BL<13>	BL<13>
* BLN<14>	BLN<14>
* BL<14>	BL<14>
* BLN<15>	BLN<15>
* VDD	VDD
* BL<15>	BL<15>
* VSS	VSS
mXI0/XI0/MM2 N_XI0/XI0/NET34_XI0/XI0/MM2_d N_XI0/XI0/NET33_XI0/XI0/MM2_g
+ N_VSS_XI0/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM3 N_XI0/XI0/NET33_XI0/XI0/MM3_d N_WL<0>_XI0/XI0/MM3_g
+ N_BLN<15>_XI0/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM0 N_XI0/XI0/NET34_XI0/XI0/MM0_d N_WL<0>_XI0/XI0/MM0_g
+ N_BL<15>_XI0/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM1 N_XI0/XI0/NET33_XI0/XI0/MM1_d N_XI0/XI0/NET34_XI0/XI0/MM1_g
+ N_VSS_XI0/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM9 N_XI0/XI0/NET36_XI0/XI0/MM9_d N_WL<1>_XI0/XI0/MM9_g
+ N_BL<15>_XI0/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM6 N_XI0/XI0/NET35_XI0/XI0/MM6_d N_XI0/XI0/NET36_XI0/XI0/MM6_g
+ N_VSS_XI0/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM7 N_XI0/XI0/NET36_XI0/XI0/MM7_d N_XI0/XI0/NET35_XI0/XI0/MM7_g
+ N_VSS_XI0/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM8 N_XI0/XI0/NET35_XI0/XI0/MM8_d N_WL<1>_XI0/XI0/MM8_g
+ N_BLN<15>_XI0/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI0/MM5 N_XI0/XI0/NET34_XI0/XI0/MM5_d N_XI0/XI0/NET33_XI0/XI0/MM5_g
+ N_VDD_XI0/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/MM4 N_XI0/XI0/NET33_XI0/XI0/MM4_d N_XI0/XI0/NET34_XI0/XI0/MM4_g
+ N_VDD_XI0/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/MM10 N_XI0/XI0/NET35_XI0/XI0/MM10_d N_XI0/XI0/NET36_XI0/XI0/MM10_g
+ N_VDD_XI0/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI0/MM11 N_XI0/XI0/NET36_XI0/XI0/MM11_d N_XI0/XI0/NET35_XI0/XI0/MM11_g
+ N_VDD_XI0/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/MM2 N_XI0/XI1/NET34_XI0/XI1/MM2_d N_XI0/XI1/NET33_XI0/XI1/MM2_g
+ N_VSS_XI0/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM3 N_XI0/XI1/NET33_XI0/XI1/MM3_d N_WL<0>_XI0/XI1/MM3_g
+ N_BLN<14>_XI0/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM0 N_XI0/XI1/NET34_XI0/XI1/MM0_d N_WL<0>_XI0/XI1/MM0_g
+ N_BL<14>_XI0/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM1 N_XI0/XI1/NET33_XI0/XI1/MM1_d N_XI0/XI1/NET34_XI0/XI1/MM1_g
+ N_VSS_XI0/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM9 N_XI0/XI1/NET36_XI0/XI1/MM9_d N_WL<1>_XI0/XI1/MM9_g
+ N_BL<14>_XI0/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM6 N_XI0/XI1/NET35_XI0/XI1/MM6_d N_XI0/XI1/NET36_XI0/XI1/MM6_g
+ N_VSS_XI0/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM7 N_XI0/XI1/NET36_XI0/XI1/MM7_d N_XI0/XI1/NET35_XI0/XI1/MM7_g
+ N_VSS_XI0/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM8 N_XI0/XI1/NET35_XI0/XI1/MM8_d N_WL<1>_XI0/XI1/MM8_g
+ N_BLN<14>_XI0/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI1/MM5 N_XI0/XI1/NET34_XI0/XI1/MM5_d N_XI0/XI1/NET33_XI0/XI1/MM5_g
+ N_VDD_XI0/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/MM4 N_XI0/XI1/NET33_XI0/XI1/MM4_d N_XI0/XI1/NET34_XI0/XI1/MM4_g
+ N_VDD_XI0/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/MM10 N_XI0/XI1/NET35_XI0/XI1/MM10_d N_XI0/XI1/NET36_XI0/XI1/MM10_g
+ N_VDD_XI0/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI1/MM11 N_XI0/XI1/NET36_XI0/XI1/MM11_d N_XI0/XI1/NET35_XI0/XI1/MM11_g
+ N_VDD_XI0/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI2/MM2 N_XI0/XI2/NET34_XI0/XI2/MM2_d N_XI0/XI2/NET33_XI0/XI2/MM2_g
+ N_VSS_XI0/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM3 N_XI0/XI2/NET33_XI0/XI2/MM3_d N_WL<0>_XI0/XI2/MM3_g
+ N_BLN<13>_XI0/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM0 N_XI0/XI2/NET34_XI0/XI2/MM0_d N_WL<0>_XI0/XI2/MM0_g
+ N_BL<13>_XI0/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM1 N_XI0/XI2/NET33_XI0/XI2/MM1_d N_XI0/XI2/NET34_XI0/XI2/MM1_g
+ N_VSS_XI0/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM9 N_XI0/XI2/NET36_XI0/XI2/MM9_d N_WL<1>_XI0/XI2/MM9_g
+ N_BL<13>_XI0/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM6 N_XI0/XI2/NET35_XI0/XI2/MM6_d N_XI0/XI2/NET36_XI0/XI2/MM6_g
+ N_VSS_XI0/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM7 N_XI0/XI2/NET36_XI0/XI2/MM7_d N_XI0/XI2/NET35_XI0/XI2/MM7_g
+ N_VSS_XI0/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM8 N_XI0/XI2/NET35_XI0/XI2/MM8_d N_WL<1>_XI0/XI2/MM8_g
+ N_BLN<13>_XI0/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI2/MM5 N_XI0/XI2/NET34_XI0/XI2/MM5_d N_XI0/XI2/NET33_XI0/XI2/MM5_g
+ N_VDD_XI0/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI2/MM4 N_XI0/XI2/NET33_XI0/XI2/MM4_d N_XI0/XI2/NET34_XI0/XI2/MM4_g
+ N_VDD_XI0/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI2/MM10 N_XI0/XI2/NET35_XI0/XI2/MM10_d N_XI0/XI2/NET36_XI0/XI2/MM10_g
+ N_VDD_XI0/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI2/MM11 N_XI0/XI2/NET36_XI0/XI2/MM11_d N_XI0/XI2/NET35_XI0/XI2/MM11_g
+ N_VDD_XI0/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI3/MM2 N_XI0/XI3/NET34_XI0/XI3/MM2_d N_XI0/XI3/NET33_XI0/XI3/MM2_g
+ N_VSS_XI0/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM3 N_XI0/XI3/NET33_XI0/XI3/MM3_d N_WL<0>_XI0/XI3/MM3_g
+ N_BLN<12>_XI0/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM0 N_XI0/XI3/NET34_XI0/XI3/MM0_d N_WL<0>_XI0/XI3/MM0_g
+ N_BL<12>_XI0/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM1 N_XI0/XI3/NET33_XI0/XI3/MM1_d N_XI0/XI3/NET34_XI0/XI3/MM1_g
+ N_VSS_XI0/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM9 N_XI0/XI3/NET36_XI0/XI3/MM9_d N_WL<1>_XI0/XI3/MM9_g
+ N_BL<12>_XI0/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM6 N_XI0/XI3/NET35_XI0/XI3/MM6_d N_XI0/XI3/NET36_XI0/XI3/MM6_g
+ N_VSS_XI0/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM7 N_XI0/XI3/NET36_XI0/XI3/MM7_d N_XI0/XI3/NET35_XI0/XI3/MM7_g
+ N_VSS_XI0/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM8 N_XI0/XI3/NET35_XI0/XI3/MM8_d N_WL<1>_XI0/XI3/MM8_g
+ N_BLN<12>_XI0/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI3/MM5 N_XI0/XI3/NET34_XI0/XI3/MM5_d N_XI0/XI3/NET33_XI0/XI3/MM5_g
+ N_VDD_XI0/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI3/MM4 N_XI0/XI3/NET33_XI0/XI3/MM4_d N_XI0/XI3/NET34_XI0/XI3/MM4_g
+ N_VDD_XI0/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI3/MM10 N_XI0/XI3/NET35_XI0/XI3/MM10_d N_XI0/XI3/NET36_XI0/XI3/MM10_g
+ N_VDD_XI0/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI3/MM11 N_XI0/XI3/NET36_XI0/XI3/MM11_d N_XI0/XI3/NET35_XI0/XI3/MM11_g
+ N_VDD_XI0/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/MM2 N_XI0/XI4/NET34_XI0/XI4/MM2_d N_XI0/XI4/NET33_XI0/XI4/MM2_g
+ N_VSS_XI0/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM3 N_XI0/XI4/NET33_XI0/XI4/MM3_d N_WL<0>_XI0/XI4/MM3_g
+ N_BLN<11>_XI0/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM0 N_XI0/XI4/NET34_XI0/XI4/MM0_d N_WL<0>_XI0/XI4/MM0_g
+ N_BL<11>_XI0/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM1 N_XI0/XI4/NET33_XI0/XI4/MM1_d N_XI0/XI4/NET34_XI0/XI4/MM1_g
+ N_VSS_XI0/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM9 N_XI0/XI4/NET36_XI0/XI4/MM9_d N_WL<1>_XI0/XI4/MM9_g
+ N_BL<11>_XI0/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM6 N_XI0/XI4/NET35_XI0/XI4/MM6_d N_XI0/XI4/NET36_XI0/XI4/MM6_g
+ N_VSS_XI0/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM7 N_XI0/XI4/NET36_XI0/XI4/MM7_d N_XI0/XI4/NET35_XI0/XI4/MM7_g
+ N_VSS_XI0/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM8 N_XI0/XI4/NET35_XI0/XI4/MM8_d N_WL<1>_XI0/XI4/MM8_g
+ N_BLN<11>_XI0/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI4/MM5 N_XI0/XI4/NET34_XI0/XI4/MM5_d N_XI0/XI4/NET33_XI0/XI4/MM5_g
+ N_VDD_XI0/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/MM4 N_XI0/XI4/NET33_XI0/XI4/MM4_d N_XI0/XI4/NET34_XI0/XI4/MM4_g
+ N_VDD_XI0/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/MM10 N_XI0/XI4/NET35_XI0/XI4/MM10_d N_XI0/XI4/NET36_XI0/XI4/MM10_g
+ N_VDD_XI0/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI4/MM11 N_XI0/XI4/NET36_XI0/XI4/MM11_d N_XI0/XI4/NET35_XI0/XI4/MM11_g
+ N_VDD_XI0/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/MM2 N_XI0/XI5/NET34_XI0/XI5/MM2_d N_XI0/XI5/NET33_XI0/XI5/MM2_g
+ N_VSS_XI0/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM3 N_XI0/XI5/NET33_XI0/XI5/MM3_d N_WL<0>_XI0/XI5/MM3_g
+ N_BLN<10>_XI0/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM0 N_XI0/XI5/NET34_XI0/XI5/MM0_d N_WL<0>_XI0/XI5/MM0_g
+ N_BL<10>_XI0/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM1 N_XI0/XI5/NET33_XI0/XI5/MM1_d N_XI0/XI5/NET34_XI0/XI5/MM1_g
+ N_VSS_XI0/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM9 N_XI0/XI5/NET36_XI0/XI5/MM9_d N_WL<1>_XI0/XI5/MM9_g
+ N_BL<10>_XI0/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM6 N_XI0/XI5/NET35_XI0/XI5/MM6_d N_XI0/XI5/NET36_XI0/XI5/MM6_g
+ N_VSS_XI0/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM7 N_XI0/XI5/NET36_XI0/XI5/MM7_d N_XI0/XI5/NET35_XI0/XI5/MM7_g
+ N_VSS_XI0/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM8 N_XI0/XI5/NET35_XI0/XI5/MM8_d N_WL<1>_XI0/XI5/MM8_g
+ N_BLN<10>_XI0/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI5/MM5 N_XI0/XI5/NET34_XI0/XI5/MM5_d N_XI0/XI5/NET33_XI0/XI5/MM5_g
+ N_VDD_XI0/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/MM4 N_XI0/XI5/NET33_XI0/XI5/MM4_d N_XI0/XI5/NET34_XI0/XI5/MM4_g
+ N_VDD_XI0/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/MM10 N_XI0/XI5/NET35_XI0/XI5/MM10_d N_XI0/XI5/NET36_XI0/XI5/MM10_g
+ N_VDD_XI0/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI5/MM11 N_XI0/XI5/NET36_XI0/XI5/MM11_d N_XI0/XI5/NET35_XI0/XI5/MM11_g
+ N_VDD_XI0/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/MM2 N_XI0/XI6/NET34_XI0/XI6/MM2_d N_XI0/XI6/NET33_XI0/XI6/MM2_g
+ N_VSS_XI0/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM3 N_XI0/XI6/NET33_XI0/XI6/MM3_d N_WL<0>_XI0/XI6/MM3_g
+ N_BLN<9>_XI0/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM0 N_XI0/XI6/NET34_XI0/XI6/MM0_d N_WL<0>_XI0/XI6/MM0_g
+ N_BL<9>_XI0/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM1 N_XI0/XI6/NET33_XI0/XI6/MM1_d N_XI0/XI6/NET34_XI0/XI6/MM1_g
+ N_VSS_XI0/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM9 N_XI0/XI6/NET36_XI0/XI6/MM9_d N_WL<1>_XI0/XI6/MM9_g
+ N_BL<9>_XI0/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM6 N_XI0/XI6/NET35_XI0/XI6/MM6_d N_XI0/XI6/NET36_XI0/XI6/MM6_g
+ N_VSS_XI0/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM7 N_XI0/XI6/NET36_XI0/XI6/MM7_d N_XI0/XI6/NET35_XI0/XI6/MM7_g
+ N_VSS_XI0/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM8 N_XI0/XI6/NET35_XI0/XI6/MM8_d N_WL<1>_XI0/XI6/MM8_g
+ N_BLN<9>_XI0/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI6/MM5 N_XI0/XI6/NET34_XI0/XI6/MM5_d N_XI0/XI6/NET33_XI0/XI6/MM5_g
+ N_VDD_XI0/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/MM4 N_XI0/XI6/NET33_XI0/XI6/MM4_d N_XI0/XI6/NET34_XI0/XI6/MM4_g
+ N_VDD_XI0/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/MM10 N_XI0/XI6/NET35_XI0/XI6/MM10_d N_XI0/XI6/NET36_XI0/XI6/MM10_g
+ N_VDD_XI0/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI6/MM11 N_XI0/XI6/NET36_XI0/XI6/MM11_d N_XI0/XI6/NET35_XI0/XI6/MM11_g
+ N_VDD_XI0/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/MM2 N_XI0/XI7/NET34_XI0/XI7/MM2_d N_XI0/XI7/NET33_XI0/XI7/MM2_g
+ N_VSS_XI0/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM3 N_XI0/XI7/NET33_XI0/XI7/MM3_d N_WL<0>_XI0/XI7/MM3_g
+ N_BLN<8>_XI0/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM0 N_XI0/XI7/NET34_XI0/XI7/MM0_d N_WL<0>_XI0/XI7/MM0_g
+ N_BL<8>_XI0/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM1 N_XI0/XI7/NET33_XI0/XI7/MM1_d N_XI0/XI7/NET34_XI0/XI7/MM1_g
+ N_VSS_XI0/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM9 N_XI0/XI7/NET36_XI0/XI7/MM9_d N_WL<1>_XI0/XI7/MM9_g
+ N_BL<8>_XI0/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM6 N_XI0/XI7/NET35_XI0/XI7/MM6_d N_XI0/XI7/NET36_XI0/XI7/MM6_g
+ N_VSS_XI0/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM7 N_XI0/XI7/NET36_XI0/XI7/MM7_d N_XI0/XI7/NET35_XI0/XI7/MM7_g
+ N_VSS_XI0/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM8 N_XI0/XI7/NET35_XI0/XI7/MM8_d N_WL<1>_XI0/XI7/MM8_g
+ N_BLN<8>_XI0/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI7/MM5 N_XI0/XI7/NET34_XI0/XI7/MM5_d N_XI0/XI7/NET33_XI0/XI7/MM5_g
+ N_VDD_XI0/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/MM4 N_XI0/XI7/NET33_XI0/XI7/MM4_d N_XI0/XI7/NET34_XI0/XI7/MM4_g
+ N_VDD_XI0/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/MM10 N_XI0/XI7/NET35_XI0/XI7/MM10_d N_XI0/XI7/NET36_XI0/XI7/MM10_g
+ N_VDD_XI0/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI7/MM11 N_XI0/XI7/NET36_XI0/XI7/MM11_d N_XI0/XI7/NET35_XI0/XI7/MM11_g
+ N_VDD_XI0/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/MM2 N_XI0/XI8/NET34_XI0/XI8/MM2_d N_XI0/XI8/NET33_XI0/XI8/MM2_g
+ N_VSS_XI0/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM3 N_XI0/XI8/NET33_XI0/XI8/MM3_d N_WL<0>_XI0/XI8/MM3_g
+ N_BLN<7>_XI0/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM0 N_XI0/XI8/NET34_XI0/XI8/MM0_d N_WL<0>_XI0/XI8/MM0_g
+ N_BL<7>_XI0/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM1 N_XI0/XI8/NET33_XI0/XI8/MM1_d N_XI0/XI8/NET34_XI0/XI8/MM1_g
+ N_VSS_XI0/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM9 N_XI0/XI8/NET36_XI0/XI8/MM9_d N_WL<1>_XI0/XI8/MM9_g
+ N_BL<7>_XI0/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM6 N_XI0/XI8/NET35_XI0/XI8/MM6_d N_XI0/XI8/NET36_XI0/XI8/MM6_g
+ N_VSS_XI0/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM7 N_XI0/XI8/NET36_XI0/XI8/MM7_d N_XI0/XI8/NET35_XI0/XI8/MM7_g
+ N_VSS_XI0/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM8 N_XI0/XI8/NET35_XI0/XI8/MM8_d N_WL<1>_XI0/XI8/MM8_g
+ N_BLN<7>_XI0/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI8/MM5 N_XI0/XI8/NET34_XI0/XI8/MM5_d N_XI0/XI8/NET33_XI0/XI8/MM5_g
+ N_VDD_XI0/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/MM4 N_XI0/XI8/NET33_XI0/XI8/MM4_d N_XI0/XI8/NET34_XI0/XI8/MM4_g
+ N_VDD_XI0/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/MM10 N_XI0/XI8/NET35_XI0/XI8/MM10_d N_XI0/XI8/NET36_XI0/XI8/MM10_g
+ N_VDD_XI0/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI8/MM11 N_XI0/XI8/NET36_XI0/XI8/MM11_d N_XI0/XI8/NET35_XI0/XI8/MM11_g
+ N_VDD_XI0/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/MM2 N_XI0/XI9/NET34_XI0/XI9/MM2_d N_XI0/XI9/NET33_XI0/XI9/MM2_g
+ N_VSS_XI0/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM3 N_XI0/XI9/NET33_XI0/XI9/MM3_d N_WL<0>_XI0/XI9/MM3_g
+ N_BLN<6>_XI0/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM0 N_XI0/XI9/NET34_XI0/XI9/MM0_d N_WL<0>_XI0/XI9/MM0_g
+ N_BL<6>_XI0/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM1 N_XI0/XI9/NET33_XI0/XI9/MM1_d N_XI0/XI9/NET34_XI0/XI9/MM1_g
+ N_VSS_XI0/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM9 N_XI0/XI9/NET36_XI0/XI9/MM9_d N_WL<1>_XI0/XI9/MM9_g
+ N_BL<6>_XI0/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM6 N_XI0/XI9/NET35_XI0/XI9/MM6_d N_XI0/XI9/NET36_XI0/XI9/MM6_g
+ N_VSS_XI0/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM7 N_XI0/XI9/NET36_XI0/XI9/MM7_d N_XI0/XI9/NET35_XI0/XI9/MM7_g
+ N_VSS_XI0/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM8 N_XI0/XI9/NET35_XI0/XI9/MM8_d N_WL<1>_XI0/XI9/MM8_g
+ N_BLN<6>_XI0/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI9/MM5 N_XI0/XI9/NET34_XI0/XI9/MM5_d N_XI0/XI9/NET33_XI0/XI9/MM5_g
+ N_VDD_XI0/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/MM4 N_XI0/XI9/NET33_XI0/XI9/MM4_d N_XI0/XI9/NET34_XI0/XI9/MM4_g
+ N_VDD_XI0/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/MM10 N_XI0/XI9/NET35_XI0/XI9/MM10_d N_XI0/XI9/NET36_XI0/XI9/MM10_g
+ N_VDD_XI0/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI9/MM11 N_XI0/XI9/NET36_XI0/XI9/MM11_d N_XI0/XI9/NET35_XI0/XI9/MM11_g
+ N_VDD_XI0/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/MM2 N_XI0/XI10/NET34_XI0/XI10/MM2_d N_XI0/XI10/NET33_XI0/XI10/MM2_g
+ N_VSS_XI0/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/MM3 N_XI0/XI10/NET33_XI0/XI10/MM3_d N_WL<0>_XI0/XI10/MM3_g
+ N_BLN<5>_XI0/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI10/MM0 N_XI0/XI10/NET34_XI0/XI10/MM0_d N_WL<0>_XI0/XI10/MM0_g
+ N_BL<5>_XI0/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/MM1 N_XI0/XI10/NET33_XI0/XI10/MM1_d N_XI0/XI10/NET34_XI0/XI10/MM1_g
+ N_VSS_XI0/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/MM9 N_XI0/XI10/NET36_XI0/XI10/MM9_d N_WL<1>_XI0/XI10/MM9_g
+ N_BL<5>_XI0/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/MM6 N_XI0/XI10/NET35_XI0/XI10/MM6_d N_XI0/XI10/NET36_XI0/XI10/MM6_g
+ N_VSS_XI0/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/MM7 N_XI0/XI10/NET36_XI0/XI10/MM7_d N_XI0/XI10/NET35_XI0/XI10/MM7_g
+ N_VSS_XI0/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI10/MM8 N_XI0/XI10/NET35_XI0/XI10/MM8_d N_WL<1>_XI0/XI10/MM8_g
+ N_BLN<5>_XI0/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI10/MM5 N_XI0/XI10/NET34_XI0/XI10/MM5_d N_XI0/XI10/NET33_XI0/XI10/MM5_g
+ N_VDD_XI0/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/MM4 N_XI0/XI10/NET33_XI0/XI10/MM4_d N_XI0/XI10/NET34_XI0/XI10/MM4_g
+ N_VDD_XI0/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/MM10 N_XI0/XI10/NET35_XI0/XI10/MM10_d N_XI0/XI10/NET36_XI0/XI10/MM10_g
+ N_VDD_XI0/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI10/MM11 N_XI0/XI10/NET36_XI0/XI10/MM11_d N_XI0/XI10/NET35_XI0/XI10/MM11_g
+ N_VDD_XI0/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/MM2 N_XI0/XI11/NET34_XI0/XI11/MM2_d N_XI0/XI11/NET33_XI0/XI11/MM2_g
+ N_VSS_XI0/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/MM3 N_XI0/XI11/NET33_XI0/XI11/MM3_d N_WL<0>_XI0/XI11/MM3_g
+ N_BLN<4>_XI0/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI11/MM0 N_XI0/XI11/NET34_XI0/XI11/MM0_d N_WL<0>_XI0/XI11/MM0_g
+ N_BL<4>_XI0/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/MM1 N_XI0/XI11/NET33_XI0/XI11/MM1_d N_XI0/XI11/NET34_XI0/XI11/MM1_g
+ N_VSS_XI0/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/MM9 N_XI0/XI11/NET36_XI0/XI11/MM9_d N_WL<1>_XI0/XI11/MM9_g
+ N_BL<4>_XI0/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/MM6 N_XI0/XI11/NET35_XI0/XI11/MM6_d N_XI0/XI11/NET36_XI0/XI11/MM6_g
+ N_VSS_XI0/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/MM7 N_XI0/XI11/NET36_XI0/XI11/MM7_d N_XI0/XI11/NET35_XI0/XI11/MM7_g
+ N_VSS_XI0/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI11/MM8 N_XI0/XI11/NET35_XI0/XI11/MM8_d N_WL<1>_XI0/XI11/MM8_g
+ N_BLN<4>_XI0/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI11/MM5 N_XI0/XI11/NET34_XI0/XI11/MM5_d N_XI0/XI11/NET33_XI0/XI11/MM5_g
+ N_VDD_XI0/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/MM4 N_XI0/XI11/NET33_XI0/XI11/MM4_d N_XI0/XI11/NET34_XI0/XI11/MM4_g
+ N_VDD_XI0/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/MM10 N_XI0/XI11/NET35_XI0/XI11/MM10_d N_XI0/XI11/NET36_XI0/XI11/MM10_g
+ N_VDD_XI0/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI11/MM11 N_XI0/XI11/NET36_XI0/XI11/MM11_d N_XI0/XI11/NET35_XI0/XI11/MM11_g
+ N_VDD_XI0/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/MM2 N_XI0/XI12/NET34_XI0/XI12/MM2_d N_XI0/XI12/NET33_XI0/XI12/MM2_g
+ N_VSS_XI0/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/MM3 N_XI0/XI12/NET33_XI0/XI12/MM3_d N_WL<0>_XI0/XI12/MM3_g
+ N_BLN<3>_XI0/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI12/MM0 N_XI0/XI12/NET34_XI0/XI12/MM0_d N_WL<0>_XI0/XI12/MM0_g
+ N_BL<3>_XI0/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/MM1 N_XI0/XI12/NET33_XI0/XI12/MM1_d N_XI0/XI12/NET34_XI0/XI12/MM1_g
+ N_VSS_XI0/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/MM9 N_XI0/XI12/NET36_XI0/XI12/MM9_d N_WL<1>_XI0/XI12/MM9_g
+ N_BL<3>_XI0/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/MM6 N_XI0/XI12/NET35_XI0/XI12/MM6_d N_XI0/XI12/NET36_XI0/XI12/MM6_g
+ N_VSS_XI0/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/MM7 N_XI0/XI12/NET36_XI0/XI12/MM7_d N_XI0/XI12/NET35_XI0/XI12/MM7_g
+ N_VSS_XI0/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI12/MM8 N_XI0/XI12/NET35_XI0/XI12/MM8_d N_WL<1>_XI0/XI12/MM8_g
+ N_BLN<3>_XI0/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI12/MM5 N_XI0/XI12/NET34_XI0/XI12/MM5_d N_XI0/XI12/NET33_XI0/XI12/MM5_g
+ N_VDD_XI0/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/MM4 N_XI0/XI12/NET33_XI0/XI12/MM4_d N_XI0/XI12/NET34_XI0/XI12/MM4_g
+ N_VDD_XI0/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/MM10 N_XI0/XI12/NET35_XI0/XI12/MM10_d N_XI0/XI12/NET36_XI0/XI12/MM10_g
+ N_VDD_XI0/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI12/MM11 N_XI0/XI12/NET36_XI0/XI12/MM11_d N_XI0/XI12/NET35_XI0/XI12/MM11_g
+ N_VDD_XI0/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/MM2 N_XI0/XI13/NET34_XI0/XI13/MM2_d N_XI0/XI13/NET33_XI0/XI13/MM2_g
+ N_VSS_XI0/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/MM3 N_XI0/XI13/NET33_XI0/XI13/MM3_d N_WL<0>_XI0/XI13/MM3_g
+ N_BLN<2>_XI0/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI13/MM0 N_XI0/XI13/NET34_XI0/XI13/MM0_d N_WL<0>_XI0/XI13/MM0_g
+ N_BL<2>_XI0/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/MM1 N_XI0/XI13/NET33_XI0/XI13/MM1_d N_XI0/XI13/NET34_XI0/XI13/MM1_g
+ N_VSS_XI0/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/MM9 N_XI0/XI13/NET36_XI0/XI13/MM9_d N_WL<1>_XI0/XI13/MM9_g
+ N_BL<2>_XI0/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/MM6 N_XI0/XI13/NET35_XI0/XI13/MM6_d N_XI0/XI13/NET36_XI0/XI13/MM6_g
+ N_VSS_XI0/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/MM7 N_XI0/XI13/NET36_XI0/XI13/MM7_d N_XI0/XI13/NET35_XI0/XI13/MM7_g
+ N_VSS_XI0/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI13/MM8 N_XI0/XI13/NET35_XI0/XI13/MM8_d N_WL<1>_XI0/XI13/MM8_g
+ N_BLN<2>_XI0/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI13/MM5 N_XI0/XI13/NET34_XI0/XI13/MM5_d N_XI0/XI13/NET33_XI0/XI13/MM5_g
+ N_VDD_XI0/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/MM4 N_XI0/XI13/NET33_XI0/XI13/MM4_d N_XI0/XI13/NET34_XI0/XI13/MM4_g
+ N_VDD_XI0/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/MM10 N_XI0/XI13/NET35_XI0/XI13/MM10_d N_XI0/XI13/NET36_XI0/XI13/MM10_g
+ N_VDD_XI0/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI13/MM11 N_XI0/XI13/NET36_XI0/XI13/MM11_d N_XI0/XI13/NET35_XI0/XI13/MM11_g
+ N_VDD_XI0/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/MM2 N_XI0/XI14/NET34_XI0/XI14/MM2_d N_XI0/XI14/NET33_XI0/XI14/MM2_g
+ N_VSS_XI0/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/MM3 N_XI0/XI14/NET33_XI0/XI14/MM3_d N_WL<0>_XI0/XI14/MM3_g
+ N_BLN<1>_XI0/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI14/MM0 N_XI0/XI14/NET34_XI0/XI14/MM0_d N_WL<0>_XI0/XI14/MM0_g
+ N_BL<1>_XI0/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/MM1 N_XI0/XI14/NET33_XI0/XI14/MM1_d N_XI0/XI14/NET34_XI0/XI14/MM1_g
+ N_VSS_XI0/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/MM9 N_XI0/XI14/NET36_XI0/XI14/MM9_d N_WL<1>_XI0/XI14/MM9_g
+ N_BL<1>_XI0/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/MM6 N_XI0/XI14/NET35_XI0/XI14/MM6_d N_XI0/XI14/NET36_XI0/XI14/MM6_g
+ N_VSS_XI0/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/MM7 N_XI0/XI14/NET36_XI0/XI14/MM7_d N_XI0/XI14/NET35_XI0/XI14/MM7_g
+ N_VSS_XI0/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI14/MM8 N_XI0/XI14/NET35_XI0/XI14/MM8_d N_WL<1>_XI0/XI14/MM8_g
+ N_BLN<1>_XI0/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI14/MM5 N_XI0/XI14/NET34_XI0/XI14/MM5_d N_XI0/XI14/NET33_XI0/XI14/MM5_g
+ N_VDD_XI0/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/MM4 N_XI0/XI14/NET33_XI0/XI14/MM4_d N_XI0/XI14/NET34_XI0/XI14/MM4_g
+ N_VDD_XI0/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/MM10 N_XI0/XI14/NET35_XI0/XI14/MM10_d N_XI0/XI14/NET36_XI0/XI14/MM10_g
+ N_VDD_XI0/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI14/MM11 N_XI0/XI14/NET36_XI0/XI14/MM11_d N_XI0/XI14/NET35_XI0/XI14/MM11_g
+ N_VDD_XI0/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/MM2 N_XI0/XI15/NET34_XI0/XI15/MM2_d N_XI0/XI15/NET33_XI0/XI15/MM2_g
+ N_VSS_XI0/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/MM3 N_XI0/XI15/NET33_XI0/XI15/MM3_d N_WL<0>_XI0/XI15/MM3_g
+ N_BLN<0>_XI0/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI15/MM0 N_XI0/XI15/NET34_XI0/XI15/MM0_d N_WL<0>_XI0/XI15/MM0_g
+ N_BL<0>_XI0/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/MM1 N_XI0/XI15/NET33_XI0/XI15/MM1_d N_XI0/XI15/NET34_XI0/XI15/MM1_g
+ N_VSS_XI0/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/MM9 N_XI0/XI15/NET36_XI0/XI15/MM9_d N_WL<1>_XI0/XI15/MM9_g
+ N_BL<0>_XI0/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/MM6 N_XI0/XI15/NET35_XI0/XI15/MM6_d N_XI0/XI15/NET36_XI0/XI15/MM6_g
+ N_VSS_XI0/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/MM7 N_XI0/XI15/NET36_XI0/XI15/MM7_d N_XI0/XI15/NET35_XI0/XI15/MM7_g
+ N_VSS_XI0/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/XI15/MM8 N_XI0/XI15/NET35_XI0/XI15/MM8_d N_WL<1>_XI0/XI15/MM8_g
+ N_BLN<0>_XI0/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI0/XI15/MM5 N_XI0/XI15/NET34_XI0/XI15/MM5_d N_XI0/XI15/NET33_XI0/XI15/MM5_g
+ N_VDD_XI0/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/MM4 N_XI0/XI15/NET33_XI0/XI15/MM4_d N_XI0/XI15/NET34_XI0/XI15/MM4_g
+ N_VDD_XI0/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/MM10 N_XI0/XI15/NET35_XI0/XI15/MM10_d N_XI0/XI15/NET36_XI0/XI15/MM10_g
+ N_VDD_XI0/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/XI15/MM11 N_XI0/XI15/NET36_XI0/XI15/MM11_d N_XI0/XI15/NET35_XI0/XI15/MM11_g
+ N_VDD_XI0/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM2 N_XI1/XI0/NET34_XI1/XI0/MM2_d N_XI1/XI0/NET33_XI1/XI0/MM2_g
+ N_VSS_XI1/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM3 N_XI1/XI0/NET33_XI1/XI0/MM3_d N_WL<2>_XI1/XI0/MM3_g
+ N_BLN<15>_XI1/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM0 N_XI1/XI0/NET34_XI1/XI0/MM0_d N_WL<2>_XI1/XI0/MM0_g
+ N_BL<15>_XI1/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM1 N_XI1/XI0/NET33_XI1/XI0/MM1_d N_XI1/XI0/NET34_XI1/XI0/MM1_g
+ N_VSS_XI1/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM9 N_XI1/XI0/NET36_XI1/XI0/MM9_d N_WL<3>_XI1/XI0/MM9_g
+ N_BL<15>_XI1/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM6 N_XI1/XI0/NET35_XI1/XI0/MM6_d N_XI1/XI0/NET36_XI1/XI0/MM6_g
+ N_VSS_XI1/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM7 N_XI1/XI0/NET36_XI1/XI0/MM7_d N_XI1/XI0/NET35_XI1/XI0/MM7_g
+ N_VSS_XI1/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM8 N_XI1/XI0/NET35_XI1/XI0/MM8_d N_WL<3>_XI1/XI0/MM8_g
+ N_BLN<15>_XI1/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI0/MM5 N_XI1/XI0/NET34_XI1/XI0/MM5_d N_XI1/XI0/NET33_XI1/XI0/MM5_g
+ N_VDD_XI1/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM4 N_XI1/XI0/NET33_XI1/XI0/MM4_d N_XI1/XI0/NET34_XI1/XI0/MM4_g
+ N_VDD_XI1/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM10 N_XI1/XI0/NET35_XI1/XI0/MM10_d N_XI1/XI0/NET36_XI1/XI0/MM10_g
+ N_VDD_XI1/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI0/MM11 N_XI1/XI0/NET36_XI1/XI0/MM11_d N_XI1/XI0/NET35_XI1/XI0/MM11_g
+ N_VDD_XI1/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM2 N_XI1/XI1/NET34_XI1/XI1/MM2_d N_XI1/XI1/NET33_XI1/XI1/MM2_g
+ N_VSS_XI1/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM3 N_XI1/XI1/NET33_XI1/XI1/MM3_d N_WL<2>_XI1/XI1/MM3_g
+ N_BLN<14>_XI1/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM0 N_XI1/XI1/NET34_XI1/XI1/MM0_d N_WL<2>_XI1/XI1/MM0_g
+ N_BL<14>_XI1/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM1 N_XI1/XI1/NET33_XI1/XI1/MM1_d N_XI1/XI1/NET34_XI1/XI1/MM1_g
+ N_VSS_XI1/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM9 N_XI1/XI1/NET36_XI1/XI1/MM9_d N_WL<3>_XI1/XI1/MM9_g
+ N_BL<14>_XI1/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM6 N_XI1/XI1/NET35_XI1/XI1/MM6_d N_XI1/XI1/NET36_XI1/XI1/MM6_g
+ N_VSS_XI1/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM7 N_XI1/XI1/NET36_XI1/XI1/MM7_d N_XI1/XI1/NET35_XI1/XI1/MM7_g
+ N_VSS_XI1/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM8 N_XI1/XI1/NET35_XI1/XI1/MM8_d N_WL<3>_XI1/XI1/MM8_g
+ N_BLN<14>_XI1/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI1/MM5 N_XI1/XI1/NET34_XI1/XI1/MM5_d N_XI1/XI1/NET33_XI1/XI1/MM5_g
+ N_VDD_XI1/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM4 N_XI1/XI1/NET33_XI1/XI1/MM4_d N_XI1/XI1/NET34_XI1/XI1/MM4_g
+ N_VDD_XI1/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM10 N_XI1/XI1/NET35_XI1/XI1/MM10_d N_XI1/XI1/NET36_XI1/XI1/MM10_g
+ N_VDD_XI1/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI1/MM11 N_XI1/XI1/NET36_XI1/XI1/MM11_d N_XI1/XI1/NET35_XI1/XI1/MM11_g
+ N_VDD_XI1/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM2 N_XI1/XI2/NET34_XI1/XI2/MM2_d N_XI1/XI2/NET33_XI1/XI2/MM2_g
+ N_VSS_XI1/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM3 N_XI1/XI2/NET33_XI1/XI2/MM3_d N_WL<2>_XI1/XI2/MM3_g
+ N_BLN<13>_XI1/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM0 N_XI1/XI2/NET34_XI1/XI2/MM0_d N_WL<2>_XI1/XI2/MM0_g
+ N_BL<13>_XI1/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM1 N_XI1/XI2/NET33_XI1/XI2/MM1_d N_XI1/XI2/NET34_XI1/XI2/MM1_g
+ N_VSS_XI1/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM9 N_XI1/XI2/NET36_XI1/XI2/MM9_d N_WL<3>_XI1/XI2/MM9_g
+ N_BL<13>_XI1/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM6 N_XI1/XI2/NET35_XI1/XI2/MM6_d N_XI1/XI2/NET36_XI1/XI2/MM6_g
+ N_VSS_XI1/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM7 N_XI1/XI2/NET36_XI1/XI2/MM7_d N_XI1/XI2/NET35_XI1/XI2/MM7_g
+ N_VSS_XI1/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM8 N_XI1/XI2/NET35_XI1/XI2/MM8_d N_WL<3>_XI1/XI2/MM8_g
+ N_BLN<13>_XI1/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI2/MM5 N_XI1/XI2/NET34_XI1/XI2/MM5_d N_XI1/XI2/NET33_XI1/XI2/MM5_g
+ N_VDD_XI1/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM4 N_XI1/XI2/NET33_XI1/XI2/MM4_d N_XI1/XI2/NET34_XI1/XI2/MM4_g
+ N_VDD_XI1/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM10 N_XI1/XI2/NET35_XI1/XI2/MM10_d N_XI1/XI2/NET36_XI1/XI2/MM10_g
+ N_VDD_XI1/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI2/MM11 N_XI1/XI2/NET36_XI1/XI2/MM11_d N_XI1/XI2/NET35_XI1/XI2/MM11_g
+ N_VDD_XI1/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM2 N_XI1/XI3/NET34_XI1/XI3/MM2_d N_XI1/XI3/NET33_XI1/XI3/MM2_g
+ N_VSS_XI1/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM3 N_XI1/XI3/NET33_XI1/XI3/MM3_d N_WL<2>_XI1/XI3/MM3_g
+ N_BLN<12>_XI1/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM0 N_XI1/XI3/NET34_XI1/XI3/MM0_d N_WL<2>_XI1/XI3/MM0_g
+ N_BL<12>_XI1/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM1 N_XI1/XI3/NET33_XI1/XI3/MM1_d N_XI1/XI3/NET34_XI1/XI3/MM1_g
+ N_VSS_XI1/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM9 N_XI1/XI3/NET36_XI1/XI3/MM9_d N_WL<3>_XI1/XI3/MM9_g
+ N_BL<12>_XI1/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM6 N_XI1/XI3/NET35_XI1/XI3/MM6_d N_XI1/XI3/NET36_XI1/XI3/MM6_g
+ N_VSS_XI1/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM7 N_XI1/XI3/NET36_XI1/XI3/MM7_d N_XI1/XI3/NET35_XI1/XI3/MM7_g
+ N_VSS_XI1/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM8 N_XI1/XI3/NET35_XI1/XI3/MM8_d N_WL<3>_XI1/XI3/MM8_g
+ N_BLN<12>_XI1/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI3/MM5 N_XI1/XI3/NET34_XI1/XI3/MM5_d N_XI1/XI3/NET33_XI1/XI3/MM5_g
+ N_VDD_XI1/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM4 N_XI1/XI3/NET33_XI1/XI3/MM4_d N_XI1/XI3/NET34_XI1/XI3/MM4_g
+ N_VDD_XI1/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM10 N_XI1/XI3/NET35_XI1/XI3/MM10_d N_XI1/XI3/NET36_XI1/XI3/MM10_g
+ N_VDD_XI1/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI3/MM11 N_XI1/XI3/NET36_XI1/XI3/MM11_d N_XI1/XI3/NET35_XI1/XI3/MM11_g
+ N_VDD_XI1/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM2 N_XI1/XI4/NET34_XI1/XI4/MM2_d N_XI1/XI4/NET33_XI1/XI4/MM2_g
+ N_VSS_XI1/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM3 N_XI1/XI4/NET33_XI1/XI4/MM3_d N_WL<2>_XI1/XI4/MM3_g
+ N_BLN<11>_XI1/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM0 N_XI1/XI4/NET34_XI1/XI4/MM0_d N_WL<2>_XI1/XI4/MM0_g
+ N_BL<11>_XI1/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM1 N_XI1/XI4/NET33_XI1/XI4/MM1_d N_XI1/XI4/NET34_XI1/XI4/MM1_g
+ N_VSS_XI1/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM9 N_XI1/XI4/NET36_XI1/XI4/MM9_d N_WL<3>_XI1/XI4/MM9_g
+ N_BL<11>_XI1/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM6 N_XI1/XI4/NET35_XI1/XI4/MM6_d N_XI1/XI4/NET36_XI1/XI4/MM6_g
+ N_VSS_XI1/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM7 N_XI1/XI4/NET36_XI1/XI4/MM7_d N_XI1/XI4/NET35_XI1/XI4/MM7_g
+ N_VSS_XI1/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM8 N_XI1/XI4/NET35_XI1/XI4/MM8_d N_WL<3>_XI1/XI4/MM8_g
+ N_BLN<11>_XI1/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI4/MM5 N_XI1/XI4/NET34_XI1/XI4/MM5_d N_XI1/XI4/NET33_XI1/XI4/MM5_g
+ N_VDD_XI1/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM4 N_XI1/XI4/NET33_XI1/XI4/MM4_d N_XI1/XI4/NET34_XI1/XI4/MM4_g
+ N_VDD_XI1/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM10 N_XI1/XI4/NET35_XI1/XI4/MM10_d N_XI1/XI4/NET36_XI1/XI4/MM10_g
+ N_VDD_XI1/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI4/MM11 N_XI1/XI4/NET36_XI1/XI4/MM11_d N_XI1/XI4/NET35_XI1/XI4/MM11_g
+ N_VDD_XI1/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM2 N_XI1/XI5/NET34_XI1/XI5/MM2_d N_XI1/XI5/NET33_XI1/XI5/MM2_g
+ N_VSS_XI1/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM3 N_XI1/XI5/NET33_XI1/XI5/MM3_d N_WL<2>_XI1/XI5/MM3_g
+ N_BLN<10>_XI1/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM0 N_XI1/XI5/NET34_XI1/XI5/MM0_d N_WL<2>_XI1/XI5/MM0_g
+ N_BL<10>_XI1/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM1 N_XI1/XI5/NET33_XI1/XI5/MM1_d N_XI1/XI5/NET34_XI1/XI5/MM1_g
+ N_VSS_XI1/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM9 N_XI1/XI5/NET36_XI1/XI5/MM9_d N_WL<3>_XI1/XI5/MM9_g
+ N_BL<10>_XI1/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM6 N_XI1/XI5/NET35_XI1/XI5/MM6_d N_XI1/XI5/NET36_XI1/XI5/MM6_g
+ N_VSS_XI1/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM7 N_XI1/XI5/NET36_XI1/XI5/MM7_d N_XI1/XI5/NET35_XI1/XI5/MM7_g
+ N_VSS_XI1/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM8 N_XI1/XI5/NET35_XI1/XI5/MM8_d N_WL<3>_XI1/XI5/MM8_g
+ N_BLN<10>_XI1/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI5/MM5 N_XI1/XI5/NET34_XI1/XI5/MM5_d N_XI1/XI5/NET33_XI1/XI5/MM5_g
+ N_VDD_XI1/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM4 N_XI1/XI5/NET33_XI1/XI5/MM4_d N_XI1/XI5/NET34_XI1/XI5/MM4_g
+ N_VDD_XI1/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM10 N_XI1/XI5/NET35_XI1/XI5/MM10_d N_XI1/XI5/NET36_XI1/XI5/MM10_g
+ N_VDD_XI1/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI5/MM11 N_XI1/XI5/NET36_XI1/XI5/MM11_d N_XI1/XI5/NET35_XI1/XI5/MM11_g
+ N_VDD_XI1/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM2 N_XI1/XI6/NET34_XI1/XI6/MM2_d N_XI1/XI6/NET33_XI1/XI6/MM2_g
+ N_VSS_XI1/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM3 N_XI1/XI6/NET33_XI1/XI6/MM3_d N_WL<2>_XI1/XI6/MM3_g
+ N_BLN<9>_XI1/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM0 N_XI1/XI6/NET34_XI1/XI6/MM0_d N_WL<2>_XI1/XI6/MM0_g
+ N_BL<9>_XI1/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM1 N_XI1/XI6/NET33_XI1/XI6/MM1_d N_XI1/XI6/NET34_XI1/XI6/MM1_g
+ N_VSS_XI1/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM9 N_XI1/XI6/NET36_XI1/XI6/MM9_d N_WL<3>_XI1/XI6/MM9_g
+ N_BL<9>_XI1/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM6 N_XI1/XI6/NET35_XI1/XI6/MM6_d N_XI1/XI6/NET36_XI1/XI6/MM6_g
+ N_VSS_XI1/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM7 N_XI1/XI6/NET36_XI1/XI6/MM7_d N_XI1/XI6/NET35_XI1/XI6/MM7_g
+ N_VSS_XI1/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM8 N_XI1/XI6/NET35_XI1/XI6/MM8_d N_WL<3>_XI1/XI6/MM8_g
+ N_BLN<9>_XI1/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI6/MM5 N_XI1/XI6/NET34_XI1/XI6/MM5_d N_XI1/XI6/NET33_XI1/XI6/MM5_g
+ N_VDD_XI1/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM4 N_XI1/XI6/NET33_XI1/XI6/MM4_d N_XI1/XI6/NET34_XI1/XI6/MM4_g
+ N_VDD_XI1/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM10 N_XI1/XI6/NET35_XI1/XI6/MM10_d N_XI1/XI6/NET36_XI1/XI6/MM10_g
+ N_VDD_XI1/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI6/MM11 N_XI1/XI6/NET36_XI1/XI6/MM11_d N_XI1/XI6/NET35_XI1/XI6/MM11_g
+ N_VDD_XI1/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM2 N_XI1/XI7/NET34_XI1/XI7/MM2_d N_XI1/XI7/NET33_XI1/XI7/MM2_g
+ N_VSS_XI1/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM3 N_XI1/XI7/NET33_XI1/XI7/MM3_d N_WL<2>_XI1/XI7/MM3_g
+ N_BLN<8>_XI1/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM0 N_XI1/XI7/NET34_XI1/XI7/MM0_d N_WL<2>_XI1/XI7/MM0_g
+ N_BL<8>_XI1/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM1 N_XI1/XI7/NET33_XI1/XI7/MM1_d N_XI1/XI7/NET34_XI1/XI7/MM1_g
+ N_VSS_XI1/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM9 N_XI1/XI7/NET36_XI1/XI7/MM9_d N_WL<3>_XI1/XI7/MM9_g
+ N_BL<8>_XI1/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM6 N_XI1/XI7/NET35_XI1/XI7/MM6_d N_XI1/XI7/NET36_XI1/XI7/MM6_g
+ N_VSS_XI1/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM7 N_XI1/XI7/NET36_XI1/XI7/MM7_d N_XI1/XI7/NET35_XI1/XI7/MM7_g
+ N_VSS_XI1/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM8 N_XI1/XI7/NET35_XI1/XI7/MM8_d N_WL<3>_XI1/XI7/MM8_g
+ N_BLN<8>_XI1/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI7/MM5 N_XI1/XI7/NET34_XI1/XI7/MM5_d N_XI1/XI7/NET33_XI1/XI7/MM5_g
+ N_VDD_XI1/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM4 N_XI1/XI7/NET33_XI1/XI7/MM4_d N_XI1/XI7/NET34_XI1/XI7/MM4_g
+ N_VDD_XI1/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM10 N_XI1/XI7/NET35_XI1/XI7/MM10_d N_XI1/XI7/NET36_XI1/XI7/MM10_g
+ N_VDD_XI1/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI7/MM11 N_XI1/XI7/NET36_XI1/XI7/MM11_d N_XI1/XI7/NET35_XI1/XI7/MM11_g
+ N_VDD_XI1/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM2 N_XI1/XI8/NET34_XI1/XI8/MM2_d N_XI1/XI8/NET33_XI1/XI8/MM2_g
+ N_VSS_XI1/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM3 N_XI1/XI8/NET33_XI1/XI8/MM3_d N_WL<2>_XI1/XI8/MM3_g
+ N_BLN<7>_XI1/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM0 N_XI1/XI8/NET34_XI1/XI8/MM0_d N_WL<2>_XI1/XI8/MM0_g
+ N_BL<7>_XI1/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM1 N_XI1/XI8/NET33_XI1/XI8/MM1_d N_XI1/XI8/NET34_XI1/XI8/MM1_g
+ N_VSS_XI1/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM9 N_XI1/XI8/NET36_XI1/XI8/MM9_d N_WL<3>_XI1/XI8/MM9_g
+ N_BL<7>_XI1/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM6 N_XI1/XI8/NET35_XI1/XI8/MM6_d N_XI1/XI8/NET36_XI1/XI8/MM6_g
+ N_VSS_XI1/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM7 N_XI1/XI8/NET36_XI1/XI8/MM7_d N_XI1/XI8/NET35_XI1/XI8/MM7_g
+ N_VSS_XI1/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM8 N_XI1/XI8/NET35_XI1/XI8/MM8_d N_WL<3>_XI1/XI8/MM8_g
+ N_BLN<7>_XI1/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI8/MM5 N_XI1/XI8/NET34_XI1/XI8/MM5_d N_XI1/XI8/NET33_XI1/XI8/MM5_g
+ N_VDD_XI1/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM4 N_XI1/XI8/NET33_XI1/XI8/MM4_d N_XI1/XI8/NET34_XI1/XI8/MM4_g
+ N_VDD_XI1/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM10 N_XI1/XI8/NET35_XI1/XI8/MM10_d N_XI1/XI8/NET36_XI1/XI8/MM10_g
+ N_VDD_XI1/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI8/MM11 N_XI1/XI8/NET36_XI1/XI8/MM11_d N_XI1/XI8/NET35_XI1/XI8/MM11_g
+ N_VDD_XI1/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM2 N_XI1/XI9/NET34_XI1/XI9/MM2_d N_XI1/XI9/NET33_XI1/XI9/MM2_g
+ N_VSS_XI1/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM3 N_XI1/XI9/NET33_XI1/XI9/MM3_d N_WL<2>_XI1/XI9/MM3_g
+ N_BLN<6>_XI1/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM0 N_XI1/XI9/NET34_XI1/XI9/MM0_d N_WL<2>_XI1/XI9/MM0_g
+ N_BL<6>_XI1/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM1 N_XI1/XI9/NET33_XI1/XI9/MM1_d N_XI1/XI9/NET34_XI1/XI9/MM1_g
+ N_VSS_XI1/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM9 N_XI1/XI9/NET36_XI1/XI9/MM9_d N_WL<3>_XI1/XI9/MM9_g
+ N_BL<6>_XI1/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM6 N_XI1/XI9/NET35_XI1/XI9/MM6_d N_XI1/XI9/NET36_XI1/XI9/MM6_g
+ N_VSS_XI1/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM7 N_XI1/XI9/NET36_XI1/XI9/MM7_d N_XI1/XI9/NET35_XI1/XI9/MM7_g
+ N_VSS_XI1/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM8 N_XI1/XI9/NET35_XI1/XI9/MM8_d N_WL<3>_XI1/XI9/MM8_g
+ N_BLN<6>_XI1/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI9/MM5 N_XI1/XI9/NET34_XI1/XI9/MM5_d N_XI1/XI9/NET33_XI1/XI9/MM5_g
+ N_VDD_XI1/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM4 N_XI1/XI9/NET33_XI1/XI9/MM4_d N_XI1/XI9/NET34_XI1/XI9/MM4_g
+ N_VDD_XI1/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM10 N_XI1/XI9/NET35_XI1/XI9/MM10_d N_XI1/XI9/NET36_XI1/XI9/MM10_g
+ N_VDD_XI1/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI9/MM11 N_XI1/XI9/NET36_XI1/XI9/MM11_d N_XI1/XI9/NET35_XI1/XI9/MM11_g
+ N_VDD_XI1/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM2 N_XI1/XI10/NET34_XI1/XI10/MM2_d N_XI1/XI10/NET33_XI1/XI10/MM2_g
+ N_VSS_XI1/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI10/MM3 N_XI1/XI10/NET33_XI1/XI10/MM3_d N_WL<2>_XI1/XI10/MM3_g
+ N_BLN<5>_XI1/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI10/MM0 N_XI1/XI10/NET34_XI1/XI10/MM0_d N_WL<2>_XI1/XI10/MM0_g
+ N_BL<5>_XI1/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI10/MM1 N_XI1/XI10/NET33_XI1/XI10/MM1_d N_XI1/XI10/NET34_XI1/XI10/MM1_g
+ N_VSS_XI1/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI10/MM9 N_XI1/XI10/NET36_XI1/XI10/MM9_d N_WL<3>_XI1/XI10/MM9_g
+ N_BL<5>_XI1/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI10/MM6 N_XI1/XI10/NET35_XI1/XI10/MM6_d N_XI1/XI10/NET36_XI1/XI10/MM6_g
+ N_VSS_XI1/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI10/MM7 N_XI1/XI10/NET36_XI1/XI10/MM7_d N_XI1/XI10/NET35_XI1/XI10/MM7_g
+ N_VSS_XI1/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI10/MM8 N_XI1/XI10/NET35_XI1/XI10/MM8_d N_WL<3>_XI1/XI10/MM8_g
+ N_BLN<5>_XI1/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI10/MM5 N_XI1/XI10/NET34_XI1/XI10/MM5_d N_XI1/XI10/NET33_XI1/XI10/MM5_g
+ N_VDD_XI1/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM4 N_XI1/XI10/NET33_XI1/XI10/MM4_d N_XI1/XI10/NET34_XI1/XI10/MM4_g
+ N_VDD_XI1/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM10 N_XI1/XI10/NET35_XI1/XI10/MM10_d N_XI1/XI10/NET36_XI1/XI10/MM10_g
+ N_VDD_XI1/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI10/MM11 N_XI1/XI10/NET36_XI1/XI10/MM11_d N_XI1/XI10/NET35_XI1/XI10/MM11_g
+ N_VDD_XI1/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM2 N_XI1/XI11/NET34_XI1/XI11/MM2_d N_XI1/XI11/NET33_XI1/XI11/MM2_g
+ N_VSS_XI1/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI11/MM3 N_XI1/XI11/NET33_XI1/XI11/MM3_d N_WL<2>_XI1/XI11/MM3_g
+ N_BLN<4>_XI1/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI11/MM0 N_XI1/XI11/NET34_XI1/XI11/MM0_d N_WL<2>_XI1/XI11/MM0_g
+ N_BL<4>_XI1/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI11/MM1 N_XI1/XI11/NET33_XI1/XI11/MM1_d N_XI1/XI11/NET34_XI1/XI11/MM1_g
+ N_VSS_XI1/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI11/MM9 N_XI1/XI11/NET36_XI1/XI11/MM9_d N_WL<3>_XI1/XI11/MM9_g
+ N_BL<4>_XI1/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI11/MM6 N_XI1/XI11/NET35_XI1/XI11/MM6_d N_XI1/XI11/NET36_XI1/XI11/MM6_g
+ N_VSS_XI1/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI11/MM7 N_XI1/XI11/NET36_XI1/XI11/MM7_d N_XI1/XI11/NET35_XI1/XI11/MM7_g
+ N_VSS_XI1/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI11/MM8 N_XI1/XI11/NET35_XI1/XI11/MM8_d N_WL<3>_XI1/XI11/MM8_g
+ N_BLN<4>_XI1/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI11/MM5 N_XI1/XI11/NET34_XI1/XI11/MM5_d N_XI1/XI11/NET33_XI1/XI11/MM5_g
+ N_VDD_XI1/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM4 N_XI1/XI11/NET33_XI1/XI11/MM4_d N_XI1/XI11/NET34_XI1/XI11/MM4_g
+ N_VDD_XI1/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM10 N_XI1/XI11/NET35_XI1/XI11/MM10_d N_XI1/XI11/NET36_XI1/XI11/MM10_g
+ N_VDD_XI1/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI11/MM11 N_XI1/XI11/NET36_XI1/XI11/MM11_d N_XI1/XI11/NET35_XI1/XI11/MM11_g
+ N_VDD_XI1/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM2 N_XI1/XI12/NET34_XI1/XI12/MM2_d N_XI1/XI12/NET33_XI1/XI12/MM2_g
+ N_VSS_XI1/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI12/MM3 N_XI1/XI12/NET33_XI1/XI12/MM3_d N_WL<2>_XI1/XI12/MM3_g
+ N_BLN<3>_XI1/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI12/MM0 N_XI1/XI12/NET34_XI1/XI12/MM0_d N_WL<2>_XI1/XI12/MM0_g
+ N_BL<3>_XI1/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI12/MM1 N_XI1/XI12/NET33_XI1/XI12/MM1_d N_XI1/XI12/NET34_XI1/XI12/MM1_g
+ N_VSS_XI1/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI12/MM9 N_XI1/XI12/NET36_XI1/XI12/MM9_d N_WL<3>_XI1/XI12/MM9_g
+ N_BL<3>_XI1/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI12/MM6 N_XI1/XI12/NET35_XI1/XI12/MM6_d N_XI1/XI12/NET36_XI1/XI12/MM6_g
+ N_VSS_XI1/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI12/MM7 N_XI1/XI12/NET36_XI1/XI12/MM7_d N_XI1/XI12/NET35_XI1/XI12/MM7_g
+ N_VSS_XI1/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI12/MM8 N_XI1/XI12/NET35_XI1/XI12/MM8_d N_WL<3>_XI1/XI12/MM8_g
+ N_BLN<3>_XI1/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI12/MM5 N_XI1/XI12/NET34_XI1/XI12/MM5_d N_XI1/XI12/NET33_XI1/XI12/MM5_g
+ N_VDD_XI1/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM4 N_XI1/XI12/NET33_XI1/XI12/MM4_d N_XI1/XI12/NET34_XI1/XI12/MM4_g
+ N_VDD_XI1/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM10 N_XI1/XI12/NET35_XI1/XI12/MM10_d N_XI1/XI12/NET36_XI1/XI12/MM10_g
+ N_VDD_XI1/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI12/MM11 N_XI1/XI12/NET36_XI1/XI12/MM11_d N_XI1/XI12/NET35_XI1/XI12/MM11_g
+ N_VDD_XI1/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM2 N_XI1/XI13/NET34_XI1/XI13/MM2_d N_XI1/XI13/NET33_XI1/XI13/MM2_g
+ N_VSS_XI1/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI13/MM3 N_XI1/XI13/NET33_XI1/XI13/MM3_d N_WL<2>_XI1/XI13/MM3_g
+ N_BLN<2>_XI1/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI13/MM0 N_XI1/XI13/NET34_XI1/XI13/MM0_d N_WL<2>_XI1/XI13/MM0_g
+ N_BL<2>_XI1/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI13/MM1 N_XI1/XI13/NET33_XI1/XI13/MM1_d N_XI1/XI13/NET34_XI1/XI13/MM1_g
+ N_VSS_XI1/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI13/MM9 N_XI1/XI13/NET36_XI1/XI13/MM9_d N_WL<3>_XI1/XI13/MM9_g
+ N_BL<2>_XI1/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI13/MM6 N_XI1/XI13/NET35_XI1/XI13/MM6_d N_XI1/XI13/NET36_XI1/XI13/MM6_g
+ N_VSS_XI1/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI13/MM7 N_XI1/XI13/NET36_XI1/XI13/MM7_d N_XI1/XI13/NET35_XI1/XI13/MM7_g
+ N_VSS_XI1/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI13/MM8 N_XI1/XI13/NET35_XI1/XI13/MM8_d N_WL<3>_XI1/XI13/MM8_g
+ N_BLN<2>_XI1/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI13/MM5 N_XI1/XI13/NET34_XI1/XI13/MM5_d N_XI1/XI13/NET33_XI1/XI13/MM5_g
+ N_VDD_XI1/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM4 N_XI1/XI13/NET33_XI1/XI13/MM4_d N_XI1/XI13/NET34_XI1/XI13/MM4_g
+ N_VDD_XI1/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM10 N_XI1/XI13/NET35_XI1/XI13/MM10_d N_XI1/XI13/NET36_XI1/XI13/MM10_g
+ N_VDD_XI1/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI13/MM11 N_XI1/XI13/NET36_XI1/XI13/MM11_d N_XI1/XI13/NET35_XI1/XI13/MM11_g
+ N_VDD_XI1/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM2 N_XI1/XI14/NET34_XI1/XI14/MM2_d N_XI1/XI14/NET33_XI1/XI14/MM2_g
+ N_VSS_XI1/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI14/MM3 N_XI1/XI14/NET33_XI1/XI14/MM3_d N_WL<2>_XI1/XI14/MM3_g
+ N_BLN<1>_XI1/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI14/MM0 N_XI1/XI14/NET34_XI1/XI14/MM0_d N_WL<2>_XI1/XI14/MM0_g
+ N_BL<1>_XI1/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI14/MM1 N_XI1/XI14/NET33_XI1/XI14/MM1_d N_XI1/XI14/NET34_XI1/XI14/MM1_g
+ N_VSS_XI1/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI14/MM9 N_XI1/XI14/NET36_XI1/XI14/MM9_d N_WL<3>_XI1/XI14/MM9_g
+ N_BL<1>_XI1/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI14/MM6 N_XI1/XI14/NET35_XI1/XI14/MM6_d N_XI1/XI14/NET36_XI1/XI14/MM6_g
+ N_VSS_XI1/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI14/MM7 N_XI1/XI14/NET36_XI1/XI14/MM7_d N_XI1/XI14/NET35_XI1/XI14/MM7_g
+ N_VSS_XI1/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI14/MM8 N_XI1/XI14/NET35_XI1/XI14/MM8_d N_WL<3>_XI1/XI14/MM8_g
+ N_BLN<1>_XI1/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI14/MM5 N_XI1/XI14/NET34_XI1/XI14/MM5_d N_XI1/XI14/NET33_XI1/XI14/MM5_g
+ N_VDD_XI1/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM4 N_XI1/XI14/NET33_XI1/XI14/MM4_d N_XI1/XI14/NET34_XI1/XI14/MM4_g
+ N_VDD_XI1/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM10 N_XI1/XI14/NET35_XI1/XI14/MM10_d N_XI1/XI14/NET36_XI1/XI14/MM10_g
+ N_VDD_XI1/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI14/MM11 N_XI1/XI14/NET36_XI1/XI14/MM11_d N_XI1/XI14/NET35_XI1/XI14/MM11_g
+ N_VDD_XI1/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM2 N_XI1/XI15/NET34_XI1/XI15/MM2_d N_XI1/XI15/NET33_XI1/XI15/MM2_g
+ N_VSS_XI1/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI15/MM3 N_XI1/XI15/NET33_XI1/XI15/MM3_d N_WL<2>_XI1/XI15/MM3_g
+ N_BLN<0>_XI1/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI15/MM0 N_XI1/XI15/NET34_XI1/XI15/MM0_d N_WL<2>_XI1/XI15/MM0_g
+ N_BL<0>_XI1/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI15/MM1 N_XI1/XI15/NET33_XI1/XI15/MM1_d N_XI1/XI15/NET34_XI1/XI15/MM1_g
+ N_VSS_XI1/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI15/MM9 N_XI1/XI15/NET36_XI1/XI15/MM9_d N_WL<3>_XI1/XI15/MM9_g
+ N_BL<0>_XI1/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI15/MM6 N_XI1/XI15/NET35_XI1/XI15/MM6_d N_XI1/XI15/NET36_XI1/XI15/MM6_g
+ N_VSS_XI1/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI15/MM7 N_XI1/XI15/NET36_XI1/XI15/MM7_d N_XI1/XI15/NET35_XI1/XI15/MM7_g
+ N_VSS_XI1/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/XI15/MM8 N_XI1/XI15/NET35_XI1/XI15/MM8_d N_WL<3>_XI1/XI15/MM8_g
+ N_BLN<0>_XI1/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI1/XI15/MM5 N_XI1/XI15/NET34_XI1/XI15/MM5_d N_XI1/XI15/NET33_XI1/XI15/MM5_g
+ N_VDD_XI1/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM4 N_XI1/XI15/NET33_XI1/XI15/MM4_d N_XI1/XI15/NET34_XI1/XI15/MM4_g
+ N_VDD_XI1/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM10 N_XI1/XI15/NET35_XI1/XI15/MM10_d N_XI1/XI15/NET36_XI1/XI15/MM10_g
+ N_VDD_XI1/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/XI15/MM11 N_XI1/XI15/NET36_XI1/XI15/MM11_d N_XI1/XI15/NET35_XI1/XI15/MM11_g
+ N_VDD_XI1/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI0/MM2 N_XI4/XI0/NET34_XI4/XI0/MM2_d N_XI4/XI0/NET33_XI4/XI0/MM2_g
+ N_VSS_XI4/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM3 N_XI4/XI0/NET33_XI4/XI0/MM3_d N_WL<4>_XI4/XI0/MM3_g
+ N_BLN<15>_XI4/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM0 N_XI4/XI0/NET34_XI4/XI0/MM0_d N_WL<4>_XI4/XI0/MM0_g
+ N_BL<15>_XI4/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM1 N_XI4/XI0/NET33_XI4/XI0/MM1_d N_XI4/XI0/NET34_XI4/XI0/MM1_g
+ N_VSS_XI4/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM9 N_XI4/XI0/NET36_XI4/XI0/MM9_d N_WL<5>_XI4/XI0/MM9_g
+ N_BL<15>_XI4/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM6 N_XI4/XI0/NET35_XI4/XI0/MM6_d N_XI4/XI0/NET36_XI4/XI0/MM6_g
+ N_VSS_XI4/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM7 N_XI4/XI0/NET36_XI4/XI0/MM7_d N_XI4/XI0/NET35_XI4/XI0/MM7_g
+ N_VSS_XI4/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM8 N_XI4/XI0/NET35_XI4/XI0/MM8_d N_WL<5>_XI4/XI0/MM8_g
+ N_BLN<15>_XI4/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI0/MM5 N_XI4/XI0/NET34_XI4/XI0/MM5_d N_XI4/XI0/NET33_XI4/XI0/MM5_g
+ N_VDD_XI4/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI0/MM4 N_XI4/XI0/NET33_XI4/XI0/MM4_d N_XI4/XI0/NET34_XI4/XI0/MM4_g
+ N_VDD_XI4/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI0/MM10 N_XI4/XI0/NET35_XI4/XI0/MM10_d N_XI4/XI0/NET36_XI4/XI0/MM10_g
+ N_VDD_XI4/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI0/MM11 N_XI4/XI0/NET36_XI4/XI0/MM11_d N_XI4/XI0/NET35_XI4/XI0/MM11_g
+ N_VDD_XI4/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI1/MM2 N_XI4/XI1/NET34_XI4/XI1/MM2_d N_XI4/XI1/NET33_XI4/XI1/MM2_g
+ N_VSS_XI4/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM3 N_XI4/XI1/NET33_XI4/XI1/MM3_d N_WL<4>_XI4/XI1/MM3_g
+ N_BLN<14>_XI4/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM0 N_XI4/XI1/NET34_XI4/XI1/MM0_d N_WL<4>_XI4/XI1/MM0_g
+ N_BL<14>_XI4/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM1 N_XI4/XI1/NET33_XI4/XI1/MM1_d N_XI4/XI1/NET34_XI4/XI1/MM1_g
+ N_VSS_XI4/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM9 N_XI4/XI1/NET36_XI4/XI1/MM9_d N_WL<5>_XI4/XI1/MM9_g
+ N_BL<14>_XI4/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM6 N_XI4/XI1/NET35_XI4/XI1/MM6_d N_XI4/XI1/NET36_XI4/XI1/MM6_g
+ N_VSS_XI4/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM7 N_XI4/XI1/NET36_XI4/XI1/MM7_d N_XI4/XI1/NET35_XI4/XI1/MM7_g
+ N_VSS_XI4/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM8 N_XI4/XI1/NET35_XI4/XI1/MM8_d N_WL<5>_XI4/XI1/MM8_g
+ N_BLN<14>_XI4/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI1/MM5 N_XI4/XI1/NET34_XI4/XI1/MM5_d N_XI4/XI1/NET33_XI4/XI1/MM5_g
+ N_VDD_XI4/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI1/MM4 N_XI4/XI1/NET33_XI4/XI1/MM4_d N_XI4/XI1/NET34_XI4/XI1/MM4_g
+ N_VDD_XI4/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI1/MM10 N_XI4/XI1/NET35_XI4/XI1/MM10_d N_XI4/XI1/NET36_XI4/XI1/MM10_g
+ N_VDD_XI4/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI1/MM11 N_XI4/XI1/NET36_XI4/XI1/MM11_d N_XI4/XI1/NET35_XI4/XI1/MM11_g
+ N_VDD_XI4/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI2/MM2 N_XI4/XI2/NET34_XI4/XI2/MM2_d N_XI4/XI2/NET33_XI4/XI2/MM2_g
+ N_VSS_XI4/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM3 N_XI4/XI2/NET33_XI4/XI2/MM3_d N_WL<4>_XI4/XI2/MM3_g
+ N_BLN<13>_XI4/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM0 N_XI4/XI2/NET34_XI4/XI2/MM0_d N_WL<4>_XI4/XI2/MM0_g
+ N_BL<13>_XI4/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM1 N_XI4/XI2/NET33_XI4/XI2/MM1_d N_XI4/XI2/NET34_XI4/XI2/MM1_g
+ N_VSS_XI4/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM9 N_XI4/XI2/NET36_XI4/XI2/MM9_d N_WL<5>_XI4/XI2/MM9_g
+ N_BL<13>_XI4/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM6 N_XI4/XI2/NET35_XI4/XI2/MM6_d N_XI4/XI2/NET36_XI4/XI2/MM6_g
+ N_VSS_XI4/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM7 N_XI4/XI2/NET36_XI4/XI2/MM7_d N_XI4/XI2/NET35_XI4/XI2/MM7_g
+ N_VSS_XI4/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM8 N_XI4/XI2/NET35_XI4/XI2/MM8_d N_WL<5>_XI4/XI2/MM8_g
+ N_BLN<13>_XI4/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI2/MM5 N_XI4/XI2/NET34_XI4/XI2/MM5_d N_XI4/XI2/NET33_XI4/XI2/MM5_g
+ N_VDD_XI4/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI2/MM4 N_XI4/XI2/NET33_XI4/XI2/MM4_d N_XI4/XI2/NET34_XI4/XI2/MM4_g
+ N_VDD_XI4/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI2/MM10 N_XI4/XI2/NET35_XI4/XI2/MM10_d N_XI4/XI2/NET36_XI4/XI2/MM10_g
+ N_VDD_XI4/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI2/MM11 N_XI4/XI2/NET36_XI4/XI2/MM11_d N_XI4/XI2/NET35_XI4/XI2/MM11_g
+ N_VDD_XI4/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI3/MM2 N_XI4/XI3/NET34_XI4/XI3/MM2_d N_XI4/XI3/NET33_XI4/XI3/MM2_g
+ N_VSS_XI4/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM3 N_XI4/XI3/NET33_XI4/XI3/MM3_d N_WL<4>_XI4/XI3/MM3_g
+ N_BLN<12>_XI4/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM0 N_XI4/XI3/NET34_XI4/XI3/MM0_d N_WL<4>_XI4/XI3/MM0_g
+ N_BL<12>_XI4/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM1 N_XI4/XI3/NET33_XI4/XI3/MM1_d N_XI4/XI3/NET34_XI4/XI3/MM1_g
+ N_VSS_XI4/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM9 N_XI4/XI3/NET36_XI4/XI3/MM9_d N_WL<5>_XI4/XI3/MM9_g
+ N_BL<12>_XI4/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM6 N_XI4/XI3/NET35_XI4/XI3/MM6_d N_XI4/XI3/NET36_XI4/XI3/MM6_g
+ N_VSS_XI4/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM7 N_XI4/XI3/NET36_XI4/XI3/MM7_d N_XI4/XI3/NET35_XI4/XI3/MM7_g
+ N_VSS_XI4/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM8 N_XI4/XI3/NET35_XI4/XI3/MM8_d N_WL<5>_XI4/XI3/MM8_g
+ N_BLN<12>_XI4/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI3/MM5 N_XI4/XI3/NET34_XI4/XI3/MM5_d N_XI4/XI3/NET33_XI4/XI3/MM5_g
+ N_VDD_XI4/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI3/MM4 N_XI4/XI3/NET33_XI4/XI3/MM4_d N_XI4/XI3/NET34_XI4/XI3/MM4_g
+ N_VDD_XI4/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI3/MM10 N_XI4/XI3/NET35_XI4/XI3/MM10_d N_XI4/XI3/NET36_XI4/XI3/MM10_g
+ N_VDD_XI4/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI3/MM11 N_XI4/XI3/NET36_XI4/XI3/MM11_d N_XI4/XI3/NET35_XI4/XI3/MM11_g
+ N_VDD_XI4/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI4/MM2 N_XI4/XI4/NET34_XI4/XI4/MM2_d N_XI4/XI4/NET33_XI4/XI4/MM2_g
+ N_VSS_XI4/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM3 N_XI4/XI4/NET33_XI4/XI4/MM3_d N_WL<4>_XI4/XI4/MM3_g
+ N_BLN<11>_XI4/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM0 N_XI4/XI4/NET34_XI4/XI4/MM0_d N_WL<4>_XI4/XI4/MM0_g
+ N_BL<11>_XI4/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM1 N_XI4/XI4/NET33_XI4/XI4/MM1_d N_XI4/XI4/NET34_XI4/XI4/MM1_g
+ N_VSS_XI4/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM9 N_XI4/XI4/NET36_XI4/XI4/MM9_d N_WL<5>_XI4/XI4/MM9_g
+ N_BL<11>_XI4/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM6 N_XI4/XI4/NET35_XI4/XI4/MM6_d N_XI4/XI4/NET36_XI4/XI4/MM6_g
+ N_VSS_XI4/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM7 N_XI4/XI4/NET36_XI4/XI4/MM7_d N_XI4/XI4/NET35_XI4/XI4/MM7_g
+ N_VSS_XI4/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM8 N_XI4/XI4/NET35_XI4/XI4/MM8_d N_WL<5>_XI4/XI4/MM8_g
+ N_BLN<11>_XI4/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI4/MM5 N_XI4/XI4/NET34_XI4/XI4/MM5_d N_XI4/XI4/NET33_XI4/XI4/MM5_g
+ N_VDD_XI4/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI4/MM4 N_XI4/XI4/NET33_XI4/XI4/MM4_d N_XI4/XI4/NET34_XI4/XI4/MM4_g
+ N_VDD_XI4/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI4/MM10 N_XI4/XI4/NET35_XI4/XI4/MM10_d N_XI4/XI4/NET36_XI4/XI4/MM10_g
+ N_VDD_XI4/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI4/MM11 N_XI4/XI4/NET36_XI4/XI4/MM11_d N_XI4/XI4/NET35_XI4/XI4/MM11_g
+ N_VDD_XI4/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI5/MM2 N_XI4/XI5/NET34_XI4/XI5/MM2_d N_XI4/XI5/NET33_XI4/XI5/MM2_g
+ N_VSS_XI4/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM3 N_XI4/XI5/NET33_XI4/XI5/MM3_d N_WL<4>_XI4/XI5/MM3_g
+ N_BLN<10>_XI4/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM0 N_XI4/XI5/NET34_XI4/XI5/MM0_d N_WL<4>_XI4/XI5/MM0_g
+ N_BL<10>_XI4/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM1 N_XI4/XI5/NET33_XI4/XI5/MM1_d N_XI4/XI5/NET34_XI4/XI5/MM1_g
+ N_VSS_XI4/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM9 N_XI4/XI5/NET36_XI4/XI5/MM9_d N_WL<5>_XI4/XI5/MM9_g
+ N_BL<10>_XI4/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM6 N_XI4/XI5/NET35_XI4/XI5/MM6_d N_XI4/XI5/NET36_XI4/XI5/MM6_g
+ N_VSS_XI4/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM7 N_XI4/XI5/NET36_XI4/XI5/MM7_d N_XI4/XI5/NET35_XI4/XI5/MM7_g
+ N_VSS_XI4/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM8 N_XI4/XI5/NET35_XI4/XI5/MM8_d N_WL<5>_XI4/XI5/MM8_g
+ N_BLN<10>_XI4/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI5/MM5 N_XI4/XI5/NET34_XI4/XI5/MM5_d N_XI4/XI5/NET33_XI4/XI5/MM5_g
+ N_VDD_XI4/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI5/MM4 N_XI4/XI5/NET33_XI4/XI5/MM4_d N_XI4/XI5/NET34_XI4/XI5/MM4_g
+ N_VDD_XI4/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI5/MM10 N_XI4/XI5/NET35_XI4/XI5/MM10_d N_XI4/XI5/NET36_XI4/XI5/MM10_g
+ N_VDD_XI4/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI5/MM11 N_XI4/XI5/NET36_XI4/XI5/MM11_d N_XI4/XI5/NET35_XI4/XI5/MM11_g
+ N_VDD_XI4/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI6/MM2 N_XI4/XI6/NET34_XI4/XI6/MM2_d N_XI4/XI6/NET33_XI4/XI6/MM2_g
+ N_VSS_XI4/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM3 N_XI4/XI6/NET33_XI4/XI6/MM3_d N_WL<4>_XI4/XI6/MM3_g
+ N_BLN<9>_XI4/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM0 N_XI4/XI6/NET34_XI4/XI6/MM0_d N_WL<4>_XI4/XI6/MM0_g
+ N_BL<9>_XI4/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM1 N_XI4/XI6/NET33_XI4/XI6/MM1_d N_XI4/XI6/NET34_XI4/XI6/MM1_g
+ N_VSS_XI4/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM9 N_XI4/XI6/NET36_XI4/XI6/MM9_d N_WL<5>_XI4/XI6/MM9_g
+ N_BL<9>_XI4/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM6 N_XI4/XI6/NET35_XI4/XI6/MM6_d N_XI4/XI6/NET36_XI4/XI6/MM6_g
+ N_VSS_XI4/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM7 N_XI4/XI6/NET36_XI4/XI6/MM7_d N_XI4/XI6/NET35_XI4/XI6/MM7_g
+ N_VSS_XI4/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM8 N_XI4/XI6/NET35_XI4/XI6/MM8_d N_WL<5>_XI4/XI6/MM8_g
+ N_BLN<9>_XI4/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI6/MM5 N_XI4/XI6/NET34_XI4/XI6/MM5_d N_XI4/XI6/NET33_XI4/XI6/MM5_g
+ N_VDD_XI4/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI6/MM4 N_XI4/XI6/NET33_XI4/XI6/MM4_d N_XI4/XI6/NET34_XI4/XI6/MM4_g
+ N_VDD_XI4/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI6/MM10 N_XI4/XI6/NET35_XI4/XI6/MM10_d N_XI4/XI6/NET36_XI4/XI6/MM10_g
+ N_VDD_XI4/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI6/MM11 N_XI4/XI6/NET36_XI4/XI6/MM11_d N_XI4/XI6/NET35_XI4/XI6/MM11_g
+ N_VDD_XI4/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI7/MM2 N_XI4/XI7/NET34_XI4/XI7/MM2_d N_XI4/XI7/NET33_XI4/XI7/MM2_g
+ N_VSS_XI4/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM3 N_XI4/XI7/NET33_XI4/XI7/MM3_d N_WL<4>_XI4/XI7/MM3_g
+ N_BLN<8>_XI4/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM0 N_XI4/XI7/NET34_XI4/XI7/MM0_d N_WL<4>_XI4/XI7/MM0_g
+ N_BL<8>_XI4/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM1 N_XI4/XI7/NET33_XI4/XI7/MM1_d N_XI4/XI7/NET34_XI4/XI7/MM1_g
+ N_VSS_XI4/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM9 N_XI4/XI7/NET36_XI4/XI7/MM9_d N_WL<5>_XI4/XI7/MM9_g
+ N_BL<8>_XI4/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM6 N_XI4/XI7/NET35_XI4/XI7/MM6_d N_XI4/XI7/NET36_XI4/XI7/MM6_g
+ N_VSS_XI4/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM7 N_XI4/XI7/NET36_XI4/XI7/MM7_d N_XI4/XI7/NET35_XI4/XI7/MM7_g
+ N_VSS_XI4/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM8 N_XI4/XI7/NET35_XI4/XI7/MM8_d N_WL<5>_XI4/XI7/MM8_g
+ N_BLN<8>_XI4/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI7/MM5 N_XI4/XI7/NET34_XI4/XI7/MM5_d N_XI4/XI7/NET33_XI4/XI7/MM5_g
+ N_VDD_XI4/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI7/MM4 N_XI4/XI7/NET33_XI4/XI7/MM4_d N_XI4/XI7/NET34_XI4/XI7/MM4_g
+ N_VDD_XI4/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI7/MM10 N_XI4/XI7/NET35_XI4/XI7/MM10_d N_XI4/XI7/NET36_XI4/XI7/MM10_g
+ N_VDD_XI4/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI7/MM11 N_XI4/XI7/NET36_XI4/XI7/MM11_d N_XI4/XI7/NET35_XI4/XI7/MM11_g
+ N_VDD_XI4/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI8/MM2 N_XI4/XI8/NET34_XI4/XI8/MM2_d N_XI4/XI8/NET33_XI4/XI8/MM2_g
+ N_VSS_XI4/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM3 N_XI4/XI8/NET33_XI4/XI8/MM3_d N_WL<4>_XI4/XI8/MM3_g
+ N_BLN<7>_XI4/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM0 N_XI4/XI8/NET34_XI4/XI8/MM0_d N_WL<4>_XI4/XI8/MM0_g
+ N_BL<7>_XI4/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM1 N_XI4/XI8/NET33_XI4/XI8/MM1_d N_XI4/XI8/NET34_XI4/XI8/MM1_g
+ N_VSS_XI4/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM9 N_XI4/XI8/NET36_XI4/XI8/MM9_d N_WL<5>_XI4/XI8/MM9_g
+ N_BL<7>_XI4/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM6 N_XI4/XI8/NET35_XI4/XI8/MM6_d N_XI4/XI8/NET36_XI4/XI8/MM6_g
+ N_VSS_XI4/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM7 N_XI4/XI8/NET36_XI4/XI8/MM7_d N_XI4/XI8/NET35_XI4/XI8/MM7_g
+ N_VSS_XI4/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM8 N_XI4/XI8/NET35_XI4/XI8/MM8_d N_WL<5>_XI4/XI8/MM8_g
+ N_BLN<7>_XI4/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI8/MM5 N_XI4/XI8/NET34_XI4/XI8/MM5_d N_XI4/XI8/NET33_XI4/XI8/MM5_g
+ N_VDD_XI4/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI8/MM4 N_XI4/XI8/NET33_XI4/XI8/MM4_d N_XI4/XI8/NET34_XI4/XI8/MM4_g
+ N_VDD_XI4/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI8/MM10 N_XI4/XI8/NET35_XI4/XI8/MM10_d N_XI4/XI8/NET36_XI4/XI8/MM10_g
+ N_VDD_XI4/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI8/MM11 N_XI4/XI8/NET36_XI4/XI8/MM11_d N_XI4/XI8/NET35_XI4/XI8/MM11_g
+ N_VDD_XI4/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI9/MM2 N_XI4/XI9/NET34_XI4/XI9/MM2_d N_XI4/XI9/NET33_XI4/XI9/MM2_g
+ N_VSS_XI4/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM3 N_XI4/XI9/NET33_XI4/XI9/MM3_d N_WL<4>_XI4/XI9/MM3_g
+ N_BLN<6>_XI4/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM0 N_XI4/XI9/NET34_XI4/XI9/MM0_d N_WL<4>_XI4/XI9/MM0_g
+ N_BL<6>_XI4/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM1 N_XI4/XI9/NET33_XI4/XI9/MM1_d N_XI4/XI9/NET34_XI4/XI9/MM1_g
+ N_VSS_XI4/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM9 N_XI4/XI9/NET36_XI4/XI9/MM9_d N_WL<5>_XI4/XI9/MM9_g
+ N_BL<6>_XI4/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM6 N_XI4/XI9/NET35_XI4/XI9/MM6_d N_XI4/XI9/NET36_XI4/XI9/MM6_g
+ N_VSS_XI4/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM7 N_XI4/XI9/NET36_XI4/XI9/MM7_d N_XI4/XI9/NET35_XI4/XI9/MM7_g
+ N_VSS_XI4/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM8 N_XI4/XI9/NET35_XI4/XI9/MM8_d N_WL<5>_XI4/XI9/MM8_g
+ N_BLN<6>_XI4/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI9/MM5 N_XI4/XI9/NET34_XI4/XI9/MM5_d N_XI4/XI9/NET33_XI4/XI9/MM5_g
+ N_VDD_XI4/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI9/MM4 N_XI4/XI9/NET33_XI4/XI9/MM4_d N_XI4/XI9/NET34_XI4/XI9/MM4_g
+ N_VDD_XI4/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI9/MM10 N_XI4/XI9/NET35_XI4/XI9/MM10_d N_XI4/XI9/NET36_XI4/XI9/MM10_g
+ N_VDD_XI4/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI9/MM11 N_XI4/XI9/NET36_XI4/XI9/MM11_d N_XI4/XI9/NET35_XI4/XI9/MM11_g
+ N_VDD_XI4/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI10/MM2 N_XI4/XI10/NET34_XI4/XI10/MM2_d N_XI4/XI10/NET33_XI4/XI10/MM2_g
+ N_VSS_XI4/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI10/MM3 N_XI4/XI10/NET33_XI4/XI10/MM3_d N_WL<4>_XI4/XI10/MM3_g
+ N_BLN<5>_XI4/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI10/MM0 N_XI4/XI10/NET34_XI4/XI10/MM0_d N_WL<4>_XI4/XI10/MM0_g
+ N_BL<5>_XI4/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI10/MM1 N_XI4/XI10/NET33_XI4/XI10/MM1_d N_XI4/XI10/NET34_XI4/XI10/MM1_g
+ N_VSS_XI4/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI10/MM9 N_XI4/XI10/NET36_XI4/XI10/MM9_d N_WL<5>_XI4/XI10/MM9_g
+ N_BL<5>_XI4/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI10/MM6 N_XI4/XI10/NET35_XI4/XI10/MM6_d N_XI4/XI10/NET36_XI4/XI10/MM6_g
+ N_VSS_XI4/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI10/MM7 N_XI4/XI10/NET36_XI4/XI10/MM7_d N_XI4/XI10/NET35_XI4/XI10/MM7_g
+ N_VSS_XI4/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI10/MM8 N_XI4/XI10/NET35_XI4/XI10/MM8_d N_WL<5>_XI4/XI10/MM8_g
+ N_BLN<5>_XI4/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI10/MM5 N_XI4/XI10/NET34_XI4/XI10/MM5_d N_XI4/XI10/NET33_XI4/XI10/MM5_g
+ N_VDD_XI4/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI10/MM4 N_XI4/XI10/NET33_XI4/XI10/MM4_d N_XI4/XI10/NET34_XI4/XI10/MM4_g
+ N_VDD_XI4/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI10/MM10 N_XI4/XI10/NET35_XI4/XI10/MM10_d N_XI4/XI10/NET36_XI4/XI10/MM10_g
+ N_VDD_XI4/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI10/MM11 N_XI4/XI10/NET36_XI4/XI10/MM11_d N_XI4/XI10/NET35_XI4/XI10/MM11_g
+ N_VDD_XI4/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI11/MM2 N_XI4/XI11/NET34_XI4/XI11/MM2_d N_XI4/XI11/NET33_XI4/XI11/MM2_g
+ N_VSS_XI4/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI11/MM3 N_XI4/XI11/NET33_XI4/XI11/MM3_d N_WL<4>_XI4/XI11/MM3_g
+ N_BLN<4>_XI4/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI11/MM0 N_XI4/XI11/NET34_XI4/XI11/MM0_d N_WL<4>_XI4/XI11/MM0_g
+ N_BL<4>_XI4/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI11/MM1 N_XI4/XI11/NET33_XI4/XI11/MM1_d N_XI4/XI11/NET34_XI4/XI11/MM1_g
+ N_VSS_XI4/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI11/MM9 N_XI4/XI11/NET36_XI4/XI11/MM9_d N_WL<5>_XI4/XI11/MM9_g
+ N_BL<4>_XI4/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI11/MM6 N_XI4/XI11/NET35_XI4/XI11/MM6_d N_XI4/XI11/NET36_XI4/XI11/MM6_g
+ N_VSS_XI4/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI11/MM7 N_XI4/XI11/NET36_XI4/XI11/MM7_d N_XI4/XI11/NET35_XI4/XI11/MM7_g
+ N_VSS_XI4/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI11/MM8 N_XI4/XI11/NET35_XI4/XI11/MM8_d N_WL<5>_XI4/XI11/MM8_g
+ N_BLN<4>_XI4/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI11/MM5 N_XI4/XI11/NET34_XI4/XI11/MM5_d N_XI4/XI11/NET33_XI4/XI11/MM5_g
+ N_VDD_XI4/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI11/MM4 N_XI4/XI11/NET33_XI4/XI11/MM4_d N_XI4/XI11/NET34_XI4/XI11/MM4_g
+ N_VDD_XI4/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI11/MM10 N_XI4/XI11/NET35_XI4/XI11/MM10_d N_XI4/XI11/NET36_XI4/XI11/MM10_g
+ N_VDD_XI4/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI11/MM11 N_XI4/XI11/NET36_XI4/XI11/MM11_d N_XI4/XI11/NET35_XI4/XI11/MM11_g
+ N_VDD_XI4/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI12/MM2 N_XI4/XI12/NET34_XI4/XI12/MM2_d N_XI4/XI12/NET33_XI4/XI12/MM2_g
+ N_VSS_XI4/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI12/MM3 N_XI4/XI12/NET33_XI4/XI12/MM3_d N_WL<4>_XI4/XI12/MM3_g
+ N_BLN<3>_XI4/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI12/MM0 N_XI4/XI12/NET34_XI4/XI12/MM0_d N_WL<4>_XI4/XI12/MM0_g
+ N_BL<3>_XI4/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI12/MM1 N_XI4/XI12/NET33_XI4/XI12/MM1_d N_XI4/XI12/NET34_XI4/XI12/MM1_g
+ N_VSS_XI4/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI12/MM9 N_XI4/XI12/NET36_XI4/XI12/MM9_d N_WL<5>_XI4/XI12/MM9_g
+ N_BL<3>_XI4/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI12/MM6 N_XI4/XI12/NET35_XI4/XI12/MM6_d N_XI4/XI12/NET36_XI4/XI12/MM6_g
+ N_VSS_XI4/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI12/MM7 N_XI4/XI12/NET36_XI4/XI12/MM7_d N_XI4/XI12/NET35_XI4/XI12/MM7_g
+ N_VSS_XI4/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI12/MM8 N_XI4/XI12/NET35_XI4/XI12/MM8_d N_WL<5>_XI4/XI12/MM8_g
+ N_BLN<3>_XI4/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI12/MM5 N_XI4/XI12/NET34_XI4/XI12/MM5_d N_XI4/XI12/NET33_XI4/XI12/MM5_g
+ N_VDD_XI4/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI12/MM4 N_XI4/XI12/NET33_XI4/XI12/MM4_d N_XI4/XI12/NET34_XI4/XI12/MM4_g
+ N_VDD_XI4/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI12/MM10 N_XI4/XI12/NET35_XI4/XI12/MM10_d N_XI4/XI12/NET36_XI4/XI12/MM10_g
+ N_VDD_XI4/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI12/MM11 N_XI4/XI12/NET36_XI4/XI12/MM11_d N_XI4/XI12/NET35_XI4/XI12/MM11_g
+ N_VDD_XI4/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI13/MM2 N_XI4/XI13/NET34_XI4/XI13/MM2_d N_XI4/XI13/NET33_XI4/XI13/MM2_g
+ N_VSS_XI4/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI13/MM3 N_XI4/XI13/NET33_XI4/XI13/MM3_d N_WL<4>_XI4/XI13/MM3_g
+ N_BLN<2>_XI4/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI13/MM0 N_XI4/XI13/NET34_XI4/XI13/MM0_d N_WL<4>_XI4/XI13/MM0_g
+ N_BL<2>_XI4/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI13/MM1 N_XI4/XI13/NET33_XI4/XI13/MM1_d N_XI4/XI13/NET34_XI4/XI13/MM1_g
+ N_VSS_XI4/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI13/MM9 N_XI4/XI13/NET36_XI4/XI13/MM9_d N_WL<5>_XI4/XI13/MM9_g
+ N_BL<2>_XI4/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI13/MM6 N_XI4/XI13/NET35_XI4/XI13/MM6_d N_XI4/XI13/NET36_XI4/XI13/MM6_g
+ N_VSS_XI4/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI13/MM7 N_XI4/XI13/NET36_XI4/XI13/MM7_d N_XI4/XI13/NET35_XI4/XI13/MM7_g
+ N_VSS_XI4/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI13/MM8 N_XI4/XI13/NET35_XI4/XI13/MM8_d N_WL<5>_XI4/XI13/MM8_g
+ N_BLN<2>_XI4/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI13/MM5 N_XI4/XI13/NET34_XI4/XI13/MM5_d N_XI4/XI13/NET33_XI4/XI13/MM5_g
+ N_VDD_XI4/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI13/MM4 N_XI4/XI13/NET33_XI4/XI13/MM4_d N_XI4/XI13/NET34_XI4/XI13/MM4_g
+ N_VDD_XI4/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI13/MM10 N_XI4/XI13/NET35_XI4/XI13/MM10_d N_XI4/XI13/NET36_XI4/XI13/MM10_g
+ N_VDD_XI4/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI13/MM11 N_XI4/XI13/NET36_XI4/XI13/MM11_d N_XI4/XI13/NET35_XI4/XI13/MM11_g
+ N_VDD_XI4/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI14/MM2 N_XI4/XI14/NET34_XI4/XI14/MM2_d N_XI4/XI14/NET33_XI4/XI14/MM2_g
+ N_VSS_XI4/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI14/MM3 N_XI4/XI14/NET33_XI4/XI14/MM3_d N_WL<4>_XI4/XI14/MM3_g
+ N_BLN<1>_XI4/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI14/MM0 N_XI4/XI14/NET34_XI4/XI14/MM0_d N_WL<4>_XI4/XI14/MM0_g
+ N_BL<1>_XI4/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI14/MM1 N_XI4/XI14/NET33_XI4/XI14/MM1_d N_XI4/XI14/NET34_XI4/XI14/MM1_g
+ N_VSS_XI4/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI14/MM9 N_XI4/XI14/NET36_XI4/XI14/MM9_d N_WL<5>_XI4/XI14/MM9_g
+ N_BL<1>_XI4/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI14/MM6 N_XI4/XI14/NET35_XI4/XI14/MM6_d N_XI4/XI14/NET36_XI4/XI14/MM6_g
+ N_VSS_XI4/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI14/MM7 N_XI4/XI14/NET36_XI4/XI14/MM7_d N_XI4/XI14/NET35_XI4/XI14/MM7_g
+ N_VSS_XI4/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI14/MM8 N_XI4/XI14/NET35_XI4/XI14/MM8_d N_WL<5>_XI4/XI14/MM8_g
+ N_BLN<1>_XI4/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI14/MM5 N_XI4/XI14/NET34_XI4/XI14/MM5_d N_XI4/XI14/NET33_XI4/XI14/MM5_g
+ N_VDD_XI4/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI14/MM4 N_XI4/XI14/NET33_XI4/XI14/MM4_d N_XI4/XI14/NET34_XI4/XI14/MM4_g
+ N_VDD_XI4/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI14/MM10 N_XI4/XI14/NET35_XI4/XI14/MM10_d N_XI4/XI14/NET36_XI4/XI14/MM10_g
+ N_VDD_XI4/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI14/MM11 N_XI4/XI14/NET36_XI4/XI14/MM11_d N_XI4/XI14/NET35_XI4/XI14/MM11_g
+ N_VDD_XI4/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI15/MM2 N_XI4/XI15/NET34_XI4/XI15/MM2_d N_XI4/XI15/NET33_XI4/XI15/MM2_g
+ N_VSS_XI4/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI15/MM3 N_XI4/XI15/NET33_XI4/XI15/MM3_d N_WL<4>_XI4/XI15/MM3_g
+ N_BLN<0>_XI4/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI15/MM0 N_XI4/XI15/NET34_XI4/XI15/MM0_d N_WL<4>_XI4/XI15/MM0_g
+ N_BL<0>_XI4/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI15/MM1 N_XI4/XI15/NET33_XI4/XI15/MM1_d N_XI4/XI15/NET34_XI4/XI15/MM1_g
+ N_VSS_XI4/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI15/MM9 N_XI4/XI15/NET36_XI4/XI15/MM9_d N_WL<5>_XI4/XI15/MM9_g
+ N_BL<0>_XI4/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI15/MM6 N_XI4/XI15/NET35_XI4/XI15/MM6_d N_XI4/XI15/NET36_XI4/XI15/MM6_g
+ N_VSS_XI4/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI15/MM7 N_XI4/XI15/NET36_XI4/XI15/MM7_d N_XI4/XI15/NET35_XI4/XI15/MM7_g
+ N_VSS_XI4/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/XI15/MM8 N_XI4/XI15/NET35_XI4/XI15/MM8_d N_WL<5>_XI4/XI15/MM8_g
+ N_BLN<0>_XI4/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI4/XI15/MM5 N_XI4/XI15/NET34_XI4/XI15/MM5_d N_XI4/XI15/NET33_XI4/XI15/MM5_g
+ N_VDD_XI4/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI15/MM4 N_XI4/XI15/NET33_XI4/XI15/MM4_d N_XI4/XI15/NET34_XI4/XI15/MM4_g
+ N_VDD_XI4/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI15/MM10 N_XI4/XI15/NET35_XI4/XI15/MM10_d N_XI4/XI15/NET36_XI4/XI15/MM10_g
+ N_VDD_XI4/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/XI15/MM11 N_XI4/XI15/NET36_XI4/XI15/MM11_d N_XI4/XI15/NET35_XI4/XI15/MM11_g
+ N_VDD_XI4/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI0/MM2 N_XI5/XI0/NET34_XI5/XI0/MM2_d N_XI5/XI0/NET33_XI5/XI0/MM2_g
+ N_VSS_XI5/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM3 N_XI5/XI0/NET33_XI5/XI0/MM3_d N_WL<6>_XI5/XI0/MM3_g
+ N_BLN<15>_XI5/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM0 N_XI5/XI0/NET34_XI5/XI0/MM0_d N_WL<6>_XI5/XI0/MM0_g
+ N_BL<15>_XI5/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM1 N_XI5/XI0/NET33_XI5/XI0/MM1_d N_XI5/XI0/NET34_XI5/XI0/MM1_g
+ N_VSS_XI5/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM9 N_XI5/XI0/NET36_XI5/XI0/MM9_d N_WL<7>_XI5/XI0/MM9_g
+ N_BL<15>_XI5/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM6 N_XI5/XI0/NET35_XI5/XI0/MM6_d N_XI5/XI0/NET36_XI5/XI0/MM6_g
+ N_VSS_XI5/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM7 N_XI5/XI0/NET36_XI5/XI0/MM7_d N_XI5/XI0/NET35_XI5/XI0/MM7_g
+ N_VSS_XI5/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM8 N_XI5/XI0/NET35_XI5/XI0/MM8_d N_WL<7>_XI5/XI0/MM8_g
+ N_BLN<15>_XI5/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI0/MM5 N_XI5/XI0/NET34_XI5/XI0/MM5_d N_XI5/XI0/NET33_XI5/XI0/MM5_g
+ N_VDD_XI5/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI0/MM4 N_XI5/XI0/NET33_XI5/XI0/MM4_d N_XI5/XI0/NET34_XI5/XI0/MM4_g
+ N_VDD_XI5/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI0/MM10 N_XI5/XI0/NET35_XI5/XI0/MM10_d N_XI5/XI0/NET36_XI5/XI0/MM10_g
+ N_VDD_XI5/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI0/MM11 N_XI5/XI0/NET36_XI5/XI0/MM11_d N_XI5/XI0/NET35_XI5/XI0/MM11_g
+ N_VDD_XI5/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI1/MM2 N_XI5/XI1/NET34_XI5/XI1/MM2_d N_XI5/XI1/NET33_XI5/XI1/MM2_g
+ N_VSS_XI5/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM3 N_XI5/XI1/NET33_XI5/XI1/MM3_d N_WL<6>_XI5/XI1/MM3_g
+ N_BLN<14>_XI5/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM0 N_XI5/XI1/NET34_XI5/XI1/MM0_d N_WL<6>_XI5/XI1/MM0_g
+ N_BL<14>_XI5/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM1 N_XI5/XI1/NET33_XI5/XI1/MM1_d N_XI5/XI1/NET34_XI5/XI1/MM1_g
+ N_VSS_XI5/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM9 N_XI5/XI1/NET36_XI5/XI1/MM9_d N_WL<7>_XI5/XI1/MM9_g
+ N_BL<14>_XI5/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM6 N_XI5/XI1/NET35_XI5/XI1/MM6_d N_XI5/XI1/NET36_XI5/XI1/MM6_g
+ N_VSS_XI5/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM7 N_XI5/XI1/NET36_XI5/XI1/MM7_d N_XI5/XI1/NET35_XI5/XI1/MM7_g
+ N_VSS_XI5/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM8 N_XI5/XI1/NET35_XI5/XI1/MM8_d N_WL<7>_XI5/XI1/MM8_g
+ N_BLN<14>_XI5/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI1/MM5 N_XI5/XI1/NET34_XI5/XI1/MM5_d N_XI5/XI1/NET33_XI5/XI1/MM5_g
+ N_VDD_XI5/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI1/MM4 N_XI5/XI1/NET33_XI5/XI1/MM4_d N_XI5/XI1/NET34_XI5/XI1/MM4_g
+ N_VDD_XI5/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI1/MM10 N_XI5/XI1/NET35_XI5/XI1/MM10_d N_XI5/XI1/NET36_XI5/XI1/MM10_g
+ N_VDD_XI5/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI1/MM11 N_XI5/XI1/NET36_XI5/XI1/MM11_d N_XI5/XI1/NET35_XI5/XI1/MM11_g
+ N_VDD_XI5/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI2/MM2 N_XI5/XI2/NET34_XI5/XI2/MM2_d N_XI5/XI2/NET33_XI5/XI2/MM2_g
+ N_VSS_XI5/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM3 N_XI5/XI2/NET33_XI5/XI2/MM3_d N_WL<6>_XI5/XI2/MM3_g
+ N_BLN<13>_XI5/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM0 N_XI5/XI2/NET34_XI5/XI2/MM0_d N_WL<6>_XI5/XI2/MM0_g
+ N_BL<13>_XI5/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM1 N_XI5/XI2/NET33_XI5/XI2/MM1_d N_XI5/XI2/NET34_XI5/XI2/MM1_g
+ N_VSS_XI5/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM9 N_XI5/XI2/NET36_XI5/XI2/MM9_d N_WL<7>_XI5/XI2/MM9_g
+ N_BL<13>_XI5/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM6 N_XI5/XI2/NET35_XI5/XI2/MM6_d N_XI5/XI2/NET36_XI5/XI2/MM6_g
+ N_VSS_XI5/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM7 N_XI5/XI2/NET36_XI5/XI2/MM7_d N_XI5/XI2/NET35_XI5/XI2/MM7_g
+ N_VSS_XI5/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM8 N_XI5/XI2/NET35_XI5/XI2/MM8_d N_WL<7>_XI5/XI2/MM8_g
+ N_BLN<13>_XI5/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI2/MM5 N_XI5/XI2/NET34_XI5/XI2/MM5_d N_XI5/XI2/NET33_XI5/XI2/MM5_g
+ N_VDD_XI5/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI2/MM4 N_XI5/XI2/NET33_XI5/XI2/MM4_d N_XI5/XI2/NET34_XI5/XI2/MM4_g
+ N_VDD_XI5/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI2/MM10 N_XI5/XI2/NET35_XI5/XI2/MM10_d N_XI5/XI2/NET36_XI5/XI2/MM10_g
+ N_VDD_XI5/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI2/MM11 N_XI5/XI2/NET36_XI5/XI2/MM11_d N_XI5/XI2/NET35_XI5/XI2/MM11_g
+ N_VDD_XI5/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI3/MM2 N_XI5/XI3/NET34_XI5/XI3/MM2_d N_XI5/XI3/NET33_XI5/XI3/MM2_g
+ N_VSS_XI5/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM3 N_XI5/XI3/NET33_XI5/XI3/MM3_d N_WL<6>_XI5/XI3/MM3_g
+ N_BLN<12>_XI5/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM0 N_XI5/XI3/NET34_XI5/XI3/MM0_d N_WL<6>_XI5/XI3/MM0_g
+ N_BL<12>_XI5/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM1 N_XI5/XI3/NET33_XI5/XI3/MM1_d N_XI5/XI3/NET34_XI5/XI3/MM1_g
+ N_VSS_XI5/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM9 N_XI5/XI3/NET36_XI5/XI3/MM9_d N_WL<7>_XI5/XI3/MM9_g
+ N_BL<12>_XI5/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM6 N_XI5/XI3/NET35_XI5/XI3/MM6_d N_XI5/XI3/NET36_XI5/XI3/MM6_g
+ N_VSS_XI5/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM7 N_XI5/XI3/NET36_XI5/XI3/MM7_d N_XI5/XI3/NET35_XI5/XI3/MM7_g
+ N_VSS_XI5/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM8 N_XI5/XI3/NET35_XI5/XI3/MM8_d N_WL<7>_XI5/XI3/MM8_g
+ N_BLN<12>_XI5/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI3/MM5 N_XI5/XI3/NET34_XI5/XI3/MM5_d N_XI5/XI3/NET33_XI5/XI3/MM5_g
+ N_VDD_XI5/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI3/MM4 N_XI5/XI3/NET33_XI5/XI3/MM4_d N_XI5/XI3/NET34_XI5/XI3/MM4_g
+ N_VDD_XI5/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI3/MM10 N_XI5/XI3/NET35_XI5/XI3/MM10_d N_XI5/XI3/NET36_XI5/XI3/MM10_g
+ N_VDD_XI5/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI3/MM11 N_XI5/XI3/NET36_XI5/XI3/MM11_d N_XI5/XI3/NET35_XI5/XI3/MM11_g
+ N_VDD_XI5/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI4/MM2 N_XI5/XI4/NET34_XI5/XI4/MM2_d N_XI5/XI4/NET33_XI5/XI4/MM2_g
+ N_VSS_XI5/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM3 N_XI5/XI4/NET33_XI5/XI4/MM3_d N_WL<6>_XI5/XI4/MM3_g
+ N_BLN<11>_XI5/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM0 N_XI5/XI4/NET34_XI5/XI4/MM0_d N_WL<6>_XI5/XI4/MM0_g
+ N_BL<11>_XI5/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM1 N_XI5/XI4/NET33_XI5/XI4/MM1_d N_XI5/XI4/NET34_XI5/XI4/MM1_g
+ N_VSS_XI5/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM9 N_XI5/XI4/NET36_XI5/XI4/MM9_d N_WL<7>_XI5/XI4/MM9_g
+ N_BL<11>_XI5/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM6 N_XI5/XI4/NET35_XI5/XI4/MM6_d N_XI5/XI4/NET36_XI5/XI4/MM6_g
+ N_VSS_XI5/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM7 N_XI5/XI4/NET36_XI5/XI4/MM7_d N_XI5/XI4/NET35_XI5/XI4/MM7_g
+ N_VSS_XI5/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM8 N_XI5/XI4/NET35_XI5/XI4/MM8_d N_WL<7>_XI5/XI4/MM8_g
+ N_BLN<11>_XI5/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI4/MM5 N_XI5/XI4/NET34_XI5/XI4/MM5_d N_XI5/XI4/NET33_XI5/XI4/MM5_g
+ N_VDD_XI5/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI4/MM4 N_XI5/XI4/NET33_XI5/XI4/MM4_d N_XI5/XI4/NET34_XI5/XI4/MM4_g
+ N_VDD_XI5/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI4/MM10 N_XI5/XI4/NET35_XI5/XI4/MM10_d N_XI5/XI4/NET36_XI5/XI4/MM10_g
+ N_VDD_XI5/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI4/MM11 N_XI5/XI4/NET36_XI5/XI4/MM11_d N_XI5/XI4/NET35_XI5/XI4/MM11_g
+ N_VDD_XI5/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI5/MM2 N_XI5/XI5/NET34_XI5/XI5/MM2_d N_XI5/XI5/NET33_XI5/XI5/MM2_g
+ N_VSS_XI5/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM3 N_XI5/XI5/NET33_XI5/XI5/MM3_d N_WL<6>_XI5/XI5/MM3_g
+ N_BLN<10>_XI5/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM0 N_XI5/XI5/NET34_XI5/XI5/MM0_d N_WL<6>_XI5/XI5/MM0_g
+ N_BL<10>_XI5/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM1 N_XI5/XI5/NET33_XI5/XI5/MM1_d N_XI5/XI5/NET34_XI5/XI5/MM1_g
+ N_VSS_XI5/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM9 N_XI5/XI5/NET36_XI5/XI5/MM9_d N_WL<7>_XI5/XI5/MM9_g
+ N_BL<10>_XI5/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM6 N_XI5/XI5/NET35_XI5/XI5/MM6_d N_XI5/XI5/NET36_XI5/XI5/MM6_g
+ N_VSS_XI5/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM7 N_XI5/XI5/NET36_XI5/XI5/MM7_d N_XI5/XI5/NET35_XI5/XI5/MM7_g
+ N_VSS_XI5/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM8 N_XI5/XI5/NET35_XI5/XI5/MM8_d N_WL<7>_XI5/XI5/MM8_g
+ N_BLN<10>_XI5/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI5/MM5 N_XI5/XI5/NET34_XI5/XI5/MM5_d N_XI5/XI5/NET33_XI5/XI5/MM5_g
+ N_VDD_XI5/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI5/MM4 N_XI5/XI5/NET33_XI5/XI5/MM4_d N_XI5/XI5/NET34_XI5/XI5/MM4_g
+ N_VDD_XI5/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI5/MM10 N_XI5/XI5/NET35_XI5/XI5/MM10_d N_XI5/XI5/NET36_XI5/XI5/MM10_g
+ N_VDD_XI5/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI5/MM11 N_XI5/XI5/NET36_XI5/XI5/MM11_d N_XI5/XI5/NET35_XI5/XI5/MM11_g
+ N_VDD_XI5/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI6/MM2 N_XI5/XI6/NET34_XI5/XI6/MM2_d N_XI5/XI6/NET33_XI5/XI6/MM2_g
+ N_VSS_XI5/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM3 N_XI5/XI6/NET33_XI5/XI6/MM3_d N_WL<6>_XI5/XI6/MM3_g
+ N_BLN<9>_XI5/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM0 N_XI5/XI6/NET34_XI5/XI6/MM0_d N_WL<6>_XI5/XI6/MM0_g
+ N_BL<9>_XI5/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM1 N_XI5/XI6/NET33_XI5/XI6/MM1_d N_XI5/XI6/NET34_XI5/XI6/MM1_g
+ N_VSS_XI5/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM9 N_XI5/XI6/NET36_XI5/XI6/MM9_d N_WL<7>_XI5/XI6/MM9_g
+ N_BL<9>_XI5/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM6 N_XI5/XI6/NET35_XI5/XI6/MM6_d N_XI5/XI6/NET36_XI5/XI6/MM6_g
+ N_VSS_XI5/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM7 N_XI5/XI6/NET36_XI5/XI6/MM7_d N_XI5/XI6/NET35_XI5/XI6/MM7_g
+ N_VSS_XI5/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM8 N_XI5/XI6/NET35_XI5/XI6/MM8_d N_WL<7>_XI5/XI6/MM8_g
+ N_BLN<9>_XI5/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI6/MM5 N_XI5/XI6/NET34_XI5/XI6/MM5_d N_XI5/XI6/NET33_XI5/XI6/MM5_g
+ N_VDD_XI5/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI6/MM4 N_XI5/XI6/NET33_XI5/XI6/MM4_d N_XI5/XI6/NET34_XI5/XI6/MM4_g
+ N_VDD_XI5/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI6/MM10 N_XI5/XI6/NET35_XI5/XI6/MM10_d N_XI5/XI6/NET36_XI5/XI6/MM10_g
+ N_VDD_XI5/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI6/MM11 N_XI5/XI6/NET36_XI5/XI6/MM11_d N_XI5/XI6/NET35_XI5/XI6/MM11_g
+ N_VDD_XI5/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI7/MM2 N_XI5/XI7/NET34_XI5/XI7/MM2_d N_XI5/XI7/NET33_XI5/XI7/MM2_g
+ N_VSS_XI5/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM3 N_XI5/XI7/NET33_XI5/XI7/MM3_d N_WL<6>_XI5/XI7/MM3_g
+ N_BLN<8>_XI5/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM0 N_XI5/XI7/NET34_XI5/XI7/MM0_d N_WL<6>_XI5/XI7/MM0_g
+ N_BL<8>_XI5/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM1 N_XI5/XI7/NET33_XI5/XI7/MM1_d N_XI5/XI7/NET34_XI5/XI7/MM1_g
+ N_VSS_XI5/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM9 N_XI5/XI7/NET36_XI5/XI7/MM9_d N_WL<7>_XI5/XI7/MM9_g
+ N_BL<8>_XI5/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM6 N_XI5/XI7/NET35_XI5/XI7/MM6_d N_XI5/XI7/NET36_XI5/XI7/MM6_g
+ N_VSS_XI5/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM7 N_XI5/XI7/NET36_XI5/XI7/MM7_d N_XI5/XI7/NET35_XI5/XI7/MM7_g
+ N_VSS_XI5/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM8 N_XI5/XI7/NET35_XI5/XI7/MM8_d N_WL<7>_XI5/XI7/MM8_g
+ N_BLN<8>_XI5/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI7/MM5 N_XI5/XI7/NET34_XI5/XI7/MM5_d N_XI5/XI7/NET33_XI5/XI7/MM5_g
+ N_VDD_XI5/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI7/MM4 N_XI5/XI7/NET33_XI5/XI7/MM4_d N_XI5/XI7/NET34_XI5/XI7/MM4_g
+ N_VDD_XI5/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI7/MM10 N_XI5/XI7/NET35_XI5/XI7/MM10_d N_XI5/XI7/NET36_XI5/XI7/MM10_g
+ N_VDD_XI5/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI7/MM11 N_XI5/XI7/NET36_XI5/XI7/MM11_d N_XI5/XI7/NET35_XI5/XI7/MM11_g
+ N_VDD_XI5/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI8/MM2 N_XI5/XI8/NET34_XI5/XI8/MM2_d N_XI5/XI8/NET33_XI5/XI8/MM2_g
+ N_VSS_XI5/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM3 N_XI5/XI8/NET33_XI5/XI8/MM3_d N_WL<6>_XI5/XI8/MM3_g
+ N_BLN<7>_XI5/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM0 N_XI5/XI8/NET34_XI5/XI8/MM0_d N_WL<6>_XI5/XI8/MM0_g
+ N_BL<7>_XI5/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM1 N_XI5/XI8/NET33_XI5/XI8/MM1_d N_XI5/XI8/NET34_XI5/XI8/MM1_g
+ N_VSS_XI5/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM9 N_XI5/XI8/NET36_XI5/XI8/MM9_d N_WL<7>_XI5/XI8/MM9_g
+ N_BL<7>_XI5/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM6 N_XI5/XI8/NET35_XI5/XI8/MM6_d N_XI5/XI8/NET36_XI5/XI8/MM6_g
+ N_VSS_XI5/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM7 N_XI5/XI8/NET36_XI5/XI8/MM7_d N_XI5/XI8/NET35_XI5/XI8/MM7_g
+ N_VSS_XI5/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM8 N_XI5/XI8/NET35_XI5/XI8/MM8_d N_WL<7>_XI5/XI8/MM8_g
+ N_BLN<7>_XI5/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI8/MM5 N_XI5/XI8/NET34_XI5/XI8/MM5_d N_XI5/XI8/NET33_XI5/XI8/MM5_g
+ N_VDD_XI5/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI8/MM4 N_XI5/XI8/NET33_XI5/XI8/MM4_d N_XI5/XI8/NET34_XI5/XI8/MM4_g
+ N_VDD_XI5/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI8/MM10 N_XI5/XI8/NET35_XI5/XI8/MM10_d N_XI5/XI8/NET36_XI5/XI8/MM10_g
+ N_VDD_XI5/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI8/MM11 N_XI5/XI8/NET36_XI5/XI8/MM11_d N_XI5/XI8/NET35_XI5/XI8/MM11_g
+ N_VDD_XI5/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI9/MM2 N_XI5/XI9/NET34_XI5/XI9/MM2_d N_XI5/XI9/NET33_XI5/XI9/MM2_g
+ N_VSS_XI5/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM3 N_XI5/XI9/NET33_XI5/XI9/MM3_d N_WL<6>_XI5/XI9/MM3_g
+ N_BLN<6>_XI5/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM0 N_XI5/XI9/NET34_XI5/XI9/MM0_d N_WL<6>_XI5/XI9/MM0_g
+ N_BL<6>_XI5/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM1 N_XI5/XI9/NET33_XI5/XI9/MM1_d N_XI5/XI9/NET34_XI5/XI9/MM1_g
+ N_VSS_XI5/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM9 N_XI5/XI9/NET36_XI5/XI9/MM9_d N_WL<7>_XI5/XI9/MM9_g
+ N_BL<6>_XI5/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM6 N_XI5/XI9/NET35_XI5/XI9/MM6_d N_XI5/XI9/NET36_XI5/XI9/MM6_g
+ N_VSS_XI5/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM7 N_XI5/XI9/NET36_XI5/XI9/MM7_d N_XI5/XI9/NET35_XI5/XI9/MM7_g
+ N_VSS_XI5/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM8 N_XI5/XI9/NET35_XI5/XI9/MM8_d N_WL<7>_XI5/XI9/MM8_g
+ N_BLN<6>_XI5/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI9/MM5 N_XI5/XI9/NET34_XI5/XI9/MM5_d N_XI5/XI9/NET33_XI5/XI9/MM5_g
+ N_VDD_XI5/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI9/MM4 N_XI5/XI9/NET33_XI5/XI9/MM4_d N_XI5/XI9/NET34_XI5/XI9/MM4_g
+ N_VDD_XI5/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI9/MM10 N_XI5/XI9/NET35_XI5/XI9/MM10_d N_XI5/XI9/NET36_XI5/XI9/MM10_g
+ N_VDD_XI5/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI9/MM11 N_XI5/XI9/NET36_XI5/XI9/MM11_d N_XI5/XI9/NET35_XI5/XI9/MM11_g
+ N_VDD_XI5/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI10/MM2 N_XI5/XI10/NET34_XI5/XI10/MM2_d N_XI5/XI10/NET33_XI5/XI10/MM2_g
+ N_VSS_XI5/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI10/MM3 N_XI5/XI10/NET33_XI5/XI10/MM3_d N_WL<6>_XI5/XI10/MM3_g
+ N_BLN<5>_XI5/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI10/MM0 N_XI5/XI10/NET34_XI5/XI10/MM0_d N_WL<6>_XI5/XI10/MM0_g
+ N_BL<5>_XI5/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI10/MM1 N_XI5/XI10/NET33_XI5/XI10/MM1_d N_XI5/XI10/NET34_XI5/XI10/MM1_g
+ N_VSS_XI5/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI10/MM9 N_XI5/XI10/NET36_XI5/XI10/MM9_d N_WL<7>_XI5/XI10/MM9_g
+ N_BL<5>_XI5/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI10/MM6 N_XI5/XI10/NET35_XI5/XI10/MM6_d N_XI5/XI10/NET36_XI5/XI10/MM6_g
+ N_VSS_XI5/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI10/MM7 N_XI5/XI10/NET36_XI5/XI10/MM7_d N_XI5/XI10/NET35_XI5/XI10/MM7_g
+ N_VSS_XI5/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI10/MM8 N_XI5/XI10/NET35_XI5/XI10/MM8_d N_WL<7>_XI5/XI10/MM8_g
+ N_BLN<5>_XI5/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI10/MM5 N_XI5/XI10/NET34_XI5/XI10/MM5_d N_XI5/XI10/NET33_XI5/XI10/MM5_g
+ N_VDD_XI5/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI10/MM4 N_XI5/XI10/NET33_XI5/XI10/MM4_d N_XI5/XI10/NET34_XI5/XI10/MM4_g
+ N_VDD_XI5/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI10/MM10 N_XI5/XI10/NET35_XI5/XI10/MM10_d N_XI5/XI10/NET36_XI5/XI10/MM10_g
+ N_VDD_XI5/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI10/MM11 N_XI5/XI10/NET36_XI5/XI10/MM11_d N_XI5/XI10/NET35_XI5/XI10/MM11_g
+ N_VDD_XI5/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI11/MM2 N_XI5/XI11/NET34_XI5/XI11/MM2_d N_XI5/XI11/NET33_XI5/XI11/MM2_g
+ N_VSS_XI5/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI11/MM3 N_XI5/XI11/NET33_XI5/XI11/MM3_d N_WL<6>_XI5/XI11/MM3_g
+ N_BLN<4>_XI5/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI11/MM0 N_XI5/XI11/NET34_XI5/XI11/MM0_d N_WL<6>_XI5/XI11/MM0_g
+ N_BL<4>_XI5/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI11/MM1 N_XI5/XI11/NET33_XI5/XI11/MM1_d N_XI5/XI11/NET34_XI5/XI11/MM1_g
+ N_VSS_XI5/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI11/MM9 N_XI5/XI11/NET36_XI5/XI11/MM9_d N_WL<7>_XI5/XI11/MM9_g
+ N_BL<4>_XI5/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI11/MM6 N_XI5/XI11/NET35_XI5/XI11/MM6_d N_XI5/XI11/NET36_XI5/XI11/MM6_g
+ N_VSS_XI5/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI11/MM7 N_XI5/XI11/NET36_XI5/XI11/MM7_d N_XI5/XI11/NET35_XI5/XI11/MM7_g
+ N_VSS_XI5/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI11/MM8 N_XI5/XI11/NET35_XI5/XI11/MM8_d N_WL<7>_XI5/XI11/MM8_g
+ N_BLN<4>_XI5/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI11/MM5 N_XI5/XI11/NET34_XI5/XI11/MM5_d N_XI5/XI11/NET33_XI5/XI11/MM5_g
+ N_VDD_XI5/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI11/MM4 N_XI5/XI11/NET33_XI5/XI11/MM4_d N_XI5/XI11/NET34_XI5/XI11/MM4_g
+ N_VDD_XI5/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI11/MM10 N_XI5/XI11/NET35_XI5/XI11/MM10_d N_XI5/XI11/NET36_XI5/XI11/MM10_g
+ N_VDD_XI5/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI11/MM11 N_XI5/XI11/NET36_XI5/XI11/MM11_d N_XI5/XI11/NET35_XI5/XI11/MM11_g
+ N_VDD_XI5/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI12/MM2 N_XI5/XI12/NET34_XI5/XI12/MM2_d N_XI5/XI12/NET33_XI5/XI12/MM2_g
+ N_VSS_XI5/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI12/MM3 N_XI5/XI12/NET33_XI5/XI12/MM3_d N_WL<6>_XI5/XI12/MM3_g
+ N_BLN<3>_XI5/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI12/MM0 N_XI5/XI12/NET34_XI5/XI12/MM0_d N_WL<6>_XI5/XI12/MM0_g
+ N_BL<3>_XI5/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI12/MM1 N_XI5/XI12/NET33_XI5/XI12/MM1_d N_XI5/XI12/NET34_XI5/XI12/MM1_g
+ N_VSS_XI5/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI12/MM9 N_XI5/XI12/NET36_XI5/XI12/MM9_d N_WL<7>_XI5/XI12/MM9_g
+ N_BL<3>_XI5/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI12/MM6 N_XI5/XI12/NET35_XI5/XI12/MM6_d N_XI5/XI12/NET36_XI5/XI12/MM6_g
+ N_VSS_XI5/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI12/MM7 N_XI5/XI12/NET36_XI5/XI12/MM7_d N_XI5/XI12/NET35_XI5/XI12/MM7_g
+ N_VSS_XI5/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI12/MM8 N_XI5/XI12/NET35_XI5/XI12/MM8_d N_WL<7>_XI5/XI12/MM8_g
+ N_BLN<3>_XI5/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI12/MM5 N_XI5/XI12/NET34_XI5/XI12/MM5_d N_XI5/XI12/NET33_XI5/XI12/MM5_g
+ N_VDD_XI5/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI12/MM4 N_XI5/XI12/NET33_XI5/XI12/MM4_d N_XI5/XI12/NET34_XI5/XI12/MM4_g
+ N_VDD_XI5/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI12/MM10 N_XI5/XI12/NET35_XI5/XI12/MM10_d N_XI5/XI12/NET36_XI5/XI12/MM10_g
+ N_VDD_XI5/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI12/MM11 N_XI5/XI12/NET36_XI5/XI12/MM11_d N_XI5/XI12/NET35_XI5/XI12/MM11_g
+ N_VDD_XI5/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI13/MM2 N_XI5/XI13/NET34_XI5/XI13/MM2_d N_XI5/XI13/NET33_XI5/XI13/MM2_g
+ N_VSS_XI5/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI13/MM3 N_XI5/XI13/NET33_XI5/XI13/MM3_d N_WL<6>_XI5/XI13/MM3_g
+ N_BLN<2>_XI5/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI13/MM0 N_XI5/XI13/NET34_XI5/XI13/MM0_d N_WL<6>_XI5/XI13/MM0_g
+ N_BL<2>_XI5/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI13/MM1 N_XI5/XI13/NET33_XI5/XI13/MM1_d N_XI5/XI13/NET34_XI5/XI13/MM1_g
+ N_VSS_XI5/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI13/MM9 N_XI5/XI13/NET36_XI5/XI13/MM9_d N_WL<7>_XI5/XI13/MM9_g
+ N_BL<2>_XI5/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI13/MM6 N_XI5/XI13/NET35_XI5/XI13/MM6_d N_XI5/XI13/NET36_XI5/XI13/MM6_g
+ N_VSS_XI5/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI13/MM7 N_XI5/XI13/NET36_XI5/XI13/MM7_d N_XI5/XI13/NET35_XI5/XI13/MM7_g
+ N_VSS_XI5/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI13/MM8 N_XI5/XI13/NET35_XI5/XI13/MM8_d N_WL<7>_XI5/XI13/MM8_g
+ N_BLN<2>_XI5/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI13/MM5 N_XI5/XI13/NET34_XI5/XI13/MM5_d N_XI5/XI13/NET33_XI5/XI13/MM5_g
+ N_VDD_XI5/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI13/MM4 N_XI5/XI13/NET33_XI5/XI13/MM4_d N_XI5/XI13/NET34_XI5/XI13/MM4_g
+ N_VDD_XI5/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI13/MM10 N_XI5/XI13/NET35_XI5/XI13/MM10_d N_XI5/XI13/NET36_XI5/XI13/MM10_g
+ N_VDD_XI5/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI13/MM11 N_XI5/XI13/NET36_XI5/XI13/MM11_d N_XI5/XI13/NET35_XI5/XI13/MM11_g
+ N_VDD_XI5/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI14/MM2 N_XI5/XI14/NET34_XI5/XI14/MM2_d N_XI5/XI14/NET33_XI5/XI14/MM2_g
+ N_VSS_XI5/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI14/MM3 N_XI5/XI14/NET33_XI5/XI14/MM3_d N_WL<6>_XI5/XI14/MM3_g
+ N_BLN<1>_XI5/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI14/MM0 N_XI5/XI14/NET34_XI5/XI14/MM0_d N_WL<6>_XI5/XI14/MM0_g
+ N_BL<1>_XI5/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI14/MM1 N_XI5/XI14/NET33_XI5/XI14/MM1_d N_XI5/XI14/NET34_XI5/XI14/MM1_g
+ N_VSS_XI5/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI14/MM9 N_XI5/XI14/NET36_XI5/XI14/MM9_d N_WL<7>_XI5/XI14/MM9_g
+ N_BL<1>_XI5/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI14/MM6 N_XI5/XI14/NET35_XI5/XI14/MM6_d N_XI5/XI14/NET36_XI5/XI14/MM6_g
+ N_VSS_XI5/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI14/MM7 N_XI5/XI14/NET36_XI5/XI14/MM7_d N_XI5/XI14/NET35_XI5/XI14/MM7_g
+ N_VSS_XI5/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI14/MM8 N_XI5/XI14/NET35_XI5/XI14/MM8_d N_WL<7>_XI5/XI14/MM8_g
+ N_BLN<1>_XI5/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI14/MM5 N_XI5/XI14/NET34_XI5/XI14/MM5_d N_XI5/XI14/NET33_XI5/XI14/MM5_g
+ N_VDD_XI5/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI14/MM4 N_XI5/XI14/NET33_XI5/XI14/MM4_d N_XI5/XI14/NET34_XI5/XI14/MM4_g
+ N_VDD_XI5/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI14/MM10 N_XI5/XI14/NET35_XI5/XI14/MM10_d N_XI5/XI14/NET36_XI5/XI14/MM10_g
+ N_VDD_XI5/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI14/MM11 N_XI5/XI14/NET36_XI5/XI14/MM11_d N_XI5/XI14/NET35_XI5/XI14/MM11_g
+ N_VDD_XI5/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI15/MM2 N_XI5/XI15/NET34_XI5/XI15/MM2_d N_XI5/XI15/NET33_XI5/XI15/MM2_g
+ N_VSS_XI5/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI15/MM3 N_XI5/XI15/NET33_XI5/XI15/MM3_d N_WL<6>_XI5/XI15/MM3_g
+ N_BLN<0>_XI5/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI15/MM0 N_XI5/XI15/NET34_XI5/XI15/MM0_d N_WL<6>_XI5/XI15/MM0_g
+ N_BL<0>_XI5/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI15/MM1 N_XI5/XI15/NET33_XI5/XI15/MM1_d N_XI5/XI15/NET34_XI5/XI15/MM1_g
+ N_VSS_XI5/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI15/MM9 N_XI5/XI15/NET36_XI5/XI15/MM9_d N_WL<7>_XI5/XI15/MM9_g
+ N_BL<0>_XI5/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI15/MM6 N_XI5/XI15/NET35_XI5/XI15/MM6_d N_XI5/XI15/NET36_XI5/XI15/MM6_g
+ N_VSS_XI5/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI15/MM7 N_XI5/XI15/NET36_XI5/XI15/MM7_d N_XI5/XI15/NET35_XI5/XI15/MM7_g
+ N_VSS_XI5/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/XI15/MM8 N_XI5/XI15/NET35_XI5/XI15/MM8_d N_WL<7>_XI5/XI15/MM8_g
+ N_BLN<0>_XI5/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI5/XI15/MM5 N_XI5/XI15/NET34_XI5/XI15/MM5_d N_XI5/XI15/NET33_XI5/XI15/MM5_g
+ N_VDD_XI5/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI15/MM4 N_XI5/XI15/NET33_XI5/XI15/MM4_d N_XI5/XI15/NET34_XI5/XI15/MM4_g
+ N_VDD_XI5/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI15/MM10 N_XI5/XI15/NET35_XI5/XI15/MM10_d N_XI5/XI15/NET36_XI5/XI15/MM10_g
+ N_VDD_XI5/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/XI15/MM11 N_XI5/XI15/NET36_XI5/XI15/MM11_d N_XI5/XI15/NET35_XI5/XI15/MM11_g
+ N_VDD_XI5/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI0/MM2 N_XI6/XI0/NET34_XI6/XI0/MM2_d N_XI6/XI0/NET33_XI6/XI0/MM2_g
+ N_VSS_XI6/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM3 N_XI6/XI0/NET33_XI6/XI0/MM3_d N_WL<8>_XI6/XI0/MM3_g
+ N_BLN<15>_XI6/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM0 N_XI6/XI0/NET34_XI6/XI0/MM0_d N_WL<8>_XI6/XI0/MM0_g
+ N_BL<15>_XI6/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM1 N_XI6/XI0/NET33_XI6/XI0/MM1_d N_XI6/XI0/NET34_XI6/XI0/MM1_g
+ N_VSS_XI6/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM9 N_XI6/XI0/NET36_XI6/XI0/MM9_d N_WL<9>_XI6/XI0/MM9_g
+ N_BL<15>_XI6/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM6 N_XI6/XI0/NET35_XI6/XI0/MM6_d N_XI6/XI0/NET36_XI6/XI0/MM6_g
+ N_VSS_XI6/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM7 N_XI6/XI0/NET36_XI6/XI0/MM7_d N_XI6/XI0/NET35_XI6/XI0/MM7_g
+ N_VSS_XI6/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM8 N_XI6/XI0/NET35_XI6/XI0/MM8_d N_WL<9>_XI6/XI0/MM8_g
+ N_BLN<15>_XI6/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI0/MM5 N_XI6/XI0/NET34_XI6/XI0/MM5_d N_XI6/XI0/NET33_XI6/XI0/MM5_g
+ N_VDD_XI6/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI0/MM4 N_XI6/XI0/NET33_XI6/XI0/MM4_d N_XI6/XI0/NET34_XI6/XI0/MM4_g
+ N_VDD_XI6/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI0/MM10 N_XI6/XI0/NET35_XI6/XI0/MM10_d N_XI6/XI0/NET36_XI6/XI0/MM10_g
+ N_VDD_XI6/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI0/MM11 N_XI6/XI0/NET36_XI6/XI0/MM11_d N_XI6/XI0/NET35_XI6/XI0/MM11_g
+ N_VDD_XI6/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI1/MM2 N_XI6/XI1/NET34_XI6/XI1/MM2_d N_XI6/XI1/NET33_XI6/XI1/MM2_g
+ N_VSS_XI6/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM3 N_XI6/XI1/NET33_XI6/XI1/MM3_d N_WL<8>_XI6/XI1/MM3_g
+ N_BLN<14>_XI6/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM0 N_XI6/XI1/NET34_XI6/XI1/MM0_d N_WL<8>_XI6/XI1/MM0_g
+ N_BL<14>_XI6/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM1 N_XI6/XI1/NET33_XI6/XI1/MM1_d N_XI6/XI1/NET34_XI6/XI1/MM1_g
+ N_VSS_XI6/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM9 N_XI6/XI1/NET36_XI6/XI1/MM9_d N_WL<9>_XI6/XI1/MM9_g
+ N_BL<14>_XI6/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM6 N_XI6/XI1/NET35_XI6/XI1/MM6_d N_XI6/XI1/NET36_XI6/XI1/MM6_g
+ N_VSS_XI6/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM7 N_XI6/XI1/NET36_XI6/XI1/MM7_d N_XI6/XI1/NET35_XI6/XI1/MM7_g
+ N_VSS_XI6/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM8 N_XI6/XI1/NET35_XI6/XI1/MM8_d N_WL<9>_XI6/XI1/MM8_g
+ N_BLN<14>_XI6/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI1/MM5 N_XI6/XI1/NET34_XI6/XI1/MM5_d N_XI6/XI1/NET33_XI6/XI1/MM5_g
+ N_VDD_XI6/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI1/MM4 N_XI6/XI1/NET33_XI6/XI1/MM4_d N_XI6/XI1/NET34_XI6/XI1/MM4_g
+ N_VDD_XI6/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI1/MM10 N_XI6/XI1/NET35_XI6/XI1/MM10_d N_XI6/XI1/NET36_XI6/XI1/MM10_g
+ N_VDD_XI6/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI1/MM11 N_XI6/XI1/NET36_XI6/XI1/MM11_d N_XI6/XI1/NET35_XI6/XI1/MM11_g
+ N_VDD_XI6/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI2/MM2 N_XI6/XI2/NET34_XI6/XI2/MM2_d N_XI6/XI2/NET33_XI6/XI2/MM2_g
+ N_VSS_XI6/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM3 N_XI6/XI2/NET33_XI6/XI2/MM3_d N_WL<8>_XI6/XI2/MM3_g
+ N_BLN<13>_XI6/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM0 N_XI6/XI2/NET34_XI6/XI2/MM0_d N_WL<8>_XI6/XI2/MM0_g
+ N_BL<13>_XI6/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM1 N_XI6/XI2/NET33_XI6/XI2/MM1_d N_XI6/XI2/NET34_XI6/XI2/MM1_g
+ N_VSS_XI6/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM9 N_XI6/XI2/NET36_XI6/XI2/MM9_d N_WL<9>_XI6/XI2/MM9_g
+ N_BL<13>_XI6/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM6 N_XI6/XI2/NET35_XI6/XI2/MM6_d N_XI6/XI2/NET36_XI6/XI2/MM6_g
+ N_VSS_XI6/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM7 N_XI6/XI2/NET36_XI6/XI2/MM7_d N_XI6/XI2/NET35_XI6/XI2/MM7_g
+ N_VSS_XI6/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM8 N_XI6/XI2/NET35_XI6/XI2/MM8_d N_WL<9>_XI6/XI2/MM8_g
+ N_BLN<13>_XI6/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI2/MM5 N_XI6/XI2/NET34_XI6/XI2/MM5_d N_XI6/XI2/NET33_XI6/XI2/MM5_g
+ N_VDD_XI6/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI2/MM4 N_XI6/XI2/NET33_XI6/XI2/MM4_d N_XI6/XI2/NET34_XI6/XI2/MM4_g
+ N_VDD_XI6/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI2/MM10 N_XI6/XI2/NET35_XI6/XI2/MM10_d N_XI6/XI2/NET36_XI6/XI2/MM10_g
+ N_VDD_XI6/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI2/MM11 N_XI6/XI2/NET36_XI6/XI2/MM11_d N_XI6/XI2/NET35_XI6/XI2/MM11_g
+ N_VDD_XI6/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI3/MM2 N_XI6/XI3/NET34_XI6/XI3/MM2_d N_XI6/XI3/NET33_XI6/XI3/MM2_g
+ N_VSS_XI6/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM3 N_XI6/XI3/NET33_XI6/XI3/MM3_d N_WL<8>_XI6/XI3/MM3_g
+ N_BLN<12>_XI6/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM0 N_XI6/XI3/NET34_XI6/XI3/MM0_d N_WL<8>_XI6/XI3/MM0_g
+ N_BL<12>_XI6/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM1 N_XI6/XI3/NET33_XI6/XI3/MM1_d N_XI6/XI3/NET34_XI6/XI3/MM1_g
+ N_VSS_XI6/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM9 N_XI6/XI3/NET36_XI6/XI3/MM9_d N_WL<9>_XI6/XI3/MM9_g
+ N_BL<12>_XI6/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM6 N_XI6/XI3/NET35_XI6/XI3/MM6_d N_XI6/XI3/NET36_XI6/XI3/MM6_g
+ N_VSS_XI6/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM7 N_XI6/XI3/NET36_XI6/XI3/MM7_d N_XI6/XI3/NET35_XI6/XI3/MM7_g
+ N_VSS_XI6/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM8 N_XI6/XI3/NET35_XI6/XI3/MM8_d N_WL<9>_XI6/XI3/MM8_g
+ N_BLN<12>_XI6/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI3/MM5 N_XI6/XI3/NET34_XI6/XI3/MM5_d N_XI6/XI3/NET33_XI6/XI3/MM5_g
+ N_VDD_XI6/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI3/MM4 N_XI6/XI3/NET33_XI6/XI3/MM4_d N_XI6/XI3/NET34_XI6/XI3/MM4_g
+ N_VDD_XI6/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI3/MM10 N_XI6/XI3/NET35_XI6/XI3/MM10_d N_XI6/XI3/NET36_XI6/XI3/MM10_g
+ N_VDD_XI6/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI3/MM11 N_XI6/XI3/NET36_XI6/XI3/MM11_d N_XI6/XI3/NET35_XI6/XI3/MM11_g
+ N_VDD_XI6/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI4/MM2 N_XI6/XI4/NET34_XI6/XI4/MM2_d N_XI6/XI4/NET33_XI6/XI4/MM2_g
+ N_VSS_XI6/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM3 N_XI6/XI4/NET33_XI6/XI4/MM3_d N_WL<8>_XI6/XI4/MM3_g
+ N_BLN<11>_XI6/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM0 N_XI6/XI4/NET34_XI6/XI4/MM0_d N_WL<8>_XI6/XI4/MM0_g
+ N_BL<11>_XI6/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM1 N_XI6/XI4/NET33_XI6/XI4/MM1_d N_XI6/XI4/NET34_XI6/XI4/MM1_g
+ N_VSS_XI6/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM9 N_XI6/XI4/NET36_XI6/XI4/MM9_d N_WL<9>_XI6/XI4/MM9_g
+ N_BL<11>_XI6/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM6 N_XI6/XI4/NET35_XI6/XI4/MM6_d N_XI6/XI4/NET36_XI6/XI4/MM6_g
+ N_VSS_XI6/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM7 N_XI6/XI4/NET36_XI6/XI4/MM7_d N_XI6/XI4/NET35_XI6/XI4/MM7_g
+ N_VSS_XI6/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM8 N_XI6/XI4/NET35_XI6/XI4/MM8_d N_WL<9>_XI6/XI4/MM8_g
+ N_BLN<11>_XI6/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI4/MM5 N_XI6/XI4/NET34_XI6/XI4/MM5_d N_XI6/XI4/NET33_XI6/XI4/MM5_g
+ N_VDD_XI6/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI4/MM4 N_XI6/XI4/NET33_XI6/XI4/MM4_d N_XI6/XI4/NET34_XI6/XI4/MM4_g
+ N_VDD_XI6/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI4/MM10 N_XI6/XI4/NET35_XI6/XI4/MM10_d N_XI6/XI4/NET36_XI6/XI4/MM10_g
+ N_VDD_XI6/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI4/MM11 N_XI6/XI4/NET36_XI6/XI4/MM11_d N_XI6/XI4/NET35_XI6/XI4/MM11_g
+ N_VDD_XI6/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI5/MM2 N_XI6/XI5/NET34_XI6/XI5/MM2_d N_XI6/XI5/NET33_XI6/XI5/MM2_g
+ N_VSS_XI6/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM3 N_XI6/XI5/NET33_XI6/XI5/MM3_d N_WL<8>_XI6/XI5/MM3_g
+ N_BLN<10>_XI6/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM0 N_XI6/XI5/NET34_XI6/XI5/MM0_d N_WL<8>_XI6/XI5/MM0_g
+ N_BL<10>_XI6/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM1 N_XI6/XI5/NET33_XI6/XI5/MM1_d N_XI6/XI5/NET34_XI6/XI5/MM1_g
+ N_VSS_XI6/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM9 N_XI6/XI5/NET36_XI6/XI5/MM9_d N_WL<9>_XI6/XI5/MM9_g
+ N_BL<10>_XI6/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM6 N_XI6/XI5/NET35_XI6/XI5/MM6_d N_XI6/XI5/NET36_XI6/XI5/MM6_g
+ N_VSS_XI6/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM7 N_XI6/XI5/NET36_XI6/XI5/MM7_d N_XI6/XI5/NET35_XI6/XI5/MM7_g
+ N_VSS_XI6/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM8 N_XI6/XI5/NET35_XI6/XI5/MM8_d N_WL<9>_XI6/XI5/MM8_g
+ N_BLN<10>_XI6/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI5/MM5 N_XI6/XI5/NET34_XI6/XI5/MM5_d N_XI6/XI5/NET33_XI6/XI5/MM5_g
+ N_VDD_XI6/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI5/MM4 N_XI6/XI5/NET33_XI6/XI5/MM4_d N_XI6/XI5/NET34_XI6/XI5/MM4_g
+ N_VDD_XI6/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI5/MM10 N_XI6/XI5/NET35_XI6/XI5/MM10_d N_XI6/XI5/NET36_XI6/XI5/MM10_g
+ N_VDD_XI6/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI5/MM11 N_XI6/XI5/NET36_XI6/XI5/MM11_d N_XI6/XI5/NET35_XI6/XI5/MM11_g
+ N_VDD_XI6/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI6/MM2 N_XI6/XI6/NET34_XI6/XI6/MM2_d N_XI6/XI6/NET33_XI6/XI6/MM2_g
+ N_VSS_XI6/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM3 N_XI6/XI6/NET33_XI6/XI6/MM3_d N_WL<8>_XI6/XI6/MM3_g
+ N_BLN<9>_XI6/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM0 N_XI6/XI6/NET34_XI6/XI6/MM0_d N_WL<8>_XI6/XI6/MM0_g
+ N_BL<9>_XI6/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM1 N_XI6/XI6/NET33_XI6/XI6/MM1_d N_XI6/XI6/NET34_XI6/XI6/MM1_g
+ N_VSS_XI6/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM9 N_XI6/XI6/NET36_XI6/XI6/MM9_d N_WL<9>_XI6/XI6/MM9_g
+ N_BL<9>_XI6/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM6 N_XI6/XI6/NET35_XI6/XI6/MM6_d N_XI6/XI6/NET36_XI6/XI6/MM6_g
+ N_VSS_XI6/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM7 N_XI6/XI6/NET36_XI6/XI6/MM7_d N_XI6/XI6/NET35_XI6/XI6/MM7_g
+ N_VSS_XI6/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM8 N_XI6/XI6/NET35_XI6/XI6/MM8_d N_WL<9>_XI6/XI6/MM8_g
+ N_BLN<9>_XI6/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI6/MM5 N_XI6/XI6/NET34_XI6/XI6/MM5_d N_XI6/XI6/NET33_XI6/XI6/MM5_g
+ N_VDD_XI6/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI6/MM4 N_XI6/XI6/NET33_XI6/XI6/MM4_d N_XI6/XI6/NET34_XI6/XI6/MM4_g
+ N_VDD_XI6/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI6/MM10 N_XI6/XI6/NET35_XI6/XI6/MM10_d N_XI6/XI6/NET36_XI6/XI6/MM10_g
+ N_VDD_XI6/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI6/MM11 N_XI6/XI6/NET36_XI6/XI6/MM11_d N_XI6/XI6/NET35_XI6/XI6/MM11_g
+ N_VDD_XI6/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI7/MM2 N_XI6/XI7/NET34_XI6/XI7/MM2_d N_XI6/XI7/NET33_XI6/XI7/MM2_g
+ N_VSS_XI6/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM3 N_XI6/XI7/NET33_XI6/XI7/MM3_d N_WL<8>_XI6/XI7/MM3_g
+ N_BLN<8>_XI6/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM0 N_XI6/XI7/NET34_XI6/XI7/MM0_d N_WL<8>_XI6/XI7/MM0_g
+ N_BL<8>_XI6/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM1 N_XI6/XI7/NET33_XI6/XI7/MM1_d N_XI6/XI7/NET34_XI6/XI7/MM1_g
+ N_VSS_XI6/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM9 N_XI6/XI7/NET36_XI6/XI7/MM9_d N_WL<9>_XI6/XI7/MM9_g
+ N_BL<8>_XI6/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM6 N_XI6/XI7/NET35_XI6/XI7/MM6_d N_XI6/XI7/NET36_XI6/XI7/MM6_g
+ N_VSS_XI6/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM7 N_XI6/XI7/NET36_XI6/XI7/MM7_d N_XI6/XI7/NET35_XI6/XI7/MM7_g
+ N_VSS_XI6/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM8 N_XI6/XI7/NET35_XI6/XI7/MM8_d N_WL<9>_XI6/XI7/MM8_g
+ N_BLN<8>_XI6/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI7/MM5 N_XI6/XI7/NET34_XI6/XI7/MM5_d N_XI6/XI7/NET33_XI6/XI7/MM5_g
+ N_VDD_XI6/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI7/MM4 N_XI6/XI7/NET33_XI6/XI7/MM4_d N_XI6/XI7/NET34_XI6/XI7/MM4_g
+ N_VDD_XI6/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI7/MM10 N_XI6/XI7/NET35_XI6/XI7/MM10_d N_XI6/XI7/NET36_XI6/XI7/MM10_g
+ N_VDD_XI6/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI7/MM11 N_XI6/XI7/NET36_XI6/XI7/MM11_d N_XI6/XI7/NET35_XI6/XI7/MM11_g
+ N_VDD_XI6/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI8/MM2 N_XI6/XI8/NET34_XI6/XI8/MM2_d N_XI6/XI8/NET33_XI6/XI8/MM2_g
+ N_VSS_XI6/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM3 N_XI6/XI8/NET33_XI6/XI8/MM3_d N_WL<8>_XI6/XI8/MM3_g
+ N_BLN<7>_XI6/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM0 N_XI6/XI8/NET34_XI6/XI8/MM0_d N_WL<8>_XI6/XI8/MM0_g
+ N_BL<7>_XI6/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM1 N_XI6/XI8/NET33_XI6/XI8/MM1_d N_XI6/XI8/NET34_XI6/XI8/MM1_g
+ N_VSS_XI6/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM9 N_XI6/XI8/NET36_XI6/XI8/MM9_d N_WL<9>_XI6/XI8/MM9_g
+ N_BL<7>_XI6/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM6 N_XI6/XI8/NET35_XI6/XI8/MM6_d N_XI6/XI8/NET36_XI6/XI8/MM6_g
+ N_VSS_XI6/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM7 N_XI6/XI8/NET36_XI6/XI8/MM7_d N_XI6/XI8/NET35_XI6/XI8/MM7_g
+ N_VSS_XI6/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM8 N_XI6/XI8/NET35_XI6/XI8/MM8_d N_WL<9>_XI6/XI8/MM8_g
+ N_BLN<7>_XI6/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI8/MM5 N_XI6/XI8/NET34_XI6/XI8/MM5_d N_XI6/XI8/NET33_XI6/XI8/MM5_g
+ N_VDD_XI6/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI8/MM4 N_XI6/XI8/NET33_XI6/XI8/MM4_d N_XI6/XI8/NET34_XI6/XI8/MM4_g
+ N_VDD_XI6/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI8/MM10 N_XI6/XI8/NET35_XI6/XI8/MM10_d N_XI6/XI8/NET36_XI6/XI8/MM10_g
+ N_VDD_XI6/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI8/MM11 N_XI6/XI8/NET36_XI6/XI8/MM11_d N_XI6/XI8/NET35_XI6/XI8/MM11_g
+ N_VDD_XI6/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI9/MM2 N_XI6/XI9/NET34_XI6/XI9/MM2_d N_XI6/XI9/NET33_XI6/XI9/MM2_g
+ N_VSS_XI6/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM3 N_XI6/XI9/NET33_XI6/XI9/MM3_d N_WL<8>_XI6/XI9/MM3_g
+ N_BLN<6>_XI6/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM0 N_XI6/XI9/NET34_XI6/XI9/MM0_d N_WL<8>_XI6/XI9/MM0_g
+ N_BL<6>_XI6/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM1 N_XI6/XI9/NET33_XI6/XI9/MM1_d N_XI6/XI9/NET34_XI6/XI9/MM1_g
+ N_VSS_XI6/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM9 N_XI6/XI9/NET36_XI6/XI9/MM9_d N_WL<9>_XI6/XI9/MM9_g
+ N_BL<6>_XI6/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM6 N_XI6/XI9/NET35_XI6/XI9/MM6_d N_XI6/XI9/NET36_XI6/XI9/MM6_g
+ N_VSS_XI6/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM7 N_XI6/XI9/NET36_XI6/XI9/MM7_d N_XI6/XI9/NET35_XI6/XI9/MM7_g
+ N_VSS_XI6/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM8 N_XI6/XI9/NET35_XI6/XI9/MM8_d N_WL<9>_XI6/XI9/MM8_g
+ N_BLN<6>_XI6/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI9/MM5 N_XI6/XI9/NET34_XI6/XI9/MM5_d N_XI6/XI9/NET33_XI6/XI9/MM5_g
+ N_VDD_XI6/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI9/MM4 N_XI6/XI9/NET33_XI6/XI9/MM4_d N_XI6/XI9/NET34_XI6/XI9/MM4_g
+ N_VDD_XI6/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI9/MM10 N_XI6/XI9/NET35_XI6/XI9/MM10_d N_XI6/XI9/NET36_XI6/XI9/MM10_g
+ N_VDD_XI6/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI9/MM11 N_XI6/XI9/NET36_XI6/XI9/MM11_d N_XI6/XI9/NET35_XI6/XI9/MM11_g
+ N_VDD_XI6/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI10/MM2 N_XI6/XI10/NET34_XI6/XI10/MM2_d N_XI6/XI10/NET33_XI6/XI10/MM2_g
+ N_VSS_XI6/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI10/MM3 N_XI6/XI10/NET33_XI6/XI10/MM3_d N_WL<8>_XI6/XI10/MM3_g
+ N_BLN<5>_XI6/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI10/MM0 N_XI6/XI10/NET34_XI6/XI10/MM0_d N_WL<8>_XI6/XI10/MM0_g
+ N_BL<5>_XI6/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI10/MM1 N_XI6/XI10/NET33_XI6/XI10/MM1_d N_XI6/XI10/NET34_XI6/XI10/MM1_g
+ N_VSS_XI6/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI10/MM9 N_XI6/XI10/NET36_XI6/XI10/MM9_d N_WL<9>_XI6/XI10/MM9_g
+ N_BL<5>_XI6/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI10/MM6 N_XI6/XI10/NET35_XI6/XI10/MM6_d N_XI6/XI10/NET36_XI6/XI10/MM6_g
+ N_VSS_XI6/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI10/MM7 N_XI6/XI10/NET36_XI6/XI10/MM7_d N_XI6/XI10/NET35_XI6/XI10/MM7_g
+ N_VSS_XI6/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI10/MM8 N_XI6/XI10/NET35_XI6/XI10/MM8_d N_WL<9>_XI6/XI10/MM8_g
+ N_BLN<5>_XI6/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI10/MM5 N_XI6/XI10/NET34_XI6/XI10/MM5_d N_XI6/XI10/NET33_XI6/XI10/MM5_g
+ N_VDD_XI6/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI10/MM4 N_XI6/XI10/NET33_XI6/XI10/MM4_d N_XI6/XI10/NET34_XI6/XI10/MM4_g
+ N_VDD_XI6/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI10/MM10 N_XI6/XI10/NET35_XI6/XI10/MM10_d N_XI6/XI10/NET36_XI6/XI10/MM10_g
+ N_VDD_XI6/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI10/MM11 N_XI6/XI10/NET36_XI6/XI10/MM11_d N_XI6/XI10/NET35_XI6/XI10/MM11_g
+ N_VDD_XI6/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI11/MM2 N_XI6/XI11/NET34_XI6/XI11/MM2_d N_XI6/XI11/NET33_XI6/XI11/MM2_g
+ N_VSS_XI6/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI11/MM3 N_XI6/XI11/NET33_XI6/XI11/MM3_d N_WL<8>_XI6/XI11/MM3_g
+ N_BLN<4>_XI6/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI11/MM0 N_XI6/XI11/NET34_XI6/XI11/MM0_d N_WL<8>_XI6/XI11/MM0_g
+ N_BL<4>_XI6/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI11/MM1 N_XI6/XI11/NET33_XI6/XI11/MM1_d N_XI6/XI11/NET34_XI6/XI11/MM1_g
+ N_VSS_XI6/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI11/MM9 N_XI6/XI11/NET36_XI6/XI11/MM9_d N_WL<9>_XI6/XI11/MM9_g
+ N_BL<4>_XI6/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI11/MM6 N_XI6/XI11/NET35_XI6/XI11/MM6_d N_XI6/XI11/NET36_XI6/XI11/MM6_g
+ N_VSS_XI6/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI11/MM7 N_XI6/XI11/NET36_XI6/XI11/MM7_d N_XI6/XI11/NET35_XI6/XI11/MM7_g
+ N_VSS_XI6/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI11/MM8 N_XI6/XI11/NET35_XI6/XI11/MM8_d N_WL<9>_XI6/XI11/MM8_g
+ N_BLN<4>_XI6/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI11/MM5 N_XI6/XI11/NET34_XI6/XI11/MM5_d N_XI6/XI11/NET33_XI6/XI11/MM5_g
+ N_VDD_XI6/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI11/MM4 N_XI6/XI11/NET33_XI6/XI11/MM4_d N_XI6/XI11/NET34_XI6/XI11/MM4_g
+ N_VDD_XI6/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI11/MM10 N_XI6/XI11/NET35_XI6/XI11/MM10_d N_XI6/XI11/NET36_XI6/XI11/MM10_g
+ N_VDD_XI6/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI11/MM11 N_XI6/XI11/NET36_XI6/XI11/MM11_d N_XI6/XI11/NET35_XI6/XI11/MM11_g
+ N_VDD_XI6/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI12/MM2 N_XI6/XI12/NET34_XI6/XI12/MM2_d N_XI6/XI12/NET33_XI6/XI12/MM2_g
+ N_VSS_XI6/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI12/MM3 N_XI6/XI12/NET33_XI6/XI12/MM3_d N_WL<8>_XI6/XI12/MM3_g
+ N_BLN<3>_XI6/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI12/MM0 N_XI6/XI12/NET34_XI6/XI12/MM0_d N_WL<8>_XI6/XI12/MM0_g
+ N_BL<3>_XI6/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI12/MM1 N_XI6/XI12/NET33_XI6/XI12/MM1_d N_XI6/XI12/NET34_XI6/XI12/MM1_g
+ N_VSS_XI6/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI12/MM9 N_XI6/XI12/NET36_XI6/XI12/MM9_d N_WL<9>_XI6/XI12/MM9_g
+ N_BL<3>_XI6/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI12/MM6 N_XI6/XI12/NET35_XI6/XI12/MM6_d N_XI6/XI12/NET36_XI6/XI12/MM6_g
+ N_VSS_XI6/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI12/MM7 N_XI6/XI12/NET36_XI6/XI12/MM7_d N_XI6/XI12/NET35_XI6/XI12/MM7_g
+ N_VSS_XI6/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI12/MM8 N_XI6/XI12/NET35_XI6/XI12/MM8_d N_WL<9>_XI6/XI12/MM8_g
+ N_BLN<3>_XI6/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI12/MM5 N_XI6/XI12/NET34_XI6/XI12/MM5_d N_XI6/XI12/NET33_XI6/XI12/MM5_g
+ N_VDD_XI6/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI12/MM4 N_XI6/XI12/NET33_XI6/XI12/MM4_d N_XI6/XI12/NET34_XI6/XI12/MM4_g
+ N_VDD_XI6/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI12/MM10 N_XI6/XI12/NET35_XI6/XI12/MM10_d N_XI6/XI12/NET36_XI6/XI12/MM10_g
+ N_VDD_XI6/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI12/MM11 N_XI6/XI12/NET36_XI6/XI12/MM11_d N_XI6/XI12/NET35_XI6/XI12/MM11_g
+ N_VDD_XI6/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI13/MM2 N_XI6/XI13/NET34_XI6/XI13/MM2_d N_XI6/XI13/NET33_XI6/XI13/MM2_g
+ N_VSS_XI6/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI13/MM3 N_XI6/XI13/NET33_XI6/XI13/MM3_d N_WL<8>_XI6/XI13/MM3_g
+ N_BLN<2>_XI6/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI13/MM0 N_XI6/XI13/NET34_XI6/XI13/MM0_d N_WL<8>_XI6/XI13/MM0_g
+ N_BL<2>_XI6/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI13/MM1 N_XI6/XI13/NET33_XI6/XI13/MM1_d N_XI6/XI13/NET34_XI6/XI13/MM1_g
+ N_VSS_XI6/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI13/MM9 N_XI6/XI13/NET36_XI6/XI13/MM9_d N_WL<9>_XI6/XI13/MM9_g
+ N_BL<2>_XI6/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI13/MM6 N_XI6/XI13/NET35_XI6/XI13/MM6_d N_XI6/XI13/NET36_XI6/XI13/MM6_g
+ N_VSS_XI6/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI13/MM7 N_XI6/XI13/NET36_XI6/XI13/MM7_d N_XI6/XI13/NET35_XI6/XI13/MM7_g
+ N_VSS_XI6/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI13/MM8 N_XI6/XI13/NET35_XI6/XI13/MM8_d N_WL<9>_XI6/XI13/MM8_g
+ N_BLN<2>_XI6/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI13/MM5 N_XI6/XI13/NET34_XI6/XI13/MM5_d N_XI6/XI13/NET33_XI6/XI13/MM5_g
+ N_VDD_XI6/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI13/MM4 N_XI6/XI13/NET33_XI6/XI13/MM4_d N_XI6/XI13/NET34_XI6/XI13/MM4_g
+ N_VDD_XI6/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI13/MM10 N_XI6/XI13/NET35_XI6/XI13/MM10_d N_XI6/XI13/NET36_XI6/XI13/MM10_g
+ N_VDD_XI6/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI13/MM11 N_XI6/XI13/NET36_XI6/XI13/MM11_d N_XI6/XI13/NET35_XI6/XI13/MM11_g
+ N_VDD_XI6/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI14/MM2 N_XI6/XI14/NET34_XI6/XI14/MM2_d N_XI6/XI14/NET33_XI6/XI14/MM2_g
+ N_VSS_XI6/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI14/MM3 N_XI6/XI14/NET33_XI6/XI14/MM3_d N_WL<8>_XI6/XI14/MM3_g
+ N_BLN<1>_XI6/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI14/MM0 N_XI6/XI14/NET34_XI6/XI14/MM0_d N_WL<8>_XI6/XI14/MM0_g
+ N_BL<1>_XI6/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI14/MM1 N_XI6/XI14/NET33_XI6/XI14/MM1_d N_XI6/XI14/NET34_XI6/XI14/MM1_g
+ N_VSS_XI6/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI14/MM9 N_XI6/XI14/NET36_XI6/XI14/MM9_d N_WL<9>_XI6/XI14/MM9_g
+ N_BL<1>_XI6/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI14/MM6 N_XI6/XI14/NET35_XI6/XI14/MM6_d N_XI6/XI14/NET36_XI6/XI14/MM6_g
+ N_VSS_XI6/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI14/MM7 N_XI6/XI14/NET36_XI6/XI14/MM7_d N_XI6/XI14/NET35_XI6/XI14/MM7_g
+ N_VSS_XI6/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI14/MM8 N_XI6/XI14/NET35_XI6/XI14/MM8_d N_WL<9>_XI6/XI14/MM8_g
+ N_BLN<1>_XI6/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI14/MM5 N_XI6/XI14/NET34_XI6/XI14/MM5_d N_XI6/XI14/NET33_XI6/XI14/MM5_g
+ N_VDD_XI6/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI14/MM4 N_XI6/XI14/NET33_XI6/XI14/MM4_d N_XI6/XI14/NET34_XI6/XI14/MM4_g
+ N_VDD_XI6/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI14/MM10 N_XI6/XI14/NET35_XI6/XI14/MM10_d N_XI6/XI14/NET36_XI6/XI14/MM10_g
+ N_VDD_XI6/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI14/MM11 N_XI6/XI14/NET36_XI6/XI14/MM11_d N_XI6/XI14/NET35_XI6/XI14/MM11_g
+ N_VDD_XI6/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI15/MM2 N_XI6/XI15/NET34_XI6/XI15/MM2_d N_XI6/XI15/NET33_XI6/XI15/MM2_g
+ N_VSS_XI6/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI15/MM3 N_XI6/XI15/NET33_XI6/XI15/MM3_d N_WL<8>_XI6/XI15/MM3_g
+ N_BLN<0>_XI6/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI15/MM0 N_XI6/XI15/NET34_XI6/XI15/MM0_d N_WL<8>_XI6/XI15/MM0_g
+ N_BL<0>_XI6/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI15/MM1 N_XI6/XI15/NET33_XI6/XI15/MM1_d N_XI6/XI15/NET34_XI6/XI15/MM1_g
+ N_VSS_XI6/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI15/MM9 N_XI6/XI15/NET36_XI6/XI15/MM9_d N_WL<9>_XI6/XI15/MM9_g
+ N_BL<0>_XI6/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI15/MM6 N_XI6/XI15/NET35_XI6/XI15/MM6_d N_XI6/XI15/NET36_XI6/XI15/MM6_g
+ N_VSS_XI6/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI15/MM7 N_XI6/XI15/NET36_XI6/XI15/MM7_d N_XI6/XI15/NET35_XI6/XI15/MM7_g
+ N_VSS_XI6/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/XI15/MM8 N_XI6/XI15/NET35_XI6/XI15/MM8_d N_WL<9>_XI6/XI15/MM8_g
+ N_BLN<0>_XI6/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI6/XI15/MM5 N_XI6/XI15/NET34_XI6/XI15/MM5_d N_XI6/XI15/NET33_XI6/XI15/MM5_g
+ N_VDD_XI6/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI15/MM4 N_XI6/XI15/NET33_XI6/XI15/MM4_d N_XI6/XI15/NET34_XI6/XI15/MM4_g
+ N_VDD_XI6/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI15/MM10 N_XI6/XI15/NET35_XI6/XI15/MM10_d N_XI6/XI15/NET36_XI6/XI15/MM10_g
+ N_VDD_XI6/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/XI15/MM11 N_XI6/XI15/NET36_XI6/XI15/MM11_d N_XI6/XI15/NET35_XI6/XI15/MM11_g
+ N_VDD_XI6/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI0/MM2 N_XI7/XI0/NET34_XI7/XI0/MM2_d N_XI7/XI0/NET33_XI7/XI0/MM2_g
+ N_VSS_XI7/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM3 N_XI7/XI0/NET33_XI7/XI0/MM3_d N_WL<10>_XI7/XI0/MM3_g
+ N_BLN<15>_XI7/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM0 N_XI7/XI0/NET34_XI7/XI0/MM0_d N_WL<10>_XI7/XI0/MM0_g
+ N_BL<15>_XI7/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM1 N_XI7/XI0/NET33_XI7/XI0/MM1_d N_XI7/XI0/NET34_XI7/XI0/MM1_g
+ N_VSS_XI7/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM9 N_XI7/XI0/NET36_XI7/XI0/MM9_d N_WL<11>_XI7/XI0/MM9_g
+ N_BL<15>_XI7/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM6 N_XI7/XI0/NET35_XI7/XI0/MM6_d N_XI7/XI0/NET36_XI7/XI0/MM6_g
+ N_VSS_XI7/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM7 N_XI7/XI0/NET36_XI7/XI0/MM7_d N_XI7/XI0/NET35_XI7/XI0/MM7_g
+ N_VSS_XI7/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM8 N_XI7/XI0/NET35_XI7/XI0/MM8_d N_WL<11>_XI7/XI0/MM8_g
+ N_BLN<15>_XI7/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI0/MM5 N_XI7/XI0/NET34_XI7/XI0/MM5_d N_XI7/XI0/NET33_XI7/XI0/MM5_g
+ N_VDD_XI7/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI0/MM4 N_XI7/XI0/NET33_XI7/XI0/MM4_d N_XI7/XI0/NET34_XI7/XI0/MM4_g
+ N_VDD_XI7/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI0/MM10 N_XI7/XI0/NET35_XI7/XI0/MM10_d N_XI7/XI0/NET36_XI7/XI0/MM10_g
+ N_VDD_XI7/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI0/MM11 N_XI7/XI0/NET36_XI7/XI0/MM11_d N_XI7/XI0/NET35_XI7/XI0/MM11_g
+ N_VDD_XI7/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI1/MM2 N_XI7/XI1/NET34_XI7/XI1/MM2_d N_XI7/XI1/NET33_XI7/XI1/MM2_g
+ N_VSS_XI7/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM3 N_XI7/XI1/NET33_XI7/XI1/MM3_d N_WL<10>_XI7/XI1/MM3_g
+ N_BLN<14>_XI7/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM0 N_XI7/XI1/NET34_XI7/XI1/MM0_d N_WL<10>_XI7/XI1/MM0_g
+ N_BL<14>_XI7/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM1 N_XI7/XI1/NET33_XI7/XI1/MM1_d N_XI7/XI1/NET34_XI7/XI1/MM1_g
+ N_VSS_XI7/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM9 N_XI7/XI1/NET36_XI7/XI1/MM9_d N_WL<11>_XI7/XI1/MM9_g
+ N_BL<14>_XI7/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM6 N_XI7/XI1/NET35_XI7/XI1/MM6_d N_XI7/XI1/NET36_XI7/XI1/MM6_g
+ N_VSS_XI7/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM7 N_XI7/XI1/NET36_XI7/XI1/MM7_d N_XI7/XI1/NET35_XI7/XI1/MM7_g
+ N_VSS_XI7/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM8 N_XI7/XI1/NET35_XI7/XI1/MM8_d N_WL<11>_XI7/XI1/MM8_g
+ N_BLN<14>_XI7/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI1/MM5 N_XI7/XI1/NET34_XI7/XI1/MM5_d N_XI7/XI1/NET33_XI7/XI1/MM5_g
+ N_VDD_XI7/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI1/MM4 N_XI7/XI1/NET33_XI7/XI1/MM4_d N_XI7/XI1/NET34_XI7/XI1/MM4_g
+ N_VDD_XI7/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI1/MM10 N_XI7/XI1/NET35_XI7/XI1/MM10_d N_XI7/XI1/NET36_XI7/XI1/MM10_g
+ N_VDD_XI7/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI1/MM11 N_XI7/XI1/NET36_XI7/XI1/MM11_d N_XI7/XI1/NET35_XI7/XI1/MM11_g
+ N_VDD_XI7/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI2/MM2 N_XI7/XI2/NET34_XI7/XI2/MM2_d N_XI7/XI2/NET33_XI7/XI2/MM2_g
+ N_VSS_XI7/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM3 N_XI7/XI2/NET33_XI7/XI2/MM3_d N_WL<10>_XI7/XI2/MM3_g
+ N_BLN<13>_XI7/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM0 N_XI7/XI2/NET34_XI7/XI2/MM0_d N_WL<10>_XI7/XI2/MM0_g
+ N_BL<13>_XI7/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM1 N_XI7/XI2/NET33_XI7/XI2/MM1_d N_XI7/XI2/NET34_XI7/XI2/MM1_g
+ N_VSS_XI7/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM9 N_XI7/XI2/NET36_XI7/XI2/MM9_d N_WL<11>_XI7/XI2/MM9_g
+ N_BL<13>_XI7/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM6 N_XI7/XI2/NET35_XI7/XI2/MM6_d N_XI7/XI2/NET36_XI7/XI2/MM6_g
+ N_VSS_XI7/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM7 N_XI7/XI2/NET36_XI7/XI2/MM7_d N_XI7/XI2/NET35_XI7/XI2/MM7_g
+ N_VSS_XI7/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM8 N_XI7/XI2/NET35_XI7/XI2/MM8_d N_WL<11>_XI7/XI2/MM8_g
+ N_BLN<13>_XI7/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI2/MM5 N_XI7/XI2/NET34_XI7/XI2/MM5_d N_XI7/XI2/NET33_XI7/XI2/MM5_g
+ N_VDD_XI7/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI2/MM4 N_XI7/XI2/NET33_XI7/XI2/MM4_d N_XI7/XI2/NET34_XI7/XI2/MM4_g
+ N_VDD_XI7/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI2/MM10 N_XI7/XI2/NET35_XI7/XI2/MM10_d N_XI7/XI2/NET36_XI7/XI2/MM10_g
+ N_VDD_XI7/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI2/MM11 N_XI7/XI2/NET36_XI7/XI2/MM11_d N_XI7/XI2/NET35_XI7/XI2/MM11_g
+ N_VDD_XI7/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI3/MM2 N_XI7/XI3/NET34_XI7/XI3/MM2_d N_XI7/XI3/NET33_XI7/XI3/MM2_g
+ N_VSS_XI7/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM3 N_XI7/XI3/NET33_XI7/XI3/MM3_d N_WL<10>_XI7/XI3/MM3_g
+ N_BLN<12>_XI7/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM0 N_XI7/XI3/NET34_XI7/XI3/MM0_d N_WL<10>_XI7/XI3/MM0_g
+ N_BL<12>_XI7/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM1 N_XI7/XI3/NET33_XI7/XI3/MM1_d N_XI7/XI3/NET34_XI7/XI3/MM1_g
+ N_VSS_XI7/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM9 N_XI7/XI3/NET36_XI7/XI3/MM9_d N_WL<11>_XI7/XI3/MM9_g
+ N_BL<12>_XI7/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM6 N_XI7/XI3/NET35_XI7/XI3/MM6_d N_XI7/XI3/NET36_XI7/XI3/MM6_g
+ N_VSS_XI7/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM7 N_XI7/XI3/NET36_XI7/XI3/MM7_d N_XI7/XI3/NET35_XI7/XI3/MM7_g
+ N_VSS_XI7/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM8 N_XI7/XI3/NET35_XI7/XI3/MM8_d N_WL<11>_XI7/XI3/MM8_g
+ N_BLN<12>_XI7/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI3/MM5 N_XI7/XI3/NET34_XI7/XI3/MM5_d N_XI7/XI3/NET33_XI7/XI3/MM5_g
+ N_VDD_XI7/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI3/MM4 N_XI7/XI3/NET33_XI7/XI3/MM4_d N_XI7/XI3/NET34_XI7/XI3/MM4_g
+ N_VDD_XI7/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI3/MM10 N_XI7/XI3/NET35_XI7/XI3/MM10_d N_XI7/XI3/NET36_XI7/XI3/MM10_g
+ N_VDD_XI7/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI3/MM11 N_XI7/XI3/NET36_XI7/XI3/MM11_d N_XI7/XI3/NET35_XI7/XI3/MM11_g
+ N_VDD_XI7/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI4/MM2 N_XI7/XI4/NET34_XI7/XI4/MM2_d N_XI7/XI4/NET33_XI7/XI4/MM2_g
+ N_VSS_XI7/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM3 N_XI7/XI4/NET33_XI7/XI4/MM3_d N_WL<10>_XI7/XI4/MM3_g
+ N_BLN<11>_XI7/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM0 N_XI7/XI4/NET34_XI7/XI4/MM0_d N_WL<10>_XI7/XI4/MM0_g
+ N_BL<11>_XI7/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM1 N_XI7/XI4/NET33_XI7/XI4/MM1_d N_XI7/XI4/NET34_XI7/XI4/MM1_g
+ N_VSS_XI7/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM9 N_XI7/XI4/NET36_XI7/XI4/MM9_d N_WL<11>_XI7/XI4/MM9_g
+ N_BL<11>_XI7/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM6 N_XI7/XI4/NET35_XI7/XI4/MM6_d N_XI7/XI4/NET36_XI7/XI4/MM6_g
+ N_VSS_XI7/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM7 N_XI7/XI4/NET36_XI7/XI4/MM7_d N_XI7/XI4/NET35_XI7/XI4/MM7_g
+ N_VSS_XI7/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM8 N_XI7/XI4/NET35_XI7/XI4/MM8_d N_WL<11>_XI7/XI4/MM8_g
+ N_BLN<11>_XI7/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI4/MM5 N_XI7/XI4/NET34_XI7/XI4/MM5_d N_XI7/XI4/NET33_XI7/XI4/MM5_g
+ N_VDD_XI7/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI4/MM4 N_XI7/XI4/NET33_XI7/XI4/MM4_d N_XI7/XI4/NET34_XI7/XI4/MM4_g
+ N_VDD_XI7/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI4/MM10 N_XI7/XI4/NET35_XI7/XI4/MM10_d N_XI7/XI4/NET36_XI7/XI4/MM10_g
+ N_VDD_XI7/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI4/MM11 N_XI7/XI4/NET36_XI7/XI4/MM11_d N_XI7/XI4/NET35_XI7/XI4/MM11_g
+ N_VDD_XI7/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI5/MM2 N_XI7/XI5/NET34_XI7/XI5/MM2_d N_XI7/XI5/NET33_XI7/XI5/MM2_g
+ N_VSS_XI7/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM3 N_XI7/XI5/NET33_XI7/XI5/MM3_d N_WL<10>_XI7/XI5/MM3_g
+ N_BLN<10>_XI7/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM0 N_XI7/XI5/NET34_XI7/XI5/MM0_d N_WL<10>_XI7/XI5/MM0_g
+ N_BL<10>_XI7/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM1 N_XI7/XI5/NET33_XI7/XI5/MM1_d N_XI7/XI5/NET34_XI7/XI5/MM1_g
+ N_VSS_XI7/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM9 N_XI7/XI5/NET36_XI7/XI5/MM9_d N_WL<11>_XI7/XI5/MM9_g
+ N_BL<10>_XI7/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM6 N_XI7/XI5/NET35_XI7/XI5/MM6_d N_XI7/XI5/NET36_XI7/XI5/MM6_g
+ N_VSS_XI7/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM7 N_XI7/XI5/NET36_XI7/XI5/MM7_d N_XI7/XI5/NET35_XI7/XI5/MM7_g
+ N_VSS_XI7/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM8 N_XI7/XI5/NET35_XI7/XI5/MM8_d N_WL<11>_XI7/XI5/MM8_g
+ N_BLN<10>_XI7/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI5/MM5 N_XI7/XI5/NET34_XI7/XI5/MM5_d N_XI7/XI5/NET33_XI7/XI5/MM5_g
+ N_VDD_XI7/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI5/MM4 N_XI7/XI5/NET33_XI7/XI5/MM4_d N_XI7/XI5/NET34_XI7/XI5/MM4_g
+ N_VDD_XI7/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI5/MM10 N_XI7/XI5/NET35_XI7/XI5/MM10_d N_XI7/XI5/NET36_XI7/XI5/MM10_g
+ N_VDD_XI7/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI5/MM11 N_XI7/XI5/NET36_XI7/XI5/MM11_d N_XI7/XI5/NET35_XI7/XI5/MM11_g
+ N_VDD_XI7/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI6/MM2 N_XI7/XI6/NET34_XI7/XI6/MM2_d N_XI7/XI6/NET33_XI7/XI6/MM2_g
+ N_VSS_XI7/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM3 N_XI7/XI6/NET33_XI7/XI6/MM3_d N_WL<10>_XI7/XI6/MM3_g
+ N_BLN<9>_XI7/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM0 N_XI7/XI6/NET34_XI7/XI6/MM0_d N_WL<10>_XI7/XI6/MM0_g
+ N_BL<9>_XI7/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM1 N_XI7/XI6/NET33_XI7/XI6/MM1_d N_XI7/XI6/NET34_XI7/XI6/MM1_g
+ N_VSS_XI7/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM9 N_XI7/XI6/NET36_XI7/XI6/MM9_d N_WL<11>_XI7/XI6/MM9_g
+ N_BL<9>_XI7/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM6 N_XI7/XI6/NET35_XI7/XI6/MM6_d N_XI7/XI6/NET36_XI7/XI6/MM6_g
+ N_VSS_XI7/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM7 N_XI7/XI6/NET36_XI7/XI6/MM7_d N_XI7/XI6/NET35_XI7/XI6/MM7_g
+ N_VSS_XI7/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM8 N_XI7/XI6/NET35_XI7/XI6/MM8_d N_WL<11>_XI7/XI6/MM8_g
+ N_BLN<9>_XI7/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI6/MM5 N_XI7/XI6/NET34_XI7/XI6/MM5_d N_XI7/XI6/NET33_XI7/XI6/MM5_g
+ N_VDD_XI7/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI6/MM4 N_XI7/XI6/NET33_XI7/XI6/MM4_d N_XI7/XI6/NET34_XI7/XI6/MM4_g
+ N_VDD_XI7/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI6/MM10 N_XI7/XI6/NET35_XI7/XI6/MM10_d N_XI7/XI6/NET36_XI7/XI6/MM10_g
+ N_VDD_XI7/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI6/MM11 N_XI7/XI6/NET36_XI7/XI6/MM11_d N_XI7/XI6/NET35_XI7/XI6/MM11_g
+ N_VDD_XI7/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI7/MM2 N_XI7/XI7/NET34_XI7/XI7/MM2_d N_XI7/XI7/NET33_XI7/XI7/MM2_g
+ N_VSS_XI7/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM3 N_XI7/XI7/NET33_XI7/XI7/MM3_d N_WL<10>_XI7/XI7/MM3_g
+ N_BLN<8>_XI7/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM0 N_XI7/XI7/NET34_XI7/XI7/MM0_d N_WL<10>_XI7/XI7/MM0_g
+ N_BL<8>_XI7/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM1 N_XI7/XI7/NET33_XI7/XI7/MM1_d N_XI7/XI7/NET34_XI7/XI7/MM1_g
+ N_VSS_XI7/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM9 N_XI7/XI7/NET36_XI7/XI7/MM9_d N_WL<11>_XI7/XI7/MM9_g
+ N_BL<8>_XI7/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM6 N_XI7/XI7/NET35_XI7/XI7/MM6_d N_XI7/XI7/NET36_XI7/XI7/MM6_g
+ N_VSS_XI7/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM7 N_XI7/XI7/NET36_XI7/XI7/MM7_d N_XI7/XI7/NET35_XI7/XI7/MM7_g
+ N_VSS_XI7/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM8 N_XI7/XI7/NET35_XI7/XI7/MM8_d N_WL<11>_XI7/XI7/MM8_g
+ N_BLN<8>_XI7/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI7/MM5 N_XI7/XI7/NET34_XI7/XI7/MM5_d N_XI7/XI7/NET33_XI7/XI7/MM5_g
+ N_VDD_XI7/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI7/MM4 N_XI7/XI7/NET33_XI7/XI7/MM4_d N_XI7/XI7/NET34_XI7/XI7/MM4_g
+ N_VDD_XI7/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI7/MM10 N_XI7/XI7/NET35_XI7/XI7/MM10_d N_XI7/XI7/NET36_XI7/XI7/MM10_g
+ N_VDD_XI7/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI7/MM11 N_XI7/XI7/NET36_XI7/XI7/MM11_d N_XI7/XI7/NET35_XI7/XI7/MM11_g
+ N_VDD_XI7/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI8/MM2 N_XI7/XI8/NET34_XI7/XI8/MM2_d N_XI7/XI8/NET33_XI7/XI8/MM2_g
+ N_VSS_XI7/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM3 N_XI7/XI8/NET33_XI7/XI8/MM3_d N_WL<10>_XI7/XI8/MM3_g
+ N_BLN<7>_XI7/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM0 N_XI7/XI8/NET34_XI7/XI8/MM0_d N_WL<10>_XI7/XI8/MM0_g
+ N_BL<7>_XI7/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM1 N_XI7/XI8/NET33_XI7/XI8/MM1_d N_XI7/XI8/NET34_XI7/XI8/MM1_g
+ N_VSS_XI7/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM9 N_XI7/XI8/NET36_XI7/XI8/MM9_d N_WL<11>_XI7/XI8/MM9_g
+ N_BL<7>_XI7/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM6 N_XI7/XI8/NET35_XI7/XI8/MM6_d N_XI7/XI8/NET36_XI7/XI8/MM6_g
+ N_VSS_XI7/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM7 N_XI7/XI8/NET36_XI7/XI8/MM7_d N_XI7/XI8/NET35_XI7/XI8/MM7_g
+ N_VSS_XI7/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM8 N_XI7/XI8/NET35_XI7/XI8/MM8_d N_WL<11>_XI7/XI8/MM8_g
+ N_BLN<7>_XI7/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI8/MM5 N_XI7/XI8/NET34_XI7/XI8/MM5_d N_XI7/XI8/NET33_XI7/XI8/MM5_g
+ N_VDD_XI7/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI8/MM4 N_XI7/XI8/NET33_XI7/XI8/MM4_d N_XI7/XI8/NET34_XI7/XI8/MM4_g
+ N_VDD_XI7/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI8/MM10 N_XI7/XI8/NET35_XI7/XI8/MM10_d N_XI7/XI8/NET36_XI7/XI8/MM10_g
+ N_VDD_XI7/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI8/MM11 N_XI7/XI8/NET36_XI7/XI8/MM11_d N_XI7/XI8/NET35_XI7/XI8/MM11_g
+ N_VDD_XI7/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI9/MM2 N_XI7/XI9/NET34_XI7/XI9/MM2_d N_XI7/XI9/NET33_XI7/XI9/MM2_g
+ N_VSS_XI7/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM3 N_XI7/XI9/NET33_XI7/XI9/MM3_d N_WL<10>_XI7/XI9/MM3_g
+ N_BLN<6>_XI7/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM0 N_XI7/XI9/NET34_XI7/XI9/MM0_d N_WL<10>_XI7/XI9/MM0_g
+ N_BL<6>_XI7/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM1 N_XI7/XI9/NET33_XI7/XI9/MM1_d N_XI7/XI9/NET34_XI7/XI9/MM1_g
+ N_VSS_XI7/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM9 N_XI7/XI9/NET36_XI7/XI9/MM9_d N_WL<11>_XI7/XI9/MM9_g
+ N_BL<6>_XI7/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM6 N_XI7/XI9/NET35_XI7/XI9/MM6_d N_XI7/XI9/NET36_XI7/XI9/MM6_g
+ N_VSS_XI7/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM7 N_XI7/XI9/NET36_XI7/XI9/MM7_d N_XI7/XI9/NET35_XI7/XI9/MM7_g
+ N_VSS_XI7/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM8 N_XI7/XI9/NET35_XI7/XI9/MM8_d N_WL<11>_XI7/XI9/MM8_g
+ N_BLN<6>_XI7/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI9/MM5 N_XI7/XI9/NET34_XI7/XI9/MM5_d N_XI7/XI9/NET33_XI7/XI9/MM5_g
+ N_VDD_XI7/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI9/MM4 N_XI7/XI9/NET33_XI7/XI9/MM4_d N_XI7/XI9/NET34_XI7/XI9/MM4_g
+ N_VDD_XI7/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI9/MM10 N_XI7/XI9/NET35_XI7/XI9/MM10_d N_XI7/XI9/NET36_XI7/XI9/MM10_g
+ N_VDD_XI7/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI9/MM11 N_XI7/XI9/NET36_XI7/XI9/MM11_d N_XI7/XI9/NET35_XI7/XI9/MM11_g
+ N_VDD_XI7/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI10/MM2 N_XI7/XI10/NET34_XI7/XI10/MM2_d N_XI7/XI10/NET33_XI7/XI10/MM2_g
+ N_VSS_XI7/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI10/MM3 N_XI7/XI10/NET33_XI7/XI10/MM3_d N_WL<10>_XI7/XI10/MM3_g
+ N_BLN<5>_XI7/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI10/MM0 N_XI7/XI10/NET34_XI7/XI10/MM0_d N_WL<10>_XI7/XI10/MM0_g
+ N_BL<5>_XI7/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI10/MM1 N_XI7/XI10/NET33_XI7/XI10/MM1_d N_XI7/XI10/NET34_XI7/XI10/MM1_g
+ N_VSS_XI7/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI10/MM9 N_XI7/XI10/NET36_XI7/XI10/MM9_d N_WL<11>_XI7/XI10/MM9_g
+ N_BL<5>_XI7/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI10/MM6 N_XI7/XI10/NET35_XI7/XI10/MM6_d N_XI7/XI10/NET36_XI7/XI10/MM6_g
+ N_VSS_XI7/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI10/MM7 N_XI7/XI10/NET36_XI7/XI10/MM7_d N_XI7/XI10/NET35_XI7/XI10/MM7_g
+ N_VSS_XI7/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI10/MM8 N_XI7/XI10/NET35_XI7/XI10/MM8_d N_WL<11>_XI7/XI10/MM8_g
+ N_BLN<5>_XI7/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI10/MM5 N_XI7/XI10/NET34_XI7/XI10/MM5_d N_XI7/XI10/NET33_XI7/XI10/MM5_g
+ N_VDD_XI7/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI10/MM4 N_XI7/XI10/NET33_XI7/XI10/MM4_d N_XI7/XI10/NET34_XI7/XI10/MM4_g
+ N_VDD_XI7/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI10/MM10 N_XI7/XI10/NET35_XI7/XI10/MM10_d N_XI7/XI10/NET36_XI7/XI10/MM10_g
+ N_VDD_XI7/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI10/MM11 N_XI7/XI10/NET36_XI7/XI10/MM11_d N_XI7/XI10/NET35_XI7/XI10/MM11_g
+ N_VDD_XI7/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI11/MM2 N_XI7/XI11/NET34_XI7/XI11/MM2_d N_XI7/XI11/NET33_XI7/XI11/MM2_g
+ N_VSS_XI7/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI11/MM3 N_XI7/XI11/NET33_XI7/XI11/MM3_d N_WL<10>_XI7/XI11/MM3_g
+ N_BLN<4>_XI7/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI11/MM0 N_XI7/XI11/NET34_XI7/XI11/MM0_d N_WL<10>_XI7/XI11/MM0_g
+ N_BL<4>_XI7/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI11/MM1 N_XI7/XI11/NET33_XI7/XI11/MM1_d N_XI7/XI11/NET34_XI7/XI11/MM1_g
+ N_VSS_XI7/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI11/MM9 N_XI7/XI11/NET36_XI7/XI11/MM9_d N_WL<11>_XI7/XI11/MM9_g
+ N_BL<4>_XI7/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI11/MM6 N_XI7/XI11/NET35_XI7/XI11/MM6_d N_XI7/XI11/NET36_XI7/XI11/MM6_g
+ N_VSS_XI7/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI11/MM7 N_XI7/XI11/NET36_XI7/XI11/MM7_d N_XI7/XI11/NET35_XI7/XI11/MM7_g
+ N_VSS_XI7/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI11/MM8 N_XI7/XI11/NET35_XI7/XI11/MM8_d N_WL<11>_XI7/XI11/MM8_g
+ N_BLN<4>_XI7/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI11/MM5 N_XI7/XI11/NET34_XI7/XI11/MM5_d N_XI7/XI11/NET33_XI7/XI11/MM5_g
+ N_VDD_XI7/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI11/MM4 N_XI7/XI11/NET33_XI7/XI11/MM4_d N_XI7/XI11/NET34_XI7/XI11/MM4_g
+ N_VDD_XI7/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI11/MM10 N_XI7/XI11/NET35_XI7/XI11/MM10_d N_XI7/XI11/NET36_XI7/XI11/MM10_g
+ N_VDD_XI7/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI11/MM11 N_XI7/XI11/NET36_XI7/XI11/MM11_d N_XI7/XI11/NET35_XI7/XI11/MM11_g
+ N_VDD_XI7/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI12/MM2 N_XI7/XI12/NET34_XI7/XI12/MM2_d N_XI7/XI12/NET33_XI7/XI12/MM2_g
+ N_VSS_XI7/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI12/MM3 N_XI7/XI12/NET33_XI7/XI12/MM3_d N_WL<10>_XI7/XI12/MM3_g
+ N_BLN<3>_XI7/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI12/MM0 N_XI7/XI12/NET34_XI7/XI12/MM0_d N_WL<10>_XI7/XI12/MM0_g
+ N_BL<3>_XI7/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI12/MM1 N_XI7/XI12/NET33_XI7/XI12/MM1_d N_XI7/XI12/NET34_XI7/XI12/MM1_g
+ N_VSS_XI7/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI12/MM9 N_XI7/XI12/NET36_XI7/XI12/MM9_d N_WL<11>_XI7/XI12/MM9_g
+ N_BL<3>_XI7/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI12/MM6 N_XI7/XI12/NET35_XI7/XI12/MM6_d N_XI7/XI12/NET36_XI7/XI12/MM6_g
+ N_VSS_XI7/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI12/MM7 N_XI7/XI12/NET36_XI7/XI12/MM7_d N_XI7/XI12/NET35_XI7/XI12/MM7_g
+ N_VSS_XI7/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI12/MM8 N_XI7/XI12/NET35_XI7/XI12/MM8_d N_WL<11>_XI7/XI12/MM8_g
+ N_BLN<3>_XI7/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI12/MM5 N_XI7/XI12/NET34_XI7/XI12/MM5_d N_XI7/XI12/NET33_XI7/XI12/MM5_g
+ N_VDD_XI7/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI12/MM4 N_XI7/XI12/NET33_XI7/XI12/MM4_d N_XI7/XI12/NET34_XI7/XI12/MM4_g
+ N_VDD_XI7/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI12/MM10 N_XI7/XI12/NET35_XI7/XI12/MM10_d N_XI7/XI12/NET36_XI7/XI12/MM10_g
+ N_VDD_XI7/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI12/MM11 N_XI7/XI12/NET36_XI7/XI12/MM11_d N_XI7/XI12/NET35_XI7/XI12/MM11_g
+ N_VDD_XI7/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI13/MM2 N_XI7/XI13/NET34_XI7/XI13/MM2_d N_XI7/XI13/NET33_XI7/XI13/MM2_g
+ N_VSS_XI7/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI13/MM3 N_XI7/XI13/NET33_XI7/XI13/MM3_d N_WL<10>_XI7/XI13/MM3_g
+ N_BLN<2>_XI7/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI13/MM0 N_XI7/XI13/NET34_XI7/XI13/MM0_d N_WL<10>_XI7/XI13/MM0_g
+ N_BL<2>_XI7/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI13/MM1 N_XI7/XI13/NET33_XI7/XI13/MM1_d N_XI7/XI13/NET34_XI7/XI13/MM1_g
+ N_VSS_XI7/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI13/MM9 N_XI7/XI13/NET36_XI7/XI13/MM9_d N_WL<11>_XI7/XI13/MM9_g
+ N_BL<2>_XI7/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI13/MM6 N_XI7/XI13/NET35_XI7/XI13/MM6_d N_XI7/XI13/NET36_XI7/XI13/MM6_g
+ N_VSS_XI7/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI13/MM7 N_XI7/XI13/NET36_XI7/XI13/MM7_d N_XI7/XI13/NET35_XI7/XI13/MM7_g
+ N_VSS_XI7/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI13/MM8 N_XI7/XI13/NET35_XI7/XI13/MM8_d N_WL<11>_XI7/XI13/MM8_g
+ N_BLN<2>_XI7/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI13/MM5 N_XI7/XI13/NET34_XI7/XI13/MM5_d N_XI7/XI13/NET33_XI7/XI13/MM5_g
+ N_VDD_XI7/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI13/MM4 N_XI7/XI13/NET33_XI7/XI13/MM4_d N_XI7/XI13/NET34_XI7/XI13/MM4_g
+ N_VDD_XI7/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI13/MM10 N_XI7/XI13/NET35_XI7/XI13/MM10_d N_XI7/XI13/NET36_XI7/XI13/MM10_g
+ N_VDD_XI7/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI13/MM11 N_XI7/XI13/NET36_XI7/XI13/MM11_d N_XI7/XI13/NET35_XI7/XI13/MM11_g
+ N_VDD_XI7/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI14/MM2 N_XI7/XI14/NET34_XI7/XI14/MM2_d N_XI7/XI14/NET33_XI7/XI14/MM2_g
+ N_VSS_XI7/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI14/MM3 N_XI7/XI14/NET33_XI7/XI14/MM3_d N_WL<10>_XI7/XI14/MM3_g
+ N_BLN<1>_XI7/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI14/MM0 N_XI7/XI14/NET34_XI7/XI14/MM0_d N_WL<10>_XI7/XI14/MM0_g
+ N_BL<1>_XI7/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI14/MM1 N_XI7/XI14/NET33_XI7/XI14/MM1_d N_XI7/XI14/NET34_XI7/XI14/MM1_g
+ N_VSS_XI7/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI14/MM9 N_XI7/XI14/NET36_XI7/XI14/MM9_d N_WL<11>_XI7/XI14/MM9_g
+ N_BL<1>_XI7/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI14/MM6 N_XI7/XI14/NET35_XI7/XI14/MM6_d N_XI7/XI14/NET36_XI7/XI14/MM6_g
+ N_VSS_XI7/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI14/MM7 N_XI7/XI14/NET36_XI7/XI14/MM7_d N_XI7/XI14/NET35_XI7/XI14/MM7_g
+ N_VSS_XI7/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI14/MM8 N_XI7/XI14/NET35_XI7/XI14/MM8_d N_WL<11>_XI7/XI14/MM8_g
+ N_BLN<1>_XI7/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI14/MM5 N_XI7/XI14/NET34_XI7/XI14/MM5_d N_XI7/XI14/NET33_XI7/XI14/MM5_g
+ N_VDD_XI7/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI14/MM4 N_XI7/XI14/NET33_XI7/XI14/MM4_d N_XI7/XI14/NET34_XI7/XI14/MM4_g
+ N_VDD_XI7/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI14/MM10 N_XI7/XI14/NET35_XI7/XI14/MM10_d N_XI7/XI14/NET36_XI7/XI14/MM10_g
+ N_VDD_XI7/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI14/MM11 N_XI7/XI14/NET36_XI7/XI14/MM11_d N_XI7/XI14/NET35_XI7/XI14/MM11_g
+ N_VDD_XI7/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI15/MM2 N_XI7/XI15/NET34_XI7/XI15/MM2_d N_XI7/XI15/NET33_XI7/XI15/MM2_g
+ N_VSS_XI7/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI15/MM3 N_XI7/XI15/NET33_XI7/XI15/MM3_d N_WL<10>_XI7/XI15/MM3_g
+ N_BLN<0>_XI7/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI15/MM0 N_XI7/XI15/NET34_XI7/XI15/MM0_d N_WL<10>_XI7/XI15/MM0_g
+ N_BL<0>_XI7/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI15/MM1 N_XI7/XI15/NET33_XI7/XI15/MM1_d N_XI7/XI15/NET34_XI7/XI15/MM1_g
+ N_VSS_XI7/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI15/MM9 N_XI7/XI15/NET36_XI7/XI15/MM9_d N_WL<11>_XI7/XI15/MM9_g
+ N_BL<0>_XI7/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI15/MM6 N_XI7/XI15/NET35_XI7/XI15/MM6_d N_XI7/XI15/NET36_XI7/XI15/MM6_g
+ N_VSS_XI7/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI15/MM7 N_XI7/XI15/NET36_XI7/XI15/MM7_d N_XI7/XI15/NET35_XI7/XI15/MM7_g
+ N_VSS_XI7/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/XI15/MM8 N_XI7/XI15/NET35_XI7/XI15/MM8_d N_WL<11>_XI7/XI15/MM8_g
+ N_BLN<0>_XI7/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI7/XI15/MM5 N_XI7/XI15/NET34_XI7/XI15/MM5_d N_XI7/XI15/NET33_XI7/XI15/MM5_g
+ N_VDD_XI7/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI15/MM4 N_XI7/XI15/NET33_XI7/XI15/MM4_d N_XI7/XI15/NET34_XI7/XI15/MM4_g
+ N_VDD_XI7/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI15/MM10 N_XI7/XI15/NET35_XI7/XI15/MM10_d N_XI7/XI15/NET36_XI7/XI15/MM10_g
+ N_VDD_XI7/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/XI15/MM11 N_XI7/XI15/NET36_XI7/XI15/MM11_d N_XI7/XI15/NET35_XI7/XI15/MM11_g
+ N_VDD_XI7/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI0/MM2 N_XI8/XI0/NET34_XI8/XI0/MM2_d N_XI8/XI0/NET33_XI8/XI0/MM2_g
+ N_VSS_XI8/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM3 N_XI8/XI0/NET33_XI8/XI0/MM3_d N_WL<12>_XI8/XI0/MM3_g
+ N_BLN<15>_XI8/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM0 N_XI8/XI0/NET34_XI8/XI0/MM0_d N_WL<12>_XI8/XI0/MM0_g
+ N_BL<15>_XI8/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM1 N_XI8/XI0/NET33_XI8/XI0/MM1_d N_XI8/XI0/NET34_XI8/XI0/MM1_g
+ N_VSS_XI8/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM9 N_XI8/XI0/NET36_XI8/XI0/MM9_d N_WL<13>_XI8/XI0/MM9_g
+ N_BL<15>_XI8/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM6 N_XI8/XI0/NET35_XI8/XI0/MM6_d N_XI8/XI0/NET36_XI8/XI0/MM6_g
+ N_VSS_XI8/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM7 N_XI8/XI0/NET36_XI8/XI0/MM7_d N_XI8/XI0/NET35_XI8/XI0/MM7_g
+ N_VSS_XI8/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM8 N_XI8/XI0/NET35_XI8/XI0/MM8_d N_WL<13>_XI8/XI0/MM8_g
+ N_BLN<15>_XI8/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI0/MM5 N_XI8/XI0/NET34_XI8/XI0/MM5_d N_XI8/XI0/NET33_XI8/XI0/MM5_g
+ N_VDD_XI8/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI0/MM4 N_XI8/XI0/NET33_XI8/XI0/MM4_d N_XI8/XI0/NET34_XI8/XI0/MM4_g
+ N_VDD_XI8/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI0/MM10 N_XI8/XI0/NET35_XI8/XI0/MM10_d N_XI8/XI0/NET36_XI8/XI0/MM10_g
+ N_VDD_XI8/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI0/MM11 N_XI8/XI0/NET36_XI8/XI0/MM11_d N_XI8/XI0/NET35_XI8/XI0/MM11_g
+ N_VDD_XI8/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI1/MM2 N_XI8/XI1/NET34_XI8/XI1/MM2_d N_XI8/XI1/NET33_XI8/XI1/MM2_g
+ N_VSS_XI8/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM3 N_XI8/XI1/NET33_XI8/XI1/MM3_d N_WL<12>_XI8/XI1/MM3_g
+ N_BLN<14>_XI8/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM0 N_XI8/XI1/NET34_XI8/XI1/MM0_d N_WL<12>_XI8/XI1/MM0_g
+ N_BL<14>_XI8/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM1 N_XI8/XI1/NET33_XI8/XI1/MM1_d N_XI8/XI1/NET34_XI8/XI1/MM1_g
+ N_VSS_XI8/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM9 N_XI8/XI1/NET36_XI8/XI1/MM9_d N_WL<13>_XI8/XI1/MM9_g
+ N_BL<14>_XI8/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM6 N_XI8/XI1/NET35_XI8/XI1/MM6_d N_XI8/XI1/NET36_XI8/XI1/MM6_g
+ N_VSS_XI8/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM7 N_XI8/XI1/NET36_XI8/XI1/MM7_d N_XI8/XI1/NET35_XI8/XI1/MM7_g
+ N_VSS_XI8/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM8 N_XI8/XI1/NET35_XI8/XI1/MM8_d N_WL<13>_XI8/XI1/MM8_g
+ N_BLN<14>_XI8/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI1/MM5 N_XI8/XI1/NET34_XI8/XI1/MM5_d N_XI8/XI1/NET33_XI8/XI1/MM5_g
+ N_VDD_XI8/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI1/MM4 N_XI8/XI1/NET33_XI8/XI1/MM4_d N_XI8/XI1/NET34_XI8/XI1/MM4_g
+ N_VDD_XI8/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI1/MM10 N_XI8/XI1/NET35_XI8/XI1/MM10_d N_XI8/XI1/NET36_XI8/XI1/MM10_g
+ N_VDD_XI8/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI1/MM11 N_XI8/XI1/NET36_XI8/XI1/MM11_d N_XI8/XI1/NET35_XI8/XI1/MM11_g
+ N_VDD_XI8/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI2/MM2 N_XI8/XI2/NET34_XI8/XI2/MM2_d N_XI8/XI2/NET33_XI8/XI2/MM2_g
+ N_VSS_XI8/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM3 N_XI8/XI2/NET33_XI8/XI2/MM3_d N_WL<12>_XI8/XI2/MM3_g
+ N_BLN<13>_XI8/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM0 N_XI8/XI2/NET34_XI8/XI2/MM0_d N_WL<12>_XI8/XI2/MM0_g
+ N_BL<13>_XI8/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM1 N_XI8/XI2/NET33_XI8/XI2/MM1_d N_XI8/XI2/NET34_XI8/XI2/MM1_g
+ N_VSS_XI8/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM9 N_XI8/XI2/NET36_XI8/XI2/MM9_d N_WL<13>_XI8/XI2/MM9_g
+ N_BL<13>_XI8/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM6 N_XI8/XI2/NET35_XI8/XI2/MM6_d N_XI8/XI2/NET36_XI8/XI2/MM6_g
+ N_VSS_XI8/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM7 N_XI8/XI2/NET36_XI8/XI2/MM7_d N_XI8/XI2/NET35_XI8/XI2/MM7_g
+ N_VSS_XI8/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM8 N_XI8/XI2/NET35_XI8/XI2/MM8_d N_WL<13>_XI8/XI2/MM8_g
+ N_BLN<13>_XI8/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI2/MM5 N_XI8/XI2/NET34_XI8/XI2/MM5_d N_XI8/XI2/NET33_XI8/XI2/MM5_g
+ N_VDD_XI8/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI2/MM4 N_XI8/XI2/NET33_XI8/XI2/MM4_d N_XI8/XI2/NET34_XI8/XI2/MM4_g
+ N_VDD_XI8/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI2/MM10 N_XI8/XI2/NET35_XI8/XI2/MM10_d N_XI8/XI2/NET36_XI8/XI2/MM10_g
+ N_VDD_XI8/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI2/MM11 N_XI8/XI2/NET36_XI8/XI2/MM11_d N_XI8/XI2/NET35_XI8/XI2/MM11_g
+ N_VDD_XI8/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI3/MM2 N_XI8/XI3/NET34_XI8/XI3/MM2_d N_XI8/XI3/NET33_XI8/XI3/MM2_g
+ N_VSS_XI8/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM3 N_XI8/XI3/NET33_XI8/XI3/MM3_d N_WL<12>_XI8/XI3/MM3_g
+ N_BLN<12>_XI8/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM0 N_XI8/XI3/NET34_XI8/XI3/MM0_d N_WL<12>_XI8/XI3/MM0_g
+ N_BL<12>_XI8/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM1 N_XI8/XI3/NET33_XI8/XI3/MM1_d N_XI8/XI3/NET34_XI8/XI3/MM1_g
+ N_VSS_XI8/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM9 N_XI8/XI3/NET36_XI8/XI3/MM9_d N_WL<13>_XI8/XI3/MM9_g
+ N_BL<12>_XI8/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM6 N_XI8/XI3/NET35_XI8/XI3/MM6_d N_XI8/XI3/NET36_XI8/XI3/MM6_g
+ N_VSS_XI8/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM7 N_XI8/XI3/NET36_XI8/XI3/MM7_d N_XI8/XI3/NET35_XI8/XI3/MM7_g
+ N_VSS_XI8/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM8 N_XI8/XI3/NET35_XI8/XI3/MM8_d N_WL<13>_XI8/XI3/MM8_g
+ N_BLN<12>_XI8/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI3/MM5 N_XI8/XI3/NET34_XI8/XI3/MM5_d N_XI8/XI3/NET33_XI8/XI3/MM5_g
+ N_VDD_XI8/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI3/MM4 N_XI8/XI3/NET33_XI8/XI3/MM4_d N_XI8/XI3/NET34_XI8/XI3/MM4_g
+ N_VDD_XI8/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI3/MM10 N_XI8/XI3/NET35_XI8/XI3/MM10_d N_XI8/XI3/NET36_XI8/XI3/MM10_g
+ N_VDD_XI8/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI3/MM11 N_XI8/XI3/NET36_XI8/XI3/MM11_d N_XI8/XI3/NET35_XI8/XI3/MM11_g
+ N_VDD_XI8/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI4/MM2 N_XI8/XI4/NET34_XI8/XI4/MM2_d N_XI8/XI4/NET33_XI8/XI4/MM2_g
+ N_VSS_XI8/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM3 N_XI8/XI4/NET33_XI8/XI4/MM3_d N_WL<12>_XI8/XI4/MM3_g
+ N_BLN<11>_XI8/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM0 N_XI8/XI4/NET34_XI8/XI4/MM0_d N_WL<12>_XI8/XI4/MM0_g
+ N_BL<11>_XI8/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM1 N_XI8/XI4/NET33_XI8/XI4/MM1_d N_XI8/XI4/NET34_XI8/XI4/MM1_g
+ N_VSS_XI8/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM9 N_XI8/XI4/NET36_XI8/XI4/MM9_d N_WL<13>_XI8/XI4/MM9_g
+ N_BL<11>_XI8/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM6 N_XI8/XI4/NET35_XI8/XI4/MM6_d N_XI8/XI4/NET36_XI8/XI4/MM6_g
+ N_VSS_XI8/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM7 N_XI8/XI4/NET36_XI8/XI4/MM7_d N_XI8/XI4/NET35_XI8/XI4/MM7_g
+ N_VSS_XI8/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM8 N_XI8/XI4/NET35_XI8/XI4/MM8_d N_WL<13>_XI8/XI4/MM8_g
+ N_BLN<11>_XI8/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI4/MM5 N_XI8/XI4/NET34_XI8/XI4/MM5_d N_XI8/XI4/NET33_XI8/XI4/MM5_g
+ N_VDD_XI8/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI4/MM4 N_XI8/XI4/NET33_XI8/XI4/MM4_d N_XI8/XI4/NET34_XI8/XI4/MM4_g
+ N_VDD_XI8/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI4/MM10 N_XI8/XI4/NET35_XI8/XI4/MM10_d N_XI8/XI4/NET36_XI8/XI4/MM10_g
+ N_VDD_XI8/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI4/MM11 N_XI8/XI4/NET36_XI8/XI4/MM11_d N_XI8/XI4/NET35_XI8/XI4/MM11_g
+ N_VDD_XI8/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI5/MM2 N_XI8/XI5/NET34_XI8/XI5/MM2_d N_XI8/XI5/NET33_XI8/XI5/MM2_g
+ N_VSS_XI8/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM3 N_XI8/XI5/NET33_XI8/XI5/MM3_d N_WL<12>_XI8/XI5/MM3_g
+ N_BLN<10>_XI8/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM0 N_XI8/XI5/NET34_XI8/XI5/MM0_d N_WL<12>_XI8/XI5/MM0_g
+ N_BL<10>_XI8/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM1 N_XI8/XI5/NET33_XI8/XI5/MM1_d N_XI8/XI5/NET34_XI8/XI5/MM1_g
+ N_VSS_XI8/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM9 N_XI8/XI5/NET36_XI8/XI5/MM9_d N_WL<13>_XI8/XI5/MM9_g
+ N_BL<10>_XI8/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM6 N_XI8/XI5/NET35_XI8/XI5/MM6_d N_XI8/XI5/NET36_XI8/XI5/MM6_g
+ N_VSS_XI8/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM7 N_XI8/XI5/NET36_XI8/XI5/MM7_d N_XI8/XI5/NET35_XI8/XI5/MM7_g
+ N_VSS_XI8/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM8 N_XI8/XI5/NET35_XI8/XI5/MM8_d N_WL<13>_XI8/XI5/MM8_g
+ N_BLN<10>_XI8/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI5/MM5 N_XI8/XI5/NET34_XI8/XI5/MM5_d N_XI8/XI5/NET33_XI8/XI5/MM5_g
+ N_VDD_XI8/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI5/MM4 N_XI8/XI5/NET33_XI8/XI5/MM4_d N_XI8/XI5/NET34_XI8/XI5/MM4_g
+ N_VDD_XI8/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI5/MM10 N_XI8/XI5/NET35_XI8/XI5/MM10_d N_XI8/XI5/NET36_XI8/XI5/MM10_g
+ N_VDD_XI8/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI5/MM11 N_XI8/XI5/NET36_XI8/XI5/MM11_d N_XI8/XI5/NET35_XI8/XI5/MM11_g
+ N_VDD_XI8/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI6/MM2 N_XI8/XI6/NET34_XI8/XI6/MM2_d N_XI8/XI6/NET33_XI8/XI6/MM2_g
+ N_VSS_XI8/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM3 N_XI8/XI6/NET33_XI8/XI6/MM3_d N_WL<12>_XI8/XI6/MM3_g
+ N_BLN<9>_XI8/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM0 N_XI8/XI6/NET34_XI8/XI6/MM0_d N_WL<12>_XI8/XI6/MM0_g
+ N_BL<9>_XI8/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM1 N_XI8/XI6/NET33_XI8/XI6/MM1_d N_XI8/XI6/NET34_XI8/XI6/MM1_g
+ N_VSS_XI8/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM9 N_XI8/XI6/NET36_XI8/XI6/MM9_d N_WL<13>_XI8/XI6/MM9_g
+ N_BL<9>_XI8/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM6 N_XI8/XI6/NET35_XI8/XI6/MM6_d N_XI8/XI6/NET36_XI8/XI6/MM6_g
+ N_VSS_XI8/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM7 N_XI8/XI6/NET36_XI8/XI6/MM7_d N_XI8/XI6/NET35_XI8/XI6/MM7_g
+ N_VSS_XI8/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM8 N_XI8/XI6/NET35_XI8/XI6/MM8_d N_WL<13>_XI8/XI6/MM8_g
+ N_BLN<9>_XI8/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI6/MM5 N_XI8/XI6/NET34_XI8/XI6/MM5_d N_XI8/XI6/NET33_XI8/XI6/MM5_g
+ N_VDD_XI8/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI6/MM4 N_XI8/XI6/NET33_XI8/XI6/MM4_d N_XI8/XI6/NET34_XI8/XI6/MM4_g
+ N_VDD_XI8/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI6/MM10 N_XI8/XI6/NET35_XI8/XI6/MM10_d N_XI8/XI6/NET36_XI8/XI6/MM10_g
+ N_VDD_XI8/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI6/MM11 N_XI8/XI6/NET36_XI8/XI6/MM11_d N_XI8/XI6/NET35_XI8/XI6/MM11_g
+ N_VDD_XI8/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI7/MM2 N_XI8/XI7/NET34_XI8/XI7/MM2_d N_XI8/XI7/NET33_XI8/XI7/MM2_g
+ N_VSS_XI8/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM3 N_XI8/XI7/NET33_XI8/XI7/MM3_d N_WL<12>_XI8/XI7/MM3_g
+ N_BLN<8>_XI8/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM0 N_XI8/XI7/NET34_XI8/XI7/MM0_d N_WL<12>_XI8/XI7/MM0_g
+ N_BL<8>_XI8/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM1 N_XI8/XI7/NET33_XI8/XI7/MM1_d N_XI8/XI7/NET34_XI8/XI7/MM1_g
+ N_VSS_XI8/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM9 N_XI8/XI7/NET36_XI8/XI7/MM9_d N_WL<13>_XI8/XI7/MM9_g
+ N_BL<8>_XI8/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM6 N_XI8/XI7/NET35_XI8/XI7/MM6_d N_XI8/XI7/NET36_XI8/XI7/MM6_g
+ N_VSS_XI8/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM7 N_XI8/XI7/NET36_XI8/XI7/MM7_d N_XI8/XI7/NET35_XI8/XI7/MM7_g
+ N_VSS_XI8/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM8 N_XI8/XI7/NET35_XI8/XI7/MM8_d N_WL<13>_XI8/XI7/MM8_g
+ N_BLN<8>_XI8/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI7/MM5 N_XI8/XI7/NET34_XI8/XI7/MM5_d N_XI8/XI7/NET33_XI8/XI7/MM5_g
+ N_VDD_XI8/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI7/MM4 N_XI8/XI7/NET33_XI8/XI7/MM4_d N_XI8/XI7/NET34_XI8/XI7/MM4_g
+ N_VDD_XI8/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI7/MM10 N_XI8/XI7/NET35_XI8/XI7/MM10_d N_XI8/XI7/NET36_XI8/XI7/MM10_g
+ N_VDD_XI8/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI7/MM11 N_XI8/XI7/NET36_XI8/XI7/MM11_d N_XI8/XI7/NET35_XI8/XI7/MM11_g
+ N_VDD_XI8/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI8/MM2 N_XI8/XI8/NET34_XI8/XI8/MM2_d N_XI8/XI8/NET33_XI8/XI8/MM2_g
+ N_VSS_XI8/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM3 N_XI8/XI8/NET33_XI8/XI8/MM3_d N_WL<12>_XI8/XI8/MM3_g
+ N_BLN<7>_XI8/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM0 N_XI8/XI8/NET34_XI8/XI8/MM0_d N_WL<12>_XI8/XI8/MM0_g
+ N_BL<7>_XI8/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM1 N_XI8/XI8/NET33_XI8/XI8/MM1_d N_XI8/XI8/NET34_XI8/XI8/MM1_g
+ N_VSS_XI8/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM9 N_XI8/XI8/NET36_XI8/XI8/MM9_d N_WL<13>_XI8/XI8/MM9_g
+ N_BL<7>_XI8/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM6 N_XI8/XI8/NET35_XI8/XI8/MM6_d N_XI8/XI8/NET36_XI8/XI8/MM6_g
+ N_VSS_XI8/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM7 N_XI8/XI8/NET36_XI8/XI8/MM7_d N_XI8/XI8/NET35_XI8/XI8/MM7_g
+ N_VSS_XI8/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM8 N_XI8/XI8/NET35_XI8/XI8/MM8_d N_WL<13>_XI8/XI8/MM8_g
+ N_BLN<7>_XI8/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI8/MM5 N_XI8/XI8/NET34_XI8/XI8/MM5_d N_XI8/XI8/NET33_XI8/XI8/MM5_g
+ N_VDD_XI8/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI8/MM4 N_XI8/XI8/NET33_XI8/XI8/MM4_d N_XI8/XI8/NET34_XI8/XI8/MM4_g
+ N_VDD_XI8/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI8/MM10 N_XI8/XI8/NET35_XI8/XI8/MM10_d N_XI8/XI8/NET36_XI8/XI8/MM10_g
+ N_VDD_XI8/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI8/MM11 N_XI8/XI8/NET36_XI8/XI8/MM11_d N_XI8/XI8/NET35_XI8/XI8/MM11_g
+ N_VDD_XI8/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI9/MM2 N_XI8/XI9/NET34_XI8/XI9/MM2_d N_XI8/XI9/NET33_XI8/XI9/MM2_g
+ N_VSS_XI8/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM3 N_XI8/XI9/NET33_XI8/XI9/MM3_d N_WL<12>_XI8/XI9/MM3_g
+ N_BLN<6>_XI8/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM0 N_XI8/XI9/NET34_XI8/XI9/MM0_d N_WL<12>_XI8/XI9/MM0_g
+ N_BL<6>_XI8/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM1 N_XI8/XI9/NET33_XI8/XI9/MM1_d N_XI8/XI9/NET34_XI8/XI9/MM1_g
+ N_VSS_XI8/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM9 N_XI8/XI9/NET36_XI8/XI9/MM9_d N_WL<13>_XI8/XI9/MM9_g
+ N_BL<6>_XI8/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM6 N_XI8/XI9/NET35_XI8/XI9/MM6_d N_XI8/XI9/NET36_XI8/XI9/MM6_g
+ N_VSS_XI8/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM7 N_XI8/XI9/NET36_XI8/XI9/MM7_d N_XI8/XI9/NET35_XI8/XI9/MM7_g
+ N_VSS_XI8/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM8 N_XI8/XI9/NET35_XI8/XI9/MM8_d N_WL<13>_XI8/XI9/MM8_g
+ N_BLN<6>_XI8/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI9/MM5 N_XI8/XI9/NET34_XI8/XI9/MM5_d N_XI8/XI9/NET33_XI8/XI9/MM5_g
+ N_VDD_XI8/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI9/MM4 N_XI8/XI9/NET33_XI8/XI9/MM4_d N_XI8/XI9/NET34_XI8/XI9/MM4_g
+ N_VDD_XI8/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI9/MM10 N_XI8/XI9/NET35_XI8/XI9/MM10_d N_XI8/XI9/NET36_XI8/XI9/MM10_g
+ N_VDD_XI8/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI9/MM11 N_XI8/XI9/NET36_XI8/XI9/MM11_d N_XI8/XI9/NET35_XI8/XI9/MM11_g
+ N_VDD_XI8/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI10/MM2 N_XI8/XI10/NET34_XI8/XI10/MM2_d N_XI8/XI10/NET33_XI8/XI10/MM2_g
+ N_VSS_XI8/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI10/MM3 N_XI8/XI10/NET33_XI8/XI10/MM3_d N_WL<12>_XI8/XI10/MM3_g
+ N_BLN<5>_XI8/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI10/MM0 N_XI8/XI10/NET34_XI8/XI10/MM0_d N_WL<12>_XI8/XI10/MM0_g
+ N_BL<5>_XI8/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI10/MM1 N_XI8/XI10/NET33_XI8/XI10/MM1_d N_XI8/XI10/NET34_XI8/XI10/MM1_g
+ N_VSS_XI8/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI10/MM9 N_XI8/XI10/NET36_XI8/XI10/MM9_d N_WL<13>_XI8/XI10/MM9_g
+ N_BL<5>_XI8/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI10/MM6 N_XI8/XI10/NET35_XI8/XI10/MM6_d N_XI8/XI10/NET36_XI8/XI10/MM6_g
+ N_VSS_XI8/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI10/MM7 N_XI8/XI10/NET36_XI8/XI10/MM7_d N_XI8/XI10/NET35_XI8/XI10/MM7_g
+ N_VSS_XI8/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI10/MM8 N_XI8/XI10/NET35_XI8/XI10/MM8_d N_WL<13>_XI8/XI10/MM8_g
+ N_BLN<5>_XI8/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI10/MM5 N_XI8/XI10/NET34_XI8/XI10/MM5_d N_XI8/XI10/NET33_XI8/XI10/MM5_g
+ N_VDD_XI8/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI10/MM4 N_XI8/XI10/NET33_XI8/XI10/MM4_d N_XI8/XI10/NET34_XI8/XI10/MM4_g
+ N_VDD_XI8/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI10/MM10 N_XI8/XI10/NET35_XI8/XI10/MM10_d N_XI8/XI10/NET36_XI8/XI10/MM10_g
+ N_VDD_XI8/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI10/MM11 N_XI8/XI10/NET36_XI8/XI10/MM11_d N_XI8/XI10/NET35_XI8/XI10/MM11_g
+ N_VDD_XI8/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI11/MM2 N_XI8/XI11/NET34_XI8/XI11/MM2_d N_XI8/XI11/NET33_XI8/XI11/MM2_g
+ N_VSS_XI8/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI11/MM3 N_XI8/XI11/NET33_XI8/XI11/MM3_d N_WL<12>_XI8/XI11/MM3_g
+ N_BLN<4>_XI8/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI11/MM0 N_XI8/XI11/NET34_XI8/XI11/MM0_d N_WL<12>_XI8/XI11/MM0_g
+ N_BL<4>_XI8/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI11/MM1 N_XI8/XI11/NET33_XI8/XI11/MM1_d N_XI8/XI11/NET34_XI8/XI11/MM1_g
+ N_VSS_XI8/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI11/MM9 N_XI8/XI11/NET36_XI8/XI11/MM9_d N_WL<13>_XI8/XI11/MM9_g
+ N_BL<4>_XI8/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI11/MM6 N_XI8/XI11/NET35_XI8/XI11/MM6_d N_XI8/XI11/NET36_XI8/XI11/MM6_g
+ N_VSS_XI8/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI11/MM7 N_XI8/XI11/NET36_XI8/XI11/MM7_d N_XI8/XI11/NET35_XI8/XI11/MM7_g
+ N_VSS_XI8/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI11/MM8 N_XI8/XI11/NET35_XI8/XI11/MM8_d N_WL<13>_XI8/XI11/MM8_g
+ N_BLN<4>_XI8/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI11/MM5 N_XI8/XI11/NET34_XI8/XI11/MM5_d N_XI8/XI11/NET33_XI8/XI11/MM5_g
+ N_VDD_XI8/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI11/MM4 N_XI8/XI11/NET33_XI8/XI11/MM4_d N_XI8/XI11/NET34_XI8/XI11/MM4_g
+ N_VDD_XI8/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI11/MM10 N_XI8/XI11/NET35_XI8/XI11/MM10_d N_XI8/XI11/NET36_XI8/XI11/MM10_g
+ N_VDD_XI8/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI11/MM11 N_XI8/XI11/NET36_XI8/XI11/MM11_d N_XI8/XI11/NET35_XI8/XI11/MM11_g
+ N_VDD_XI8/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI12/MM2 N_XI8/XI12/NET34_XI8/XI12/MM2_d N_XI8/XI12/NET33_XI8/XI12/MM2_g
+ N_VSS_XI8/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI12/MM3 N_XI8/XI12/NET33_XI8/XI12/MM3_d N_WL<12>_XI8/XI12/MM3_g
+ N_BLN<3>_XI8/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI12/MM0 N_XI8/XI12/NET34_XI8/XI12/MM0_d N_WL<12>_XI8/XI12/MM0_g
+ N_BL<3>_XI8/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI12/MM1 N_XI8/XI12/NET33_XI8/XI12/MM1_d N_XI8/XI12/NET34_XI8/XI12/MM1_g
+ N_VSS_XI8/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI12/MM9 N_XI8/XI12/NET36_XI8/XI12/MM9_d N_WL<13>_XI8/XI12/MM9_g
+ N_BL<3>_XI8/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI12/MM6 N_XI8/XI12/NET35_XI8/XI12/MM6_d N_XI8/XI12/NET36_XI8/XI12/MM6_g
+ N_VSS_XI8/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI12/MM7 N_XI8/XI12/NET36_XI8/XI12/MM7_d N_XI8/XI12/NET35_XI8/XI12/MM7_g
+ N_VSS_XI8/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI12/MM8 N_XI8/XI12/NET35_XI8/XI12/MM8_d N_WL<13>_XI8/XI12/MM8_g
+ N_BLN<3>_XI8/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI12/MM5 N_XI8/XI12/NET34_XI8/XI12/MM5_d N_XI8/XI12/NET33_XI8/XI12/MM5_g
+ N_VDD_XI8/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI12/MM4 N_XI8/XI12/NET33_XI8/XI12/MM4_d N_XI8/XI12/NET34_XI8/XI12/MM4_g
+ N_VDD_XI8/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI12/MM10 N_XI8/XI12/NET35_XI8/XI12/MM10_d N_XI8/XI12/NET36_XI8/XI12/MM10_g
+ N_VDD_XI8/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI12/MM11 N_XI8/XI12/NET36_XI8/XI12/MM11_d N_XI8/XI12/NET35_XI8/XI12/MM11_g
+ N_VDD_XI8/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI13/MM2 N_XI8/XI13/NET34_XI8/XI13/MM2_d N_XI8/XI13/NET33_XI8/XI13/MM2_g
+ N_VSS_XI8/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI13/MM3 N_XI8/XI13/NET33_XI8/XI13/MM3_d N_WL<12>_XI8/XI13/MM3_g
+ N_BLN<2>_XI8/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI13/MM0 N_XI8/XI13/NET34_XI8/XI13/MM0_d N_WL<12>_XI8/XI13/MM0_g
+ N_BL<2>_XI8/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI13/MM1 N_XI8/XI13/NET33_XI8/XI13/MM1_d N_XI8/XI13/NET34_XI8/XI13/MM1_g
+ N_VSS_XI8/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI13/MM9 N_XI8/XI13/NET36_XI8/XI13/MM9_d N_WL<13>_XI8/XI13/MM9_g
+ N_BL<2>_XI8/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI13/MM6 N_XI8/XI13/NET35_XI8/XI13/MM6_d N_XI8/XI13/NET36_XI8/XI13/MM6_g
+ N_VSS_XI8/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI13/MM7 N_XI8/XI13/NET36_XI8/XI13/MM7_d N_XI8/XI13/NET35_XI8/XI13/MM7_g
+ N_VSS_XI8/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI13/MM8 N_XI8/XI13/NET35_XI8/XI13/MM8_d N_WL<13>_XI8/XI13/MM8_g
+ N_BLN<2>_XI8/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI13/MM5 N_XI8/XI13/NET34_XI8/XI13/MM5_d N_XI8/XI13/NET33_XI8/XI13/MM5_g
+ N_VDD_XI8/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI13/MM4 N_XI8/XI13/NET33_XI8/XI13/MM4_d N_XI8/XI13/NET34_XI8/XI13/MM4_g
+ N_VDD_XI8/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI13/MM10 N_XI8/XI13/NET35_XI8/XI13/MM10_d N_XI8/XI13/NET36_XI8/XI13/MM10_g
+ N_VDD_XI8/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI13/MM11 N_XI8/XI13/NET36_XI8/XI13/MM11_d N_XI8/XI13/NET35_XI8/XI13/MM11_g
+ N_VDD_XI8/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI14/MM2 N_XI8/XI14/NET34_XI8/XI14/MM2_d N_XI8/XI14/NET33_XI8/XI14/MM2_g
+ N_VSS_XI8/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI14/MM3 N_XI8/XI14/NET33_XI8/XI14/MM3_d N_WL<12>_XI8/XI14/MM3_g
+ N_BLN<1>_XI8/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI14/MM0 N_XI8/XI14/NET34_XI8/XI14/MM0_d N_WL<12>_XI8/XI14/MM0_g
+ N_BL<1>_XI8/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI14/MM1 N_XI8/XI14/NET33_XI8/XI14/MM1_d N_XI8/XI14/NET34_XI8/XI14/MM1_g
+ N_VSS_XI8/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI14/MM9 N_XI8/XI14/NET36_XI8/XI14/MM9_d N_WL<13>_XI8/XI14/MM9_g
+ N_BL<1>_XI8/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI14/MM6 N_XI8/XI14/NET35_XI8/XI14/MM6_d N_XI8/XI14/NET36_XI8/XI14/MM6_g
+ N_VSS_XI8/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI14/MM7 N_XI8/XI14/NET36_XI8/XI14/MM7_d N_XI8/XI14/NET35_XI8/XI14/MM7_g
+ N_VSS_XI8/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI14/MM8 N_XI8/XI14/NET35_XI8/XI14/MM8_d N_WL<13>_XI8/XI14/MM8_g
+ N_BLN<1>_XI8/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI14/MM5 N_XI8/XI14/NET34_XI8/XI14/MM5_d N_XI8/XI14/NET33_XI8/XI14/MM5_g
+ N_VDD_XI8/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI14/MM4 N_XI8/XI14/NET33_XI8/XI14/MM4_d N_XI8/XI14/NET34_XI8/XI14/MM4_g
+ N_VDD_XI8/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI14/MM10 N_XI8/XI14/NET35_XI8/XI14/MM10_d N_XI8/XI14/NET36_XI8/XI14/MM10_g
+ N_VDD_XI8/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI14/MM11 N_XI8/XI14/NET36_XI8/XI14/MM11_d N_XI8/XI14/NET35_XI8/XI14/MM11_g
+ N_VDD_XI8/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI15/MM2 N_XI8/XI15/NET34_XI8/XI15/MM2_d N_XI8/XI15/NET33_XI8/XI15/MM2_g
+ N_VSS_XI8/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI15/MM3 N_XI8/XI15/NET33_XI8/XI15/MM3_d N_WL<12>_XI8/XI15/MM3_g
+ N_BLN<0>_XI8/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI15/MM0 N_XI8/XI15/NET34_XI8/XI15/MM0_d N_WL<12>_XI8/XI15/MM0_g
+ N_BL<0>_XI8/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI15/MM1 N_XI8/XI15/NET33_XI8/XI15/MM1_d N_XI8/XI15/NET34_XI8/XI15/MM1_g
+ N_VSS_XI8/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI15/MM9 N_XI8/XI15/NET36_XI8/XI15/MM9_d N_WL<13>_XI8/XI15/MM9_g
+ N_BL<0>_XI8/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI15/MM6 N_XI8/XI15/NET35_XI8/XI15/MM6_d N_XI8/XI15/NET36_XI8/XI15/MM6_g
+ N_VSS_XI8/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI15/MM7 N_XI8/XI15/NET36_XI8/XI15/MM7_d N_XI8/XI15/NET35_XI8/XI15/MM7_g
+ N_VSS_XI8/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/XI15/MM8 N_XI8/XI15/NET35_XI8/XI15/MM8_d N_WL<13>_XI8/XI15/MM8_g
+ N_BLN<0>_XI8/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI8/XI15/MM5 N_XI8/XI15/NET34_XI8/XI15/MM5_d N_XI8/XI15/NET33_XI8/XI15/MM5_g
+ N_VDD_XI8/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI15/MM4 N_XI8/XI15/NET33_XI8/XI15/MM4_d N_XI8/XI15/NET34_XI8/XI15/MM4_g
+ N_VDD_XI8/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI15/MM10 N_XI8/XI15/NET35_XI8/XI15/MM10_d N_XI8/XI15/NET36_XI8/XI15/MM10_g
+ N_VDD_XI8/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/XI15/MM11 N_XI8/XI15/NET36_XI8/XI15/MM11_d N_XI8/XI15/NET35_XI8/XI15/MM11_g
+ N_VDD_XI8/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI0/MM2 N_XI9/XI0/NET34_XI9/XI0/MM2_d N_XI9/XI0/NET33_XI9/XI0/MM2_g
+ N_VSS_XI9/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM3 N_XI9/XI0/NET33_XI9/XI0/MM3_d N_WL<14>_XI9/XI0/MM3_g
+ N_BLN<15>_XI9/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM0 N_XI9/XI0/NET34_XI9/XI0/MM0_d N_WL<14>_XI9/XI0/MM0_g
+ N_BL<15>_XI9/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM1 N_XI9/XI0/NET33_XI9/XI0/MM1_d N_XI9/XI0/NET34_XI9/XI0/MM1_g
+ N_VSS_XI9/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM9 N_XI9/XI0/NET36_XI9/XI0/MM9_d N_WL<15>_XI9/XI0/MM9_g
+ N_BL<15>_XI9/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM6 N_XI9/XI0/NET35_XI9/XI0/MM6_d N_XI9/XI0/NET36_XI9/XI0/MM6_g
+ N_VSS_XI9/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM7 N_XI9/XI0/NET36_XI9/XI0/MM7_d N_XI9/XI0/NET35_XI9/XI0/MM7_g
+ N_VSS_XI9/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM8 N_XI9/XI0/NET35_XI9/XI0/MM8_d N_WL<15>_XI9/XI0/MM8_g
+ N_BLN<15>_XI9/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI0/MM5 N_XI9/XI0/NET34_XI9/XI0/MM5_d N_XI9/XI0/NET33_XI9/XI0/MM5_g
+ N_VDD_XI9/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI0/MM4 N_XI9/XI0/NET33_XI9/XI0/MM4_d N_XI9/XI0/NET34_XI9/XI0/MM4_g
+ N_VDD_XI9/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI0/MM10 N_XI9/XI0/NET35_XI9/XI0/MM10_d N_XI9/XI0/NET36_XI9/XI0/MM10_g
+ N_VDD_XI9/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI0/MM11 N_XI9/XI0/NET36_XI9/XI0/MM11_d N_XI9/XI0/NET35_XI9/XI0/MM11_g
+ N_VDD_XI9/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI1/MM2 N_XI9/XI1/NET34_XI9/XI1/MM2_d N_XI9/XI1/NET33_XI9/XI1/MM2_g
+ N_VSS_XI9/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM3 N_XI9/XI1/NET33_XI9/XI1/MM3_d N_WL<14>_XI9/XI1/MM3_g
+ N_BLN<14>_XI9/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM0 N_XI9/XI1/NET34_XI9/XI1/MM0_d N_WL<14>_XI9/XI1/MM0_g
+ N_BL<14>_XI9/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM1 N_XI9/XI1/NET33_XI9/XI1/MM1_d N_XI9/XI1/NET34_XI9/XI1/MM1_g
+ N_VSS_XI9/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM9 N_XI9/XI1/NET36_XI9/XI1/MM9_d N_WL<15>_XI9/XI1/MM9_g
+ N_BL<14>_XI9/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM6 N_XI9/XI1/NET35_XI9/XI1/MM6_d N_XI9/XI1/NET36_XI9/XI1/MM6_g
+ N_VSS_XI9/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM7 N_XI9/XI1/NET36_XI9/XI1/MM7_d N_XI9/XI1/NET35_XI9/XI1/MM7_g
+ N_VSS_XI9/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM8 N_XI9/XI1/NET35_XI9/XI1/MM8_d N_WL<15>_XI9/XI1/MM8_g
+ N_BLN<14>_XI9/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI1/MM5 N_XI9/XI1/NET34_XI9/XI1/MM5_d N_XI9/XI1/NET33_XI9/XI1/MM5_g
+ N_VDD_XI9/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI1/MM4 N_XI9/XI1/NET33_XI9/XI1/MM4_d N_XI9/XI1/NET34_XI9/XI1/MM4_g
+ N_VDD_XI9/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI1/MM10 N_XI9/XI1/NET35_XI9/XI1/MM10_d N_XI9/XI1/NET36_XI9/XI1/MM10_g
+ N_VDD_XI9/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI1/MM11 N_XI9/XI1/NET36_XI9/XI1/MM11_d N_XI9/XI1/NET35_XI9/XI1/MM11_g
+ N_VDD_XI9/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI2/MM2 N_XI9/XI2/NET34_XI9/XI2/MM2_d N_XI9/XI2/NET33_XI9/XI2/MM2_g
+ N_VSS_XI9/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM3 N_XI9/XI2/NET33_XI9/XI2/MM3_d N_WL<14>_XI9/XI2/MM3_g
+ N_BLN<13>_XI9/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM0 N_XI9/XI2/NET34_XI9/XI2/MM0_d N_WL<14>_XI9/XI2/MM0_g
+ N_BL<13>_XI9/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM1 N_XI9/XI2/NET33_XI9/XI2/MM1_d N_XI9/XI2/NET34_XI9/XI2/MM1_g
+ N_VSS_XI9/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM9 N_XI9/XI2/NET36_XI9/XI2/MM9_d N_WL<15>_XI9/XI2/MM9_g
+ N_BL<13>_XI9/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM6 N_XI9/XI2/NET35_XI9/XI2/MM6_d N_XI9/XI2/NET36_XI9/XI2/MM6_g
+ N_VSS_XI9/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM7 N_XI9/XI2/NET36_XI9/XI2/MM7_d N_XI9/XI2/NET35_XI9/XI2/MM7_g
+ N_VSS_XI9/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM8 N_XI9/XI2/NET35_XI9/XI2/MM8_d N_WL<15>_XI9/XI2/MM8_g
+ N_BLN<13>_XI9/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI2/MM5 N_XI9/XI2/NET34_XI9/XI2/MM5_d N_XI9/XI2/NET33_XI9/XI2/MM5_g
+ N_VDD_XI9/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI2/MM4 N_XI9/XI2/NET33_XI9/XI2/MM4_d N_XI9/XI2/NET34_XI9/XI2/MM4_g
+ N_VDD_XI9/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI2/MM10 N_XI9/XI2/NET35_XI9/XI2/MM10_d N_XI9/XI2/NET36_XI9/XI2/MM10_g
+ N_VDD_XI9/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI2/MM11 N_XI9/XI2/NET36_XI9/XI2/MM11_d N_XI9/XI2/NET35_XI9/XI2/MM11_g
+ N_VDD_XI9/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI3/MM2 N_XI9/XI3/NET34_XI9/XI3/MM2_d N_XI9/XI3/NET33_XI9/XI3/MM2_g
+ N_VSS_XI9/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM3 N_XI9/XI3/NET33_XI9/XI3/MM3_d N_WL<14>_XI9/XI3/MM3_g
+ N_BLN<12>_XI9/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM0 N_XI9/XI3/NET34_XI9/XI3/MM0_d N_WL<14>_XI9/XI3/MM0_g
+ N_BL<12>_XI9/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM1 N_XI9/XI3/NET33_XI9/XI3/MM1_d N_XI9/XI3/NET34_XI9/XI3/MM1_g
+ N_VSS_XI9/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM9 N_XI9/XI3/NET36_XI9/XI3/MM9_d N_WL<15>_XI9/XI3/MM9_g
+ N_BL<12>_XI9/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM6 N_XI9/XI3/NET35_XI9/XI3/MM6_d N_XI9/XI3/NET36_XI9/XI3/MM6_g
+ N_VSS_XI9/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM7 N_XI9/XI3/NET36_XI9/XI3/MM7_d N_XI9/XI3/NET35_XI9/XI3/MM7_g
+ N_VSS_XI9/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM8 N_XI9/XI3/NET35_XI9/XI3/MM8_d N_WL<15>_XI9/XI3/MM8_g
+ N_BLN<12>_XI9/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI3/MM5 N_XI9/XI3/NET34_XI9/XI3/MM5_d N_XI9/XI3/NET33_XI9/XI3/MM5_g
+ N_VDD_XI9/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI3/MM4 N_XI9/XI3/NET33_XI9/XI3/MM4_d N_XI9/XI3/NET34_XI9/XI3/MM4_g
+ N_VDD_XI9/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI3/MM10 N_XI9/XI3/NET35_XI9/XI3/MM10_d N_XI9/XI3/NET36_XI9/XI3/MM10_g
+ N_VDD_XI9/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI3/MM11 N_XI9/XI3/NET36_XI9/XI3/MM11_d N_XI9/XI3/NET35_XI9/XI3/MM11_g
+ N_VDD_XI9/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI4/MM2 N_XI9/XI4/NET34_XI9/XI4/MM2_d N_XI9/XI4/NET33_XI9/XI4/MM2_g
+ N_VSS_XI9/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM3 N_XI9/XI4/NET33_XI9/XI4/MM3_d N_WL<14>_XI9/XI4/MM3_g
+ N_BLN<11>_XI9/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM0 N_XI9/XI4/NET34_XI9/XI4/MM0_d N_WL<14>_XI9/XI4/MM0_g
+ N_BL<11>_XI9/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM1 N_XI9/XI4/NET33_XI9/XI4/MM1_d N_XI9/XI4/NET34_XI9/XI4/MM1_g
+ N_VSS_XI9/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM9 N_XI9/XI4/NET36_XI9/XI4/MM9_d N_WL<15>_XI9/XI4/MM9_g
+ N_BL<11>_XI9/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM6 N_XI9/XI4/NET35_XI9/XI4/MM6_d N_XI9/XI4/NET36_XI9/XI4/MM6_g
+ N_VSS_XI9/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM7 N_XI9/XI4/NET36_XI9/XI4/MM7_d N_XI9/XI4/NET35_XI9/XI4/MM7_g
+ N_VSS_XI9/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM8 N_XI9/XI4/NET35_XI9/XI4/MM8_d N_WL<15>_XI9/XI4/MM8_g
+ N_BLN<11>_XI9/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI4/MM5 N_XI9/XI4/NET34_XI9/XI4/MM5_d N_XI9/XI4/NET33_XI9/XI4/MM5_g
+ N_VDD_XI9/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI4/MM4 N_XI9/XI4/NET33_XI9/XI4/MM4_d N_XI9/XI4/NET34_XI9/XI4/MM4_g
+ N_VDD_XI9/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI4/MM10 N_XI9/XI4/NET35_XI9/XI4/MM10_d N_XI9/XI4/NET36_XI9/XI4/MM10_g
+ N_VDD_XI9/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI4/MM11 N_XI9/XI4/NET36_XI9/XI4/MM11_d N_XI9/XI4/NET35_XI9/XI4/MM11_g
+ N_VDD_XI9/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI5/MM2 N_XI9/XI5/NET34_XI9/XI5/MM2_d N_XI9/XI5/NET33_XI9/XI5/MM2_g
+ N_VSS_XI9/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM3 N_XI9/XI5/NET33_XI9/XI5/MM3_d N_WL<14>_XI9/XI5/MM3_g
+ N_BLN<10>_XI9/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM0 N_XI9/XI5/NET34_XI9/XI5/MM0_d N_WL<14>_XI9/XI5/MM0_g
+ N_BL<10>_XI9/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM1 N_XI9/XI5/NET33_XI9/XI5/MM1_d N_XI9/XI5/NET34_XI9/XI5/MM1_g
+ N_VSS_XI9/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM9 N_XI9/XI5/NET36_XI9/XI5/MM9_d N_WL<15>_XI9/XI5/MM9_g
+ N_BL<10>_XI9/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM6 N_XI9/XI5/NET35_XI9/XI5/MM6_d N_XI9/XI5/NET36_XI9/XI5/MM6_g
+ N_VSS_XI9/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM7 N_XI9/XI5/NET36_XI9/XI5/MM7_d N_XI9/XI5/NET35_XI9/XI5/MM7_g
+ N_VSS_XI9/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM8 N_XI9/XI5/NET35_XI9/XI5/MM8_d N_WL<15>_XI9/XI5/MM8_g
+ N_BLN<10>_XI9/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI5/MM5 N_XI9/XI5/NET34_XI9/XI5/MM5_d N_XI9/XI5/NET33_XI9/XI5/MM5_g
+ N_VDD_XI9/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI5/MM4 N_XI9/XI5/NET33_XI9/XI5/MM4_d N_XI9/XI5/NET34_XI9/XI5/MM4_g
+ N_VDD_XI9/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI5/MM10 N_XI9/XI5/NET35_XI9/XI5/MM10_d N_XI9/XI5/NET36_XI9/XI5/MM10_g
+ N_VDD_XI9/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI5/MM11 N_XI9/XI5/NET36_XI9/XI5/MM11_d N_XI9/XI5/NET35_XI9/XI5/MM11_g
+ N_VDD_XI9/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI6/MM2 N_XI9/XI6/NET34_XI9/XI6/MM2_d N_XI9/XI6/NET33_XI9/XI6/MM2_g
+ N_VSS_XI9/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM3 N_XI9/XI6/NET33_XI9/XI6/MM3_d N_WL<14>_XI9/XI6/MM3_g
+ N_BLN<9>_XI9/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM0 N_XI9/XI6/NET34_XI9/XI6/MM0_d N_WL<14>_XI9/XI6/MM0_g
+ N_BL<9>_XI9/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM1 N_XI9/XI6/NET33_XI9/XI6/MM1_d N_XI9/XI6/NET34_XI9/XI6/MM1_g
+ N_VSS_XI9/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM9 N_XI9/XI6/NET36_XI9/XI6/MM9_d N_WL<15>_XI9/XI6/MM9_g
+ N_BL<9>_XI9/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM6 N_XI9/XI6/NET35_XI9/XI6/MM6_d N_XI9/XI6/NET36_XI9/XI6/MM6_g
+ N_VSS_XI9/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM7 N_XI9/XI6/NET36_XI9/XI6/MM7_d N_XI9/XI6/NET35_XI9/XI6/MM7_g
+ N_VSS_XI9/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM8 N_XI9/XI6/NET35_XI9/XI6/MM8_d N_WL<15>_XI9/XI6/MM8_g
+ N_BLN<9>_XI9/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI6/MM5 N_XI9/XI6/NET34_XI9/XI6/MM5_d N_XI9/XI6/NET33_XI9/XI6/MM5_g
+ N_VDD_XI9/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI6/MM4 N_XI9/XI6/NET33_XI9/XI6/MM4_d N_XI9/XI6/NET34_XI9/XI6/MM4_g
+ N_VDD_XI9/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI6/MM10 N_XI9/XI6/NET35_XI9/XI6/MM10_d N_XI9/XI6/NET36_XI9/XI6/MM10_g
+ N_VDD_XI9/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI6/MM11 N_XI9/XI6/NET36_XI9/XI6/MM11_d N_XI9/XI6/NET35_XI9/XI6/MM11_g
+ N_VDD_XI9/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI7/MM2 N_XI9/XI7/NET34_XI9/XI7/MM2_d N_XI9/XI7/NET33_XI9/XI7/MM2_g
+ N_VSS_XI9/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM3 N_XI9/XI7/NET33_XI9/XI7/MM3_d N_WL<14>_XI9/XI7/MM3_g
+ N_BLN<8>_XI9/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM0 N_XI9/XI7/NET34_XI9/XI7/MM0_d N_WL<14>_XI9/XI7/MM0_g
+ N_BL<8>_XI9/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM1 N_XI9/XI7/NET33_XI9/XI7/MM1_d N_XI9/XI7/NET34_XI9/XI7/MM1_g
+ N_VSS_XI9/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM9 N_XI9/XI7/NET36_XI9/XI7/MM9_d N_WL<15>_XI9/XI7/MM9_g
+ N_BL<8>_XI9/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM6 N_XI9/XI7/NET35_XI9/XI7/MM6_d N_XI9/XI7/NET36_XI9/XI7/MM6_g
+ N_VSS_XI9/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM7 N_XI9/XI7/NET36_XI9/XI7/MM7_d N_XI9/XI7/NET35_XI9/XI7/MM7_g
+ N_VSS_XI9/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM8 N_XI9/XI7/NET35_XI9/XI7/MM8_d N_WL<15>_XI9/XI7/MM8_g
+ N_BLN<8>_XI9/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI7/MM5 N_XI9/XI7/NET34_XI9/XI7/MM5_d N_XI9/XI7/NET33_XI9/XI7/MM5_g
+ N_VDD_XI9/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI7/MM4 N_XI9/XI7/NET33_XI9/XI7/MM4_d N_XI9/XI7/NET34_XI9/XI7/MM4_g
+ N_VDD_XI9/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI7/MM10 N_XI9/XI7/NET35_XI9/XI7/MM10_d N_XI9/XI7/NET36_XI9/XI7/MM10_g
+ N_VDD_XI9/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI7/MM11 N_XI9/XI7/NET36_XI9/XI7/MM11_d N_XI9/XI7/NET35_XI9/XI7/MM11_g
+ N_VDD_XI9/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI8/MM2 N_XI9/XI8/NET34_XI9/XI8/MM2_d N_XI9/XI8/NET33_XI9/XI8/MM2_g
+ N_VSS_XI9/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM3 N_XI9/XI8/NET33_XI9/XI8/MM3_d N_WL<14>_XI9/XI8/MM3_g
+ N_BLN<7>_XI9/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM0 N_XI9/XI8/NET34_XI9/XI8/MM0_d N_WL<14>_XI9/XI8/MM0_g
+ N_BL<7>_XI9/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM1 N_XI9/XI8/NET33_XI9/XI8/MM1_d N_XI9/XI8/NET34_XI9/XI8/MM1_g
+ N_VSS_XI9/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM9 N_XI9/XI8/NET36_XI9/XI8/MM9_d N_WL<15>_XI9/XI8/MM9_g
+ N_BL<7>_XI9/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM6 N_XI9/XI8/NET35_XI9/XI8/MM6_d N_XI9/XI8/NET36_XI9/XI8/MM6_g
+ N_VSS_XI9/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM7 N_XI9/XI8/NET36_XI9/XI8/MM7_d N_XI9/XI8/NET35_XI9/XI8/MM7_g
+ N_VSS_XI9/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM8 N_XI9/XI8/NET35_XI9/XI8/MM8_d N_WL<15>_XI9/XI8/MM8_g
+ N_BLN<7>_XI9/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI8/MM5 N_XI9/XI8/NET34_XI9/XI8/MM5_d N_XI9/XI8/NET33_XI9/XI8/MM5_g
+ N_VDD_XI9/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI8/MM4 N_XI9/XI8/NET33_XI9/XI8/MM4_d N_XI9/XI8/NET34_XI9/XI8/MM4_g
+ N_VDD_XI9/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI8/MM10 N_XI9/XI8/NET35_XI9/XI8/MM10_d N_XI9/XI8/NET36_XI9/XI8/MM10_g
+ N_VDD_XI9/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI8/MM11 N_XI9/XI8/NET36_XI9/XI8/MM11_d N_XI9/XI8/NET35_XI9/XI8/MM11_g
+ N_VDD_XI9/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI9/MM2 N_XI9/XI9/NET34_XI9/XI9/MM2_d N_XI9/XI9/NET33_XI9/XI9/MM2_g
+ N_VSS_XI9/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM3 N_XI9/XI9/NET33_XI9/XI9/MM3_d N_WL<14>_XI9/XI9/MM3_g
+ N_BLN<6>_XI9/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM0 N_XI9/XI9/NET34_XI9/XI9/MM0_d N_WL<14>_XI9/XI9/MM0_g
+ N_BL<6>_XI9/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM1 N_XI9/XI9/NET33_XI9/XI9/MM1_d N_XI9/XI9/NET34_XI9/XI9/MM1_g
+ N_VSS_XI9/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM9 N_XI9/XI9/NET36_XI9/XI9/MM9_d N_WL<15>_XI9/XI9/MM9_g
+ N_BL<6>_XI9/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM6 N_XI9/XI9/NET35_XI9/XI9/MM6_d N_XI9/XI9/NET36_XI9/XI9/MM6_g
+ N_VSS_XI9/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM7 N_XI9/XI9/NET36_XI9/XI9/MM7_d N_XI9/XI9/NET35_XI9/XI9/MM7_g
+ N_VSS_XI9/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM8 N_XI9/XI9/NET35_XI9/XI9/MM8_d N_WL<15>_XI9/XI9/MM8_g
+ N_BLN<6>_XI9/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI9/MM5 N_XI9/XI9/NET34_XI9/XI9/MM5_d N_XI9/XI9/NET33_XI9/XI9/MM5_g
+ N_VDD_XI9/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI9/MM4 N_XI9/XI9/NET33_XI9/XI9/MM4_d N_XI9/XI9/NET34_XI9/XI9/MM4_g
+ N_VDD_XI9/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI9/MM10 N_XI9/XI9/NET35_XI9/XI9/MM10_d N_XI9/XI9/NET36_XI9/XI9/MM10_g
+ N_VDD_XI9/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI9/MM11 N_XI9/XI9/NET36_XI9/XI9/MM11_d N_XI9/XI9/NET35_XI9/XI9/MM11_g
+ N_VDD_XI9/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI10/MM2 N_XI9/XI10/NET34_XI9/XI10/MM2_d N_XI9/XI10/NET33_XI9/XI10/MM2_g
+ N_VSS_XI9/XI10/MM2_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI10/MM3 N_XI9/XI10/NET33_XI9/XI10/MM3_d N_WL<14>_XI9/XI10/MM3_g
+ N_BLN<5>_XI9/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI10/MM0 N_XI9/XI10/NET34_XI9/XI10/MM0_d N_WL<14>_XI9/XI10/MM0_g
+ N_BL<5>_XI9/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI10/MM1 N_XI9/XI10/NET33_XI9/XI10/MM1_d N_XI9/XI10/NET34_XI9/XI10/MM1_g
+ N_VSS_XI9/XI10/MM1_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI10/MM9 N_XI9/XI10/NET36_XI9/XI10/MM9_d N_WL<15>_XI9/XI10/MM9_g
+ N_BL<5>_XI9/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI10/MM6 N_XI9/XI10/NET35_XI9/XI10/MM6_d N_XI9/XI10/NET36_XI9/XI10/MM6_g
+ N_VSS_XI9/XI10/MM6_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI10/MM7 N_XI9/XI10/NET36_XI9/XI10/MM7_d N_XI9/XI10/NET35_XI9/XI10/MM7_g
+ N_VSS_XI9/XI10/MM7_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI10/MM8 N_XI9/XI10/NET35_XI9/XI10/MM8_d N_WL<15>_XI9/XI10/MM8_g
+ N_BLN<5>_XI9/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI10/MM5 N_XI9/XI10/NET34_XI9/XI10/MM5_d N_XI9/XI10/NET33_XI9/XI10/MM5_g
+ N_VDD_XI9/XI10/MM5_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI10/MM4 N_XI9/XI10/NET33_XI9/XI10/MM4_d N_XI9/XI10/NET34_XI9/XI10/MM4_g
+ N_VDD_XI9/XI10/MM4_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI10/MM10 N_XI9/XI10/NET35_XI9/XI10/MM10_d N_XI9/XI10/NET36_XI9/XI10/MM10_g
+ N_VDD_XI9/XI10/MM10_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI10/MM11 N_XI9/XI10/NET36_XI9/XI10/MM11_d N_XI9/XI10/NET35_XI9/XI10/MM11_g
+ N_VDD_XI9/XI10/MM11_s N_VDD_XI0/XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI11/MM2 N_XI9/XI11/NET34_XI9/XI11/MM2_d N_XI9/XI11/NET33_XI9/XI11/MM2_g
+ N_VSS_XI9/XI11/MM2_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI11/MM3 N_XI9/XI11/NET33_XI9/XI11/MM3_d N_WL<14>_XI9/XI11/MM3_g
+ N_BLN<4>_XI9/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI11/MM0 N_XI9/XI11/NET34_XI9/XI11/MM0_d N_WL<14>_XI9/XI11/MM0_g
+ N_BL<4>_XI9/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI11/MM1 N_XI9/XI11/NET33_XI9/XI11/MM1_d N_XI9/XI11/NET34_XI9/XI11/MM1_g
+ N_VSS_XI9/XI11/MM1_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI11/MM9 N_XI9/XI11/NET36_XI9/XI11/MM9_d N_WL<15>_XI9/XI11/MM9_g
+ N_BL<4>_XI9/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI11/MM6 N_XI9/XI11/NET35_XI9/XI11/MM6_d N_XI9/XI11/NET36_XI9/XI11/MM6_g
+ N_VSS_XI9/XI11/MM6_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI11/MM7 N_XI9/XI11/NET36_XI9/XI11/MM7_d N_XI9/XI11/NET35_XI9/XI11/MM7_g
+ N_VSS_XI9/XI11/MM7_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI11/MM8 N_XI9/XI11/NET35_XI9/XI11/MM8_d N_WL<15>_XI9/XI11/MM8_g
+ N_BLN<4>_XI9/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI11/MM5 N_XI9/XI11/NET34_XI9/XI11/MM5_d N_XI9/XI11/NET33_XI9/XI11/MM5_g
+ N_VDD_XI9/XI11/MM5_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI11/MM4 N_XI9/XI11/NET33_XI9/XI11/MM4_d N_XI9/XI11/NET34_XI9/XI11/MM4_g
+ N_VDD_XI9/XI11/MM4_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI11/MM10 N_XI9/XI11/NET35_XI9/XI11/MM10_d N_XI9/XI11/NET36_XI9/XI11/MM10_g
+ N_VDD_XI9/XI11/MM10_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI11/MM11 N_XI9/XI11/NET36_XI9/XI11/MM11_d N_XI9/XI11/NET35_XI9/XI11/MM11_g
+ N_VDD_XI9/XI11/MM11_s N_VDD_XI0/XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI12/MM2 N_XI9/XI12/NET34_XI9/XI12/MM2_d N_XI9/XI12/NET33_XI9/XI12/MM2_g
+ N_VSS_XI9/XI12/MM2_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI12/MM3 N_XI9/XI12/NET33_XI9/XI12/MM3_d N_WL<14>_XI9/XI12/MM3_g
+ N_BLN<3>_XI9/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI12/MM0 N_XI9/XI12/NET34_XI9/XI12/MM0_d N_WL<14>_XI9/XI12/MM0_g
+ N_BL<3>_XI9/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI12/MM1 N_XI9/XI12/NET33_XI9/XI12/MM1_d N_XI9/XI12/NET34_XI9/XI12/MM1_g
+ N_VSS_XI9/XI12/MM1_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI12/MM9 N_XI9/XI12/NET36_XI9/XI12/MM9_d N_WL<15>_XI9/XI12/MM9_g
+ N_BL<3>_XI9/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI12/MM6 N_XI9/XI12/NET35_XI9/XI12/MM6_d N_XI9/XI12/NET36_XI9/XI12/MM6_g
+ N_VSS_XI9/XI12/MM6_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI12/MM7 N_XI9/XI12/NET36_XI9/XI12/MM7_d N_XI9/XI12/NET35_XI9/XI12/MM7_g
+ N_VSS_XI9/XI12/MM7_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI12/MM8 N_XI9/XI12/NET35_XI9/XI12/MM8_d N_WL<15>_XI9/XI12/MM8_g
+ N_BLN<3>_XI9/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI12/MM5 N_XI9/XI12/NET34_XI9/XI12/MM5_d N_XI9/XI12/NET33_XI9/XI12/MM5_g
+ N_VDD_XI9/XI12/MM5_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI12/MM4 N_XI9/XI12/NET33_XI9/XI12/MM4_d N_XI9/XI12/NET34_XI9/XI12/MM4_g
+ N_VDD_XI9/XI12/MM4_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI12/MM10 N_XI9/XI12/NET35_XI9/XI12/MM10_d N_XI9/XI12/NET36_XI9/XI12/MM10_g
+ N_VDD_XI9/XI12/MM10_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI12/MM11 N_XI9/XI12/NET36_XI9/XI12/MM11_d N_XI9/XI12/NET35_XI9/XI12/MM11_g
+ N_VDD_XI9/XI12/MM11_s N_VDD_XI0/XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI13/MM2 N_XI9/XI13/NET34_XI9/XI13/MM2_d N_XI9/XI13/NET33_XI9/XI13/MM2_g
+ N_VSS_XI9/XI13/MM2_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI13/MM3 N_XI9/XI13/NET33_XI9/XI13/MM3_d N_WL<14>_XI9/XI13/MM3_g
+ N_BLN<2>_XI9/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI13/MM0 N_XI9/XI13/NET34_XI9/XI13/MM0_d N_WL<14>_XI9/XI13/MM0_g
+ N_BL<2>_XI9/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI13/MM1 N_XI9/XI13/NET33_XI9/XI13/MM1_d N_XI9/XI13/NET34_XI9/XI13/MM1_g
+ N_VSS_XI9/XI13/MM1_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI13/MM9 N_XI9/XI13/NET36_XI9/XI13/MM9_d N_WL<15>_XI9/XI13/MM9_g
+ N_BL<2>_XI9/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI13/MM6 N_XI9/XI13/NET35_XI9/XI13/MM6_d N_XI9/XI13/NET36_XI9/XI13/MM6_g
+ N_VSS_XI9/XI13/MM6_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI13/MM7 N_XI9/XI13/NET36_XI9/XI13/MM7_d N_XI9/XI13/NET35_XI9/XI13/MM7_g
+ N_VSS_XI9/XI13/MM7_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI13/MM8 N_XI9/XI13/NET35_XI9/XI13/MM8_d N_WL<15>_XI9/XI13/MM8_g
+ N_BLN<2>_XI9/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI13/MM5 N_XI9/XI13/NET34_XI9/XI13/MM5_d N_XI9/XI13/NET33_XI9/XI13/MM5_g
+ N_VDD_XI9/XI13/MM5_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI13/MM4 N_XI9/XI13/NET33_XI9/XI13/MM4_d N_XI9/XI13/NET34_XI9/XI13/MM4_g
+ N_VDD_XI9/XI13/MM4_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI13/MM10 N_XI9/XI13/NET35_XI9/XI13/MM10_d N_XI9/XI13/NET36_XI9/XI13/MM10_g
+ N_VDD_XI9/XI13/MM10_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI13/MM11 N_XI9/XI13/NET36_XI9/XI13/MM11_d N_XI9/XI13/NET35_XI9/XI13/MM11_g
+ N_VDD_XI9/XI13/MM11_s N_VDD_XI0/XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI14/MM2 N_XI9/XI14/NET34_XI9/XI14/MM2_d N_XI9/XI14/NET33_XI9/XI14/MM2_g
+ N_VSS_XI9/XI14/MM2_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI14/MM3 N_XI9/XI14/NET33_XI9/XI14/MM3_d N_WL<14>_XI9/XI14/MM3_g
+ N_BLN<1>_XI9/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI14/MM0 N_XI9/XI14/NET34_XI9/XI14/MM0_d N_WL<14>_XI9/XI14/MM0_g
+ N_BL<1>_XI9/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI14/MM1 N_XI9/XI14/NET33_XI9/XI14/MM1_d N_XI9/XI14/NET34_XI9/XI14/MM1_g
+ N_VSS_XI9/XI14/MM1_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI14/MM9 N_XI9/XI14/NET36_XI9/XI14/MM9_d N_WL<15>_XI9/XI14/MM9_g
+ N_BL<1>_XI9/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI14/MM6 N_XI9/XI14/NET35_XI9/XI14/MM6_d N_XI9/XI14/NET36_XI9/XI14/MM6_g
+ N_VSS_XI9/XI14/MM6_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI14/MM7 N_XI9/XI14/NET36_XI9/XI14/MM7_d N_XI9/XI14/NET35_XI9/XI14/MM7_g
+ N_VSS_XI9/XI14/MM7_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI14/MM8 N_XI9/XI14/NET35_XI9/XI14/MM8_d N_WL<15>_XI9/XI14/MM8_g
+ N_BLN<1>_XI9/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI14/MM5 N_XI9/XI14/NET34_XI9/XI14/MM5_d N_XI9/XI14/NET33_XI9/XI14/MM5_g
+ N_VDD_XI9/XI14/MM5_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI14/MM4 N_XI9/XI14/NET33_XI9/XI14/MM4_d N_XI9/XI14/NET34_XI9/XI14/MM4_g
+ N_VDD_XI9/XI14/MM4_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI14/MM10 N_XI9/XI14/NET35_XI9/XI14/MM10_d N_XI9/XI14/NET36_XI9/XI14/MM10_g
+ N_VDD_XI9/XI14/MM10_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI14/MM11 N_XI9/XI14/NET36_XI9/XI14/MM11_d N_XI9/XI14/NET35_XI9/XI14/MM11_g
+ N_VDD_XI9/XI14/MM11_s N_VDD_XI0/XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI15/MM2 N_XI9/XI15/NET34_XI9/XI15/MM2_d N_XI9/XI15/NET33_XI9/XI15/MM2_g
+ N_VSS_XI9/XI15/MM2_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI15/MM3 N_XI9/XI15/NET33_XI9/XI15/MM3_d N_WL<14>_XI9/XI15/MM3_g
+ N_BLN<0>_XI9/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI15/MM0 N_XI9/XI15/NET34_XI9/XI15/MM0_d N_WL<14>_XI9/XI15/MM0_g
+ N_BL<0>_XI9/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI15/MM1 N_XI9/XI15/NET33_XI9/XI15/MM1_d N_XI9/XI15/NET34_XI9/XI15/MM1_g
+ N_VSS_XI9/XI15/MM1_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI15/MM9 N_XI9/XI15/NET36_XI9/XI15/MM9_d N_WL<15>_XI9/XI15/MM9_g
+ N_BL<0>_XI9/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI15/MM6 N_XI9/XI15/NET35_XI9/XI15/MM6_d N_XI9/XI15/NET36_XI9/XI15/MM6_g
+ N_VSS_XI9/XI15/MM6_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI15/MM7 N_XI9/XI15/NET36_XI9/XI15/MM7_d N_XI9/XI15/NET35_XI9/XI15/MM7_g
+ N_VSS_XI9/XI15/MM7_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/XI15/MM8 N_XI9/XI15/NET35_XI9/XI15/MM8_d N_WL<15>_XI9/XI15/MM8_g
+ N_BLN<0>_XI9/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI9/XI15/MM5 N_XI9/XI15/NET34_XI9/XI15/MM5_d N_XI9/XI15/NET33_XI9/XI15/MM5_g
+ N_VDD_XI9/XI15/MM5_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI15/MM4 N_XI9/XI15/NET33_XI9/XI15/MM4_d N_XI9/XI15/NET34_XI9/XI15/MM4_g
+ N_VDD_XI9/XI15/MM4_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI15/MM10 N_XI9/XI15/NET35_XI9/XI15/MM10_d N_XI9/XI15/NET36_XI9/XI15/MM10_g
+ N_VDD_XI9/XI15/MM10_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/XI15/MM11 N_XI9/XI15/NET36_XI9/XI15/MM11_d N_XI9/XI15/NET35_XI9/XI15/MM11_g
+ N_VDD_XI9/XI15/MM11_s N_VDD_XI0/XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI0/MM2 N_XI10/XI0/NET34_XI10/XI0/MM2_d N_XI10/XI0/NET33_XI10/XI0/MM2_g
+ N_VSS_XI10/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI0/MM3 N_XI10/XI0/NET33_XI10/XI0/MM3_d N_WL<16>_XI10/XI0/MM3_g
+ N_BLN<15>_XI10/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI0/MM0 N_XI10/XI0/NET34_XI10/XI0/MM0_d N_WL<16>_XI10/XI0/MM0_g
+ N_BL<15>_XI10/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI0/MM1 N_XI10/XI0/NET33_XI10/XI0/MM1_d N_XI10/XI0/NET34_XI10/XI0/MM1_g
+ N_VSS_XI10/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI0/MM9 N_XI10/XI0/NET36_XI10/XI0/MM9_d N_WL<17>_XI10/XI0/MM9_g
+ N_BL<15>_XI10/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI0/MM6 N_XI10/XI0/NET35_XI10/XI0/MM6_d N_XI10/XI0/NET36_XI10/XI0/MM6_g
+ N_VSS_XI10/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI0/MM7 N_XI10/XI0/NET36_XI10/XI0/MM7_d N_XI10/XI0/NET35_XI10/XI0/MM7_g
+ N_VSS_XI10/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI0/MM8 N_XI10/XI0/NET35_XI10/XI0/MM8_d N_WL<17>_XI10/XI0/MM8_g
+ N_BLN<15>_XI10/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI0/MM5 N_XI10/XI0/NET34_XI10/XI0/MM5_d N_XI10/XI0/NET33_XI10/XI0/MM5_g
+ N_VDD_XI10/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI0/MM4 N_XI10/XI0/NET33_XI10/XI0/MM4_d N_XI10/XI0/NET34_XI10/XI0/MM4_g
+ N_VDD_XI10/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI0/MM10 N_XI10/XI0/NET35_XI10/XI0/MM10_d N_XI10/XI0/NET36_XI10/XI0/MM10_g
+ N_VDD_XI10/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI0/MM11 N_XI10/XI0/NET36_XI10/XI0/MM11_d N_XI10/XI0/NET35_XI10/XI0/MM11_g
+ N_VDD_XI10/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI1/MM2 N_XI10/XI1/NET34_XI10/XI1/MM2_d N_XI10/XI1/NET33_XI10/XI1/MM2_g
+ N_VSS_XI10/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI1/MM3 N_XI10/XI1/NET33_XI10/XI1/MM3_d N_WL<16>_XI10/XI1/MM3_g
+ N_BLN<14>_XI10/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI1/MM0 N_XI10/XI1/NET34_XI10/XI1/MM0_d N_WL<16>_XI10/XI1/MM0_g
+ N_BL<14>_XI10/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI1/MM1 N_XI10/XI1/NET33_XI10/XI1/MM1_d N_XI10/XI1/NET34_XI10/XI1/MM1_g
+ N_VSS_XI10/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI1/MM9 N_XI10/XI1/NET36_XI10/XI1/MM9_d N_WL<17>_XI10/XI1/MM9_g
+ N_BL<14>_XI10/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI1/MM6 N_XI10/XI1/NET35_XI10/XI1/MM6_d N_XI10/XI1/NET36_XI10/XI1/MM6_g
+ N_VSS_XI10/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI1/MM7 N_XI10/XI1/NET36_XI10/XI1/MM7_d N_XI10/XI1/NET35_XI10/XI1/MM7_g
+ N_VSS_XI10/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI1/MM8 N_XI10/XI1/NET35_XI10/XI1/MM8_d N_WL<17>_XI10/XI1/MM8_g
+ N_BLN<14>_XI10/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI1/MM5 N_XI10/XI1/NET34_XI10/XI1/MM5_d N_XI10/XI1/NET33_XI10/XI1/MM5_g
+ N_VDD_XI10/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI1/MM4 N_XI10/XI1/NET33_XI10/XI1/MM4_d N_XI10/XI1/NET34_XI10/XI1/MM4_g
+ N_VDD_XI10/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI1/MM10 N_XI10/XI1/NET35_XI10/XI1/MM10_d N_XI10/XI1/NET36_XI10/XI1/MM10_g
+ N_VDD_XI10/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI1/MM11 N_XI10/XI1/NET36_XI10/XI1/MM11_d N_XI10/XI1/NET35_XI10/XI1/MM11_g
+ N_VDD_XI10/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI2/MM2 N_XI10/XI2/NET34_XI10/XI2/MM2_d N_XI10/XI2/NET33_XI10/XI2/MM2_g
+ N_VSS_XI10/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI2/MM3 N_XI10/XI2/NET33_XI10/XI2/MM3_d N_WL<16>_XI10/XI2/MM3_g
+ N_BLN<13>_XI10/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI2/MM0 N_XI10/XI2/NET34_XI10/XI2/MM0_d N_WL<16>_XI10/XI2/MM0_g
+ N_BL<13>_XI10/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI2/MM1 N_XI10/XI2/NET33_XI10/XI2/MM1_d N_XI10/XI2/NET34_XI10/XI2/MM1_g
+ N_VSS_XI10/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI2/MM9 N_XI10/XI2/NET36_XI10/XI2/MM9_d N_WL<17>_XI10/XI2/MM9_g
+ N_BL<13>_XI10/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI2/MM6 N_XI10/XI2/NET35_XI10/XI2/MM6_d N_XI10/XI2/NET36_XI10/XI2/MM6_g
+ N_VSS_XI10/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI2/MM7 N_XI10/XI2/NET36_XI10/XI2/MM7_d N_XI10/XI2/NET35_XI10/XI2/MM7_g
+ N_VSS_XI10/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI2/MM8 N_XI10/XI2/NET35_XI10/XI2/MM8_d N_WL<17>_XI10/XI2/MM8_g
+ N_BLN<13>_XI10/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI2/MM5 N_XI10/XI2/NET34_XI10/XI2/MM5_d N_XI10/XI2/NET33_XI10/XI2/MM5_g
+ N_VDD_XI10/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI2/MM4 N_XI10/XI2/NET33_XI10/XI2/MM4_d N_XI10/XI2/NET34_XI10/XI2/MM4_g
+ N_VDD_XI10/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI2/MM10 N_XI10/XI2/NET35_XI10/XI2/MM10_d N_XI10/XI2/NET36_XI10/XI2/MM10_g
+ N_VDD_XI10/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI2/MM11 N_XI10/XI2/NET36_XI10/XI2/MM11_d N_XI10/XI2/NET35_XI10/XI2/MM11_g
+ N_VDD_XI10/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI3/MM2 N_XI10/XI3/NET34_XI10/XI3/MM2_d N_XI10/XI3/NET33_XI10/XI3/MM2_g
+ N_VSS_XI10/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI3/MM3 N_XI10/XI3/NET33_XI10/XI3/MM3_d N_WL<16>_XI10/XI3/MM3_g
+ N_BLN<12>_XI10/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI3/MM0 N_XI10/XI3/NET34_XI10/XI3/MM0_d N_WL<16>_XI10/XI3/MM0_g
+ N_BL<12>_XI10/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI3/MM1 N_XI10/XI3/NET33_XI10/XI3/MM1_d N_XI10/XI3/NET34_XI10/XI3/MM1_g
+ N_VSS_XI10/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI3/MM9 N_XI10/XI3/NET36_XI10/XI3/MM9_d N_WL<17>_XI10/XI3/MM9_g
+ N_BL<12>_XI10/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI3/MM6 N_XI10/XI3/NET35_XI10/XI3/MM6_d N_XI10/XI3/NET36_XI10/XI3/MM6_g
+ N_VSS_XI10/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI3/MM7 N_XI10/XI3/NET36_XI10/XI3/MM7_d N_XI10/XI3/NET35_XI10/XI3/MM7_g
+ N_VSS_XI10/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI3/MM8 N_XI10/XI3/NET35_XI10/XI3/MM8_d N_WL<17>_XI10/XI3/MM8_g
+ N_BLN<12>_XI10/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI3/MM5 N_XI10/XI3/NET34_XI10/XI3/MM5_d N_XI10/XI3/NET33_XI10/XI3/MM5_g
+ N_VDD_XI10/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI3/MM4 N_XI10/XI3/NET33_XI10/XI3/MM4_d N_XI10/XI3/NET34_XI10/XI3/MM4_g
+ N_VDD_XI10/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI3/MM10 N_XI10/XI3/NET35_XI10/XI3/MM10_d N_XI10/XI3/NET36_XI10/XI3/MM10_g
+ N_VDD_XI10/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI3/MM11 N_XI10/XI3/NET36_XI10/XI3/MM11_d N_XI10/XI3/NET35_XI10/XI3/MM11_g
+ N_VDD_XI10/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI4/MM2 N_XI10/XI4/NET34_XI10/XI4/MM2_d N_XI10/XI4/NET33_XI10/XI4/MM2_g
+ N_VSS_XI10/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI4/MM3 N_XI10/XI4/NET33_XI10/XI4/MM3_d N_WL<16>_XI10/XI4/MM3_g
+ N_BLN<11>_XI10/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI4/MM0 N_XI10/XI4/NET34_XI10/XI4/MM0_d N_WL<16>_XI10/XI4/MM0_g
+ N_BL<11>_XI10/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI4/MM1 N_XI10/XI4/NET33_XI10/XI4/MM1_d N_XI10/XI4/NET34_XI10/XI4/MM1_g
+ N_VSS_XI10/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI4/MM9 N_XI10/XI4/NET36_XI10/XI4/MM9_d N_WL<17>_XI10/XI4/MM9_g
+ N_BL<11>_XI10/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI4/MM6 N_XI10/XI4/NET35_XI10/XI4/MM6_d N_XI10/XI4/NET36_XI10/XI4/MM6_g
+ N_VSS_XI10/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI4/MM7 N_XI10/XI4/NET36_XI10/XI4/MM7_d N_XI10/XI4/NET35_XI10/XI4/MM7_g
+ N_VSS_XI10/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI4/MM8 N_XI10/XI4/NET35_XI10/XI4/MM8_d N_WL<17>_XI10/XI4/MM8_g
+ N_BLN<11>_XI10/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI4/MM5 N_XI10/XI4/NET34_XI10/XI4/MM5_d N_XI10/XI4/NET33_XI10/XI4/MM5_g
+ N_VDD_XI10/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI4/MM4 N_XI10/XI4/NET33_XI10/XI4/MM4_d N_XI10/XI4/NET34_XI10/XI4/MM4_g
+ N_VDD_XI10/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI4/MM10 N_XI10/XI4/NET35_XI10/XI4/MM10_d N_XI10/XI4/NET36_XI10/XI4/MM10_g
+ N_VDD_XI10/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI4/MM11 N_XI10/XI4/NET36_XI10/XI4/MM11_d N_XI10/XI4/NET35_XI10/XI4/MM11_g
+ N_VDD_XI10/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI5/MM2 N_XI10/XI5/NET34_XI10/XI5/MM2_d N_XI10/XI5/NET33_XI10/XI5/MM2_g
+ N_VSS_XI10/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI5/MM3 N_XI10/XI5/NET33_XI10/XI5/MM3_d N_WL<16>_XI10/XI5/MM3_g
+ N_BLN<10>_XI10/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI5/MM0 N_XI10/XI5/NET34_XI10/XI5/MM0_d N_WL<16>_XI10/XI5/MM0_g
+ N_BL<10>_XI10/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI5/MM1 N_XI10/XI5/NET33_XI10/XI5/MM1_d N_XI10/XI5/NET34_XI10/XI5/MM1_g
+ N_VSS_XI10/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI5/MM9 N_XI10/XI5/NET36_XI10/XI5/MM9_d N_WL<17>_XI10/XI5/MM9_g
+ N_BL<10>_XI10/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI5/MM6 N_XI10/XI5/NET35_XI10/XI5/MM6_d N_XI10/XI5/NET36_XI10/XI5/MM6_g
+ N_VSS_XI10/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI5/MM7 N_XI10/XI5/NET36_XI10/XI5/MM7_d N_XI10/XI5/NET35_XI10/XI5/MM7_g
+ N_VSS_XI10/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI5/MM8 N_XI10/XI5/NET35_XI10/XI5/MM8_d N_WL<17>_XI10/XI5/MM8_g
+ N_BLN<10>_XI10/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI5/MM5 N_XI10/XI5/NET34_XI10/XI5/MM5_d N_XI10/XI5/NET33_XI10/XI5/MM5_g
+ N_VDD_XI10/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI5/MM4 N_XI10/XI5/NET33_XI10/XI5/MM4_d N_XI10/XI5/NET34_XI10/XI5/MM4_g
+ N_VDD_XI10/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI5/MM10 N_XI10/XI5/NET35_XI10/XI5/MM10_d N_XI10/XI5/NET36_XI10/XI5/MM10_g
+ N_VDD_XI10/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI5/MM11 N_XI10/XI5/NET36_XI10/XI5/MM11_d N_XI10/XI5/NET35_XI10/XI5/MM11_g
+ N_VDD_XI10/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI6/MM2 N_XI10/XI6/NET34_XI10/XI6/MM2_d N_XI10/XI6/NET33_XI10/XI6/MM2_g
+ N_VSS_XI10/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM3 N_XI10/XI6/NET33_XI10/XI6/MM3_d N_WL<16>_XI10/XI6/MM3_g
+ N_BLN<9>_XI10/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM0 N_XI10/XI6/NET34_XI10/XI6/MM0_d N_WL<16>_XI10/XI6/MM0_g
+ N_BL<9>_XI10/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM1 N_XI10/XI6/NET33_XI10/XI6/MM1_d N_XI10/XI6/NET34_XI10/XI6/MM1_g
+ N_VSS_XI10/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM9 N_XI10/XI6/NET36_XI10/XI6/MM9_d N_WL<17>_XI10/XI6/MM9_g
+ N_BL<9>_XI10/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM6 N_XI10/XI6/NET35_XI10/XI6/MM6_d N_XI10/XI6/NET36_XI10/XI6/MM6_g
+ N_VSS_XI10/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM7 N_XI10/XI6/NET36_XI10/XI6/MM7_d N_XI10/XI6/NET35_XI10/XI6/MM7_g
+ N_VSS_XI10/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM8 N_XI10/XI6/NET35_XI10/XI6/MM8_d N_WL<17>_XI10/XI6/MM8_g
+ N_BLN<9>_XI10/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI6/MM5 N_XI10/XI6/NET34_XI10/XI6/MM5_d N_XI10/XI6/NET33_XI10/XI6/MM5_g
+ N_VDD_XI10/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI6/MM4 N_XI10/XI6/NET33_XI10/XI6/MM4_d N_XI10/XI6/NET34_XI10/XI6/MM4_g
+ N_VDD_XI10/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI6/MM10 N_XI10/XI6/NET35_XI10/XI6/MM10_d N_XI10/XI6/NET36_XI10/XI6/MM10_g
+ N_VDD_XI10/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI6/MM11 N_XI10/XI6/NET36_XI10/XI6/MM11_d N_XI10/XI6/NET35_XI10/XI6/MM11_g
+ N_VDD_XI10/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI7/MM2 N_XI10/XI7/NET34_XI10/XI7/MM2_d N_XI10/XI7/NET33_XI10/XI7/MM2_g
+ N_VSS_XI10/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM3 N_XI10/XI7/NET33_XI10/XI7/MM3_d N_WL<16>_XI10/XI7/MM3_g
+ N_BLN<8>_XI10/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM0 N_XI10/XI7/NET34_XI10/XI7/MM0_d N_WL<16>_XI10/XI7/MM0_g
+ N_BL<8>_XI10/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM1 N_XI10/XI7/NET33_XI10/XI7/MM1_d N_XI10/XI7/NET34_XI10/XI7/MM1_g
+ N_VSS_XI10/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM9 N_XI10/XI7/NET36_XI10/XI7/MM9_d N_WL<17>_XI10/XI7/MM9_g
+ N_BL<8>_XI10/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM6 N_XI10/XI7/NET35_XI10/XI7/MM6_d N_XI10/XI7/NET36_XI10/XI7/MM6_g
+ N_VSS_XI10/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM7 N_XI10/XI7/NET36_XI10/XI7/MM7_d N_XI10/XI7/NET35_XI10/XI7/MM7_g
+ N_VSS_XI10/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM8 N_XI10/XI7/NET35_XI10/XI7/MM8_d N_WL<17>_XI10/XI7/MM8_g
+ N_BLN<8>_XI10/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI7/MM5 N_XI10/XI7/NET34_XI10/XI7/MM5_d N_XI10/XI7/NET33_XI10/XI7/MM5_g
+ N_VDD_XI10/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI7/MM4 N_XI10/XI7/NET33_XI10/XI7/MM4_d N_XI10/XI7/NET34_XI10/XI7/MM4_g
+ N_VDD_XI10/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI7/MM10 N_XI10/XI7/NET35_XI10/XI7/MM10_d N_XI10/XI7/NET36_XI10/XI7/MM10_g
+ N_VDD_XI10/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI7/MM11 N_XI10/XI7/NET36_XI10/XI7/MM11_d N_XI10/XI7/NET35_XI10/XI7/MM11_g
+ N_VDD_XI10/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI8/MM2 N_XI10/XI8/NET34_XI10/XI8/MM2_d N_XI10/XI8/NET33_XI10/XI8/MM2_g
+ N_VSS_XI10/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM3 N_XI10/XI8/NET33_XI10/XI8/MM3_d N_WL<16>_XI10/XI8/MM3_g
+ N_BLN<7>_XI10/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM0 N_XI10/XI8/NET34_XI10/XI8/MM0_d N_WL<16>_XI10/XI8/MM0_g
+ N_BL<7>_XI10/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM1 N_XI10/XI8/NET33_XI10/XI8/MM1_d N_XI10/XI8/NET34_XI10/XI8/MM1_g
+ N_VSS_XI10/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM9 N_XI10/XI8/NET36_XI10/XI8/MM9_d N_WL<17>_XI10/XI8/MM9_g
+ N_BL<7>_XI10/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM6 N_XI10/XI8/NET35_XI10/XI8/MM6_d N_XI10/XI8/NET36_XI10/XI8/MM6_g
+ N_VSS_XI10/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM7 N_XI10/XI8/NET36_XI10/XI8/MM7_d N_XI10/XI8/NET35_XI10/XI8/MM7_g
+ N_VSS_XI10/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM8 N_XI10/XI8/NET35_XI10/XI8/MM8_d N_WL<17>_XI10/XI8/MM8_g
+ N_BLN<7>_XI10/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI8/MM5 N_XI10/XI8/NET34_XI10/XI8/MM5_d N_XI10/XI8/NET33_XI10/XI8/MM5_g
+ N_VDD_XI10/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI8/MM4 N_XI10/XI8/NET33_XI10/XI8/MM4_d N_XI10/XI8/NET34_XI10/XI8/MM4_g
+ N_VDD_XI10/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI8/MM10 N_XI10/XI8/NET35_XI10/XI8/MM10_d N_XI10/XI8/NET36_XI10/XI8/MM10_g
+ N_VDD_XI10/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI8/MM11 N_XI10/XI8/NET36_XI10/XI8/MM11_d N_XI10/XI8/NET35_XI10/XI8/MM11_g
+ N_VDD_XI10/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI9/MM2 N_XI10/XI9/NET34_XI10/XI9/MM2_d N_XI10/XI9/NET33_XI10/XI9/MM2_g
+ N_VSS_XI10/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM3 N_XI10/XI9/NET33_XI10/XI9/MM3_d N_WL<16>_XI10/XI9/MM3_g
+ N_BLN<6>_XI10/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM0 N_XI10/XI9/NET34_XI10/XI9/MM0_d N_WL<16>_XI10/XI9/MM0_g
+ N_BL<6>_XI10/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM1 N_XI10/XI9/NET33_XI10/XI9/MM1_d N_XI10/XI9/NET34_XI10/XI9/MM1_g
+ N_VSS_XI10/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM9 N_XI10/XI9/NET36_XI10/XI9/MM9_d N_WL<17>_XI10/XI9/MM9_g
+ N_BL<6>_XI10/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM6 N_XI10/XI9/NET35_XI10/XI9/MM6_d N_XI10/XI9/NET36_XI10/XI9/MM6_g
+ N_VSS_XI10/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM7 N_XI10/XI9/NET36_XI10/XI9/MM7_d N_XI10/XI9/NET35_XI10/XI9/MM7_g
+ N_VSS_XI10/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM8 N_XI10/XI9/NET35_XI10/XI9/MM8_d N_WL<17>_XI10/XI9/MM8_g
+ N_BLN<6>_XI10/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI9/MM5 N_XI10/XI9/NET34_XI10/XI9/MM5_d N_XI10/XI9/NET33_XI10/XI9/MM5_g
+ N_VDD_XI10/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI9/MM4 N_XI10/XI9/NET33_XI10/XI9/MM4_d N_XI10/XI9/NET34_XI10/XI9/MM4_g
+ N_VDD_XI10/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI9/MM10 N_XI10/XI9/NET35_XI10/XI9/MM10_d N_XI10/XI9/NET36_XI10/XI9/MM10_g
+ N_VDD_XI10/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI9/MM11 N_XI10/XI9/NET36_XI10/XI9/MM11_d N_XI10/XI9/NET35_XI10/XI9/MM11_g
+ N_VDD_XI10/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI10/MM2 N_XI10/XI10/NET34_XI10/XI10/MM2_d
+ N_XI10/XI10/NET33_XI10/XI10/MM2_g N_VSS_XI10/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI10/MM3 N_XI10/XI10/NET33_XI10/XI10/MM3_d N_WL<16>_XI10/XI10/MM3_g
+ N_BLN<5>_XI10/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI10/MM0 N_XI10/XI10/NET34_XI10/XI10/MM0_d N_WL<16>_XI10/XI10/MM0_g
+ N_BL<5>_XI10/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI10/MM1 N_XI10/XI10/NET33_XI10/XI10/MM1_d
+ N_XI10/XI10/NET34_XI10/XI10/MM1_g N_VSS_XI10/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI10/MM9 N_XI10/XI10/NET36_XI10/XI10/MM9_d N_WL<17>_XI10/XI10/MM9_g
+ N_BL<5>_XI10/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI10/MM6 N_XI10/XI10/NET35_XI10/XI10/MM6_d
+ N_XI10/XI10/NET36_XI10/XI10/MM6_g N_VSS_XI10/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI10/MM7 N_XI10/XI10/NET36_XI10/XI10/MM7_d
+ N_XI10/XI10/NET35_XI10/XI10/MM7_g N_VSS_XI10/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI10/MM8 N_XI10/XI10/NET35_XI10/XI10/MM8_d N_WL<17>_XI10/XI10/MM8_g
+ N_BLN<5>_XI10/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI10/MM5 N_XI10/XI10/NET34_XI10/XI10/MM5_d
+ N_XI10/XI10/NET33_XI10/XI10/MM5_g N_VDD_XI10/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI10/MM4 N_XI10/XI10/NET33_XI10/XI10/MM4_d
+ N_XI10/XI10/NET34_XI10/XI10/MM4_g N_VDD_XI10/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI10/MM10 N_XI10/XI10/NET35_XI10/XI10/MM10_d
+ N_XI10/XI10/NET36_XI10/XI10/MM10_g N_VDD_XI10/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI10/MM11 N_XI10/XI10/NET36_XI10/XI10/MM11_d
+ N_XI10/XI10/NET35_XI10/XI10/MM11_g N_VDD_XI10/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI11/MM2 N_XI10/XI11/NET34_XI10/XI11/MM2_d
+ N_XI10/XI11/NET33_XI10/XI11/MM2_g N_VSS_XI10/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI11/MM3 N_XI10/XI11/NET33_XI10/XI11/MM3_d N_WL<16>_XI10/XI11/MM3_g
+ N_BLN<4>_XI10/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI11/MM0 N_XI10/XI11/NET34_XI10/XI11/MM0_d N_WL<16>_XI10/XI11/MM0_g
+ N_BL<4>_XI10/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI11/MM1 N_XI10/XI11/NET33_XI10/XI11/MM1_d
+ N_XI10/XI11/NET34_XI10/XI11/MM1_g N_VSS_XI10/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI11/MM9 N_XI10/XI11/NET36_XI10/XI11/MM9_d N_WL<17>_XI10/XI11/MM9_g
+ N_BL<4>_XI10/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI11/MM6 N_XI10/XI11/NET35_XI10/XI11/MM6_d
+ N_XI10/XI11/NET36_XI10/XI11/MM6_g N_VSS_XI10/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI11/MM7 N_XI10/XI11/NET36_XI10/XI11/MM7_d
+ N_XI10/XI11/NET35_XI10/XI11/MM7_g N_VSS_XI10/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI11/MM8 N_XI10/XI11/NET35_XI10/XI11/MM8_d N_WL<17>_XI10/XI11/MM8_g
+ N_BLN<4>_XI10/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI11/MM5 N_XI10/XI11/NET34_XI10/XI11/MM5_d
+ N_XI10/XI11/NET33_XI10/XI11/MM5_g N_VDD_XI10/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI11/MM4 N_XI10/XI11/NET33_XI10/XI11/MM4_d
+ N_XI10/XI11/NET34_XI10/XI11/MM4_g N_VDD_XI10/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI11/MM10 N_XI10/XI11/NET35_XI10/XI11/MM10_d
+ N_XI10/XI11/NET36_XI10/XI11/MM10_g N_VDD_XI10/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI11/MM11 N_XI10/XI11/NET36_XI10/XI11/MM11_d
+ N_XI10/XI11/NET35_XI10/XI11/MM11_g N_VDD_XI10/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI12/MM2 N_XI10/XI12/NET34_XI10/XI12/MM2_d
+ N_XI10/XI12/NET33_XI10/XI12/MM2_g N_VSS_XI10/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI12/MM3 N_XI10/XI12/NET33_XI10/XI12/MM3_d N_WL<16>_XI10/XI12/MM3_g
+ N_BLN<3>_XI10/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI12/MM0 N_XI10/XI12/NET34_XI10/XI12/MM0_d N_WL<16>_XI10/XI12/MM0_g
+ N_BL<3>_XI10/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI12/MM1 N_XI10/XI12/NET33_XI10/XI12/MM1_d
+ N_XI10/XI12/NET34_XI10/XI12/MM1_g N_VSS_XI10/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI12/MM9 N_XI10/XI12/NET36_XI10/XI12/MM9_d N_WL<17>_XI10/XI12/MM9_g
+ N_BL<3>_XI10/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI12/MM6 N_XI10/XI12/NET35_XI10/XI12/MM6_d
+ N_XI10/XI12/NET36_XI10/XI12/MM6_g N_VSS_XI10/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI12/MM7 N_XI10/XI12/NET36_XI10/XI12/MM7_d
+ N_XI10/XI12/NET35_XI10/XI12/MM7_g N_VSS_XI10/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI12/MM8 N_XI10/XI12/NET35_XI10/XI12/MM8_d N_WL<17>_XI10/XI12/MM8_g
+ N_BLN<3>_XI10/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI12/MM5 N_XI10/XI12/NET34_XI10/XI12/MM5_d
+ N_XI10/XI12/NET33_XI10/XI12/MM5_g N_VDD_XI10/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI12/MM4 N_XI10/XI12/NET33_XI10/XI12/MM4_d
+ N_XI10/XI12/NET34_XI10/XI12/MM4_g N_VDD_XI10/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI12/MM10 N_XI10/XI12/NET35_XI10/XI12/MM10_d
+ N_XI10/XI12/NET36_XI10/XI12/MM10_g N_VDD_XI10/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI12/MM11 N_XI10/XI12/NET36_XI10/XI12/MM11_d
+ N_XI10/XI12/NET35_XI10/XI12/MM11_g N_VDD_XI10/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI13/MM2 N_XI10/XI13/NET34_XI10/XI13/MM2_d
+ N_XI10/XI13/NET33_XI10/XI13/MM2_g N_VSS_XI10/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI13/MM3 N_XI10/XI13/NET33_XI10/XI13/MM3_d N_WL<16>_XI10/XI13/MM3_g
+ N_BLN<2>_XI10/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI13/MM0 N_XI10/XI13/NET34_XI10/XI13/MM0_d N_WL<16>_XI10/XI13/MM0_g
+ N_BL<2>_XI10/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI13/MM1 N_XI10/XI13/NET33_XI10/XI13/MM1_d
+ N_XI10/XI13/NET34_XI10/XI13/MM1_g N_VSS_XI10/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI13/MM9 N_XI10/XI13/NET36_XI10/XI13/MM9_d N_WL<17>_XI10/XI13/MM9_g
+ N_BL<2>_XI10/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI13/MM6 N_XI10/XI13/NET35_XI10/XI13/MM6_d
+ N_XI10/XI13/NET36_XI10/XI13/MM6_g N_VSS_XI10/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI13/MM7 N_XI10/XI13/NET36_XI10/XI13/MM7_d
+ N_XI10/XI13/NET35_XI10/XI13/MM7_g N_VSS_XI10/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI13/MM8 N_XI10/XI13/NET35_XI10/XI13/MM8_d N_WL<17>_XI10/XI13/MM8_g
+ N_BLN<2>_XI10/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI13/MM5 N_XI10/XI13/NET34_XI10/XI13/MM5_d
+ N_XI10/XI13/NET33_XI10/XI13/MM5_g N_VDD_XI10/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI13/MM4 N_XI10/XI13/NET33_XI10/XI13/MM4_d
+ N_XI10/XI13/NET34_XI10/XI13/MM4_g N_VDD_XI10/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI13/MM10 N_XI10/XI13/NET35_XI10/XI13/MM10_d
+ N_XI10/XI13/NET36_XI10/XI13/MM10_g N_VDD_XI10/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI13/MM11 N_XI10/XI13/NET36_XI10/XI13/MM11_d
+ N_XI10/XI13/NET35_XI10/XI13/MM11_g N_VDD_XI10/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI14/MM2 N_XI10/XI14/NET34_XI10/XI14/MM2_d
+ N_XI10/XI14/NET33_XI10/XI14/MM2_g N_VSS_XI10/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI14/MM3 N_XI10/XI14/NET33_XI10/XI14/MM3_d N_WL<16>_XI10/XI14/MM3_g
+ N_BLN<1>_XI10/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI14/MM0 N_XI10/XI14/NET34_XI10/XI14/MM0_d N_WL<16>_XI10/XI14/MM0_g
+ N_BL<1>_XI10/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI14/MM1 N_XI10/XI14/NET33_XI10/XI14/MM1_d
+ N_XI10/XI14/NET34_XI10/XI14/MM1_g N_VSS_XI10/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI14/MM9 N_XI10/XI14/NET36_XI10/XI14/MM9_d N_WL<17>_XI10/XI14/MM9_g
+ N_BL<1>_XI10/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI14/MM6 N_XI10/XI14/NET35_XI10/XI14/MM6_d
+ N_XI10/XI14/NET36_XI10/XI14/MM6_g N_VSS_XI10/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI14/MM7 N_XI10/XI14/NET36_XI10/XI14/MM7_d
+ N_XI10/XI14/NET35_XI10/XI14/MM7_g N_VSS_XI10/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI14/MM8 N_XI10/XI14/NET35_XI10/XI14/MM8_d N_WL<17>_XI10/XI14/MM8_g
+ N_BLN<1>_XI10/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI14/MM5 N_XI10/XI14/NET34_XI10/XI14/MM5_d
+ N_XI10/XI14/NET33_XI10/XI14/MM5_g N_VDD_XI10/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI14/MM4 N_XI10/XI14/NET33_XI10/XI14/MM4_d
+ N_XI10/XI14/NET34_XI10/XI14/MM4_g N_VDD_XI10/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI14/MM10 N_XI10/XI14/NET35_XI10/XI14/MM10_d
+ N_XI10/XI14/NET36_XI10/XI14/MM10_g N_VDD_XI10/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI14/MM11 N_XI10/XI14/NET36_XI10/XI14/MM11_d
+ N_XI10/XI14/NET35_XI10/XI14/MM11_g N_VDD_XI10/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI15/MM2 N_XI10/XI15/NET34_XI10/XI15/MM2_d
+ N_XI10/XI15/NET33_XI10/XI15/MM2_g N_VSS_XI10/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI15/MM3 N_XI10/XI15/NET33_XI10/XI15/MM3_d N_WL<16>_XI10/XI15/MM3_g
+ N_BLN<0>_XI10/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI15/MM0 N_XI10/XI15/NET34_XI10/XI15/MM0_d N_WL<16>_XI10/XI15/MM0_g
+ N_BL<0>_XI10/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI15/MM1 N_XI10/XI15/NET33_XI10/XI15/MM1_d
+ N_XI10/XI15/NET34_XI10/XI15/MM1_g N_VSS_XI10/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI15/MM9 N_XI10/XI15/NET36_XI10/XI15/MM9_d N_WL<17>_XI10/XI15/MM9_g
+ N_BL<0>_XI10/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI15/MM6 N_XI10/XI15/NET35_XI10/XI15/MM6_d
+ N_XI10/XI15/NET36_XI10/XI15/MM6_g N_VSS_XI10/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI15/MM7 N_XI10/XI15/NET36_XI10/XI15/MM7_d
+ N_XI10/XI15/NET35_XI10/XI15/MM7_g N_VSS_XI10/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/XI15/MM8 N_XI10/XI15/NET35_XI10/XI15/MM8_d N_WL<17>_XI10/XI15/MM8_g
+ N_BLN<0>_XI10/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI10/XI15/MM5 N_XI10/XI15/NET34_XI10/XI15/MM5_d
+ N_XI10/XI15/NET33_XI10/XI15/MM5_g N_VDD_XI10/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI15/MM4 N_XI10/XI15/NET33_XI10/XI15/MM4_d
+ N_XI10/XI15/NET34_XI10/XI15/MM4_g N_VDD_XI10/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI15/MM10 N_XI10/XI15/NET35_XI10/XI15/MM10_d
+ N_XI10/XI15/NET36_XI10/XI15/MM10_g N_VDD_XI10/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/XI15/MM11 N_XI10/XI15/NET36_XI10/XI15/MM11_d
+ N_XI10/XI15/NET35_XI10/XI15/MM11_g N_VDD_XI10/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI0/MM2 N_XI11/XI0/NET34_XI11/XI0/MM2_d N_XI11/XI0/NET33_XI11/XI0/MM2_g
+ N_VSS_XI11/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI0/MM3 N_XI11/XI0/NET33_XI11/XI0/MM3_d N_WL<18>_XI11/XI0/MM3_g
+ N_BLN<15>_XI11/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI0/MM0 N_XI11/XI0/NET34_XI11/XI0/MM0_d N_WL<18>_XI11/XI0/MM0_g
+ N_BL<15>_XI11/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI0/MM1 N_XI11/XI0/NET33_XI11/XI0/MM1_d N_XI11/XI0/NET34_XI11/XI0/MM1_g
+ N_VSS_XI11/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI0/MM9 N_XI11/XI0/NET36_XI11/XI0/MM9_d N_WL<19>_XI11/XI0/MM9_g
+ N_BL<15>_XI11/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI0/MM6 N_XI11/XI0/NET35_XI11/XI0/MM6_d N_XI11/XI0/NET36_XI11/XI0/MM6_g
+ N_VSS_XI11/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI0/MM7 N_XI11/XI0/NET36_XI11/XI0/MM7_d N_XI11/XI0/NET35_XI11/XI0/MM7_g
+ N_VSS_XI11/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI0/MM8 N_XI11/XI0/NET35_XI11/XI0/MM8_d N_WL<19>_XI11/XI0/MM8_g
+ N_BLN<15>_XI11/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI0/MM5 N_XI11/XI0/NET34_XI11/XI0/MM5_d N_XI11/XI0/NET33_XI11/XI0/MM5_g
+ N_VDD_XI11/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI0/MM4 N_XI11/XI0/NET33_XI11/XI0/MM4_d N_XI11/XI0/NET34_XI11/XI0/MM4_g
+ N_VDD_XI11/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI0/MM10 N_XI11/XI0/NET35_XI11/XI0/MM10_d N_XI11/XI0/NET36_XI11/XI0/MM10_g
+ N_VDD_XI11/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI0/MM11 N_XI11/XI0/NET36_XI11/XI0/MM11_d N_XI11/XI0/NET35_XI11/XI0/MM11_g
+ N_VDD_XI11/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI1/MM2 N_XI11/XI1/NET34_XI11/XI1/MM2_d N_XI11/XI1/NET33_XI11/XI1/MM2_g
+ N_VSS_XI11/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI1/MM3 N_XI11/XI1/NET33_XI11/XI1/MM3_d N_WL<18>_XI11/XI1/MM3_g
+ N_BLN<14>_XI11/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI1/MM0 N_XI11/XI1/NET34_XI11/XI1/MM0_d N_WL<18>_XI11/XI1/MM0_g
+ N_BL<14>_XI11/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI1/MM1 N_XI11/XI1/NET33_XI11/XI1/MM1_d N_XI11/XI1/NET34_XI11/XI1/MM1_g
+ N_VSS_XI11/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI1/MM9 N_XI11/XI1/NET36_XI11/XI1/MM9_d N_WL<19>_XI11/XI1/MM9_g
+ N_BL<14>_XI11/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI1/MM6 N_XI11/XI1/NET35_XI11/XI1/MM6_d N_XI11/XI1/NET36_XI11/XI1/MM6_g
+ N_VSS_XI11/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI1/MM7 N_XI11/XI1/NET36_XI11/XI1/MM7_d N_XI11/XI1/NET35_XI11/XI1/MM7_g
+ N_VSS_XI11/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI1/MM8 N_XI11/XI1/NET35_XI11/XI1/MM8_d N_WL<19>_XI11/XI1/MM8_g
+ N_BLN<14>_XI11/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI1/MM5 N_XI11/XI1/NET34_XI11/XI1/MM5_d N_XI11/XI1/NET33_XI11/XI1/MM5_g
+ N_VDD_XI11/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI1/MM4 N_XI11/XI1/NET33_XI11/XI1/MM4_d N_XI11/XI1/NET34_XI11/XI1/MM4_g
+ N_VDD_XI11/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI1/MM10 N_XI11/XI1/NET35_XI11/XI1/MM10_d N_XI11/XI1/NET36_XI11/XI1/MM10_g
+ N_VDD_XI11/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI1/MM11 N_XI11/XI1/NET36_XI11/XI1/MM11_d N_XI11/XI1/NET35_XI11/XI1/MM11_g
+ N_VDD_XI11/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI2/MM2 N_XI11/XI2/NET34_XI11/XI2/MM2_d N_XI11/XI2/NET33_XI11/XI2/MM2_g
+ N_VSS_XI11/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI2/MM3 N_XI11/XI2/NET33_XI11/XI2/MM3_d N_WL<18>_XI11/XI2/MM3_g
+ N_BLN<13>_XI11/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI2/MM0 N_XI11/XI2/NET34_XI11/XI2/MM0_d N_WL<18>_XI11/XI2/MM0_g
+ N_BL<13>_XI11/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI2/MM1 N_XI11/XI2/NET33_XI11/XI2/MM1_d N_XI11/XI2/NET34_XI11/XI2/MM1_g
+ N_VSS_XI11/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI2/MM9 N_XI11/XI2/NET36_XI11/XI2/MM9_d N_WL<19>_XI11/XI2/MM9_g
+ N_BL<13>_XI11/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI2/MM6 N_XI11/XI2/NET35_XI11/XI2/MM6_d N_XI11/XI2/NET36_XI11/XI2/MM6_g
+ N_VSS_XI11/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI2/MM7 N_XI11/XI2/NET36_XI11/XI2/MM7_d N_XI11/XI2/NET35_XI11/XI2/MM7_g
+ N_VSS_XI11/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI2/MM8 N_XI11/XI2/NET35_XI11/XI2/MM8_d N_WL<19>_XI11/XI2/MM8_g
+ N_BLN<13>_XI11/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI2/MM5 N_XI11/XI2/NET34_XI11/XI2/MM5_d N_XI11/XI2/NET33_XI11/XI2/MM5_g
+ N_VDD_XI11/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI2/MM4 N_XI11/XI2/NET33_XI11/XI2/MM4_d N_XI11/XI2/NET34_XI11/XI2/MM4_g
+ N_VDD_XI11/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI2/MM10 N_XI11/XI2/NET35_XI11/XI2/MM10_d N_XI11/XI2/NET36_XI11/XI2/MM10_g
+ N_VDD_XI11/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI2/MM11 N_XI11/XI2/NET36_XI11/XI2/MM11_d N_XI11/XI2/NET35_XI11/XI2/MM11_g
+ N_VDD_XI11/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI3/MM2 N_XI11/XI3/NET34_XI11/XI3/MM2_d N_XI11/XI3/NET33_XI11/XI3/MM2_g
+ N_VSS_XI11/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI3/MM3 N_XI11/XI3/NET33_XI11/XI3/MM3_d N_WL<18>_XI11/XI3/MM3_g
+ N_BLN<12>_XI11/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI3/MM0 N_XI11/XI3/NET34_XI11/XI3/MM0_d N_WL<18>_XI11/XI3/MM0_g
+ N_BL<12>_XI11/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI3/MM1 N_XI11/XI3/NET33_XI11/XI3/MM1_d N_XI11/XI3/NET34_XI11/XI3/MM1_g
+ N_VSS_XI11/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI3/MM9 N_XI11/XI3/NET36_XI11/XI3/MM9_d N_WL<19>_XI11/XI3/MM9_g
+ N_BL<12>_XI11/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI3/MM6 N_XI11/XI3/NET35_XI11/XI3/MM6_d N_XI11/XI3/NET36_XI11/XI3/MM6_g
+ N_VSS_XI11/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI3/MM7 N_XI11/XI3/NET36_XI11/XI3/MM7_d N_XI11/XI3/NET35_XI11/XI3/MM7_g
+ N_VSS_XI11/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI3/MM8 N_XI11/XI3/NET35_XI11/XI3/MM8_d N_WL<19>_XI11/XI3/MM8_g
+ N_BLN<12>_XI11/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI3/MM5 N_XI11/XI3/NET34_XI11/XI3/MM5_d N_XI11/XI3/NET33_XI11/XI3/MM5_g
+ N_VDD_XI11/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI3/MM4 N_XI11/XI3/NET33_XI11/XI3/MM4_d N_XI11/XI3/NET34_XI11/XI3/MM4_g
+ N_VDD_XI11/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI3/MM10 N_XI11/XI3/NET35_XI11/XI3/MM10_d N_XI11/XI3/NET36_XI11/XI3/MM10_g
+ N_VDD_XI11/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI3/MM11 N_XI11/XI3/NET36_XI11/XI3/MM11_d N_XI11/XI3/NET35_XI11/XI3/MM11_g
+ N_VDD_XI11/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI4/MM2 N_XI11/XI4/NET34_XI11/XI4/MM2_d N_XI11/XI4/NET33_XI11/XI4/MM2_g
+ N_VSS_XI11/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI4/MM3 N_XI11/XI4/NET33_XI11/XI4/MM3_d N_WL<18>_XI11/XI4/MM3_g
+ N_BLN<11>_XI11/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI4/MM0 N_XI11/XI4/NET34_XI11/XI4/MM0_d N_WL<18>_XI11/XI4/MM0_g
+ N_BL<11>_XI11/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI4/MM1 N_XI11/XI4/NET33_XI11/XI4/MM1_d N_XI11/XI4/NET34_XI11/XI4/MM1_g
+ N_VSS_XI11/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI4/MM9 N_XI11/XI4/NET36_XI11/XI4/MM9_d N_WL<19>_XI11/XI4/MM9_g
+ N_BL<11>_XI11/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI4/MM6 N_XI11/XI4/NET35_XI11/XI4/MM6_d N_XI11/XI4/NET36_XI11/XI4/MM6_g
+ N_VSS_XI11/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI4/MM7 N_XI11/XI4/NET36_XI11/XI4/MM7_d N_XI11/XI4/NET35_XI11/XI4/MM7_g
+ N_VSS_XI11/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI4/MM8 N_XI11/XI4/NET35_XI11/XI4/MM8_d N_WL<19>_XI11/XI4/MM8_g
+ N_BLN<11>_XI11/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI4/MM5 N_XI11/XI4/NET34_XI11/XI4/MM5_d N_XI11/XI4/NET33_XI11/XI4/MM5_g
+ N_VDD_XI11/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI4/MM4 N_XI11/XI4/NET33_XI11/XI4/MM4_d N_XI11/XI4/NET34_XI11/XI4/MM4_g
+ N_VDD_XI11/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI4/MM10 N_XI11/XI4/NET35_XI11/XI4/MM10_d N_XI11/XI4/NET36_XI11/XI4/MM10_g
+ N_VDD_XI11/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI4/MM11 N_XI11/XI4/NET36_XI11/XI4/MM11_d N_XI11/XI4/NET35_XI11/XI4/MM11_g
+ N_VDD_XI11/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI5/MM2 N_XI11/XI5/NET34_XI11/XI5/MM2_d N_XI11/XI5/NET33_XI11/XI5/MM2_g
+ N_VSS_XI11/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI5/MM3 N_XI11/XI5/NET33_XI11/XI5/MM3_d N_WL<18>_XI11/XI5/MM3_g
+ N_BLN<10>_XI11/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI5/MM0 N_XI11/XI5/NET34_XI11/XI5/MM0_d N_WL<18>_XI11/XI5/MM0_g
+ N_BL<10>_XI11/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI5/MM1 N_XI11/XI5/NET33_XI11/XI5/MM1_d N_XI11/XI5/NET34_XI11/XI5/MM1_g
+ N_VSS_XI11/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI5/MM9 N_XI11/XI5/NET36_XI11/XI5/MM9_d N_WL<19>_XI11/XI5/MM9_g
+ N_BL<10>_XI11/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI5/MM6 N_XI11/XI5/NET35_XI11/XI5/MM6_d N_XI11/XI5/NET36_XI11/XI5/MM6_g
+ N_VSS_XI11/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI5/MM7 N_XI11/XI5/NET36_XI11/XI5/MM7_d N_XI11/XI5/NET35_XI11/XI5/MM7_g
+ N_VSS_XI11/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI5/MM8 N_XI11/XI5/NET35_XI11/XI5/MM8_d N_WL<19>_XI11/XI5/MM8_g
+ N_BLN<10>_XI11/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI5/MM5 N_XI11/XI5/NET34_XI11/XI5/MM5_d N_XI11/XI5/NET33_XI11/XI5/MM5_g
+ N_VDD_XI11/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI5/MM4 N_XI11/XI5/NET33_XI11/XI5/MM4_d N_XI11/XI5/NET34_XI11/XI5/MM4_g
+ N_VDD_XI11/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI5/MM10 N_XI11/XI5/NET35_XI11/XI5/MM10_d N_XI11/XI5/NET36_XI11/XI5/MM10_g
+ N_VDD_XI11/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI5/MM11 N_XI11/XI5/NET36_XI11/XI5/MM11_d N_XI11/XI5/NET35_XI11/XI5/MM11_g
+ N_VDD_XI11/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI6/MM2 N_XI11/XI6/NET34_XI11/XI6/MM2_d N_XI11/XI6/NET33_XI11/XI6/MM2_g
+ N_VSS_XI11/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM3 N_XI11/XI6/NET33_XI11/XI6/MM3_d N_WL<18>_XI11/XI6/MM3_g
+ N_BLN<9>_XI11/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM0 N_XI11/XI6/NET34_XI11/XI6/MM0_d N_WL<18>_XI11/XI6/MM0_g
+ N_BL<9>_XI11/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM1 N_XI11/XI6/NET33_XI11/XI6/MM1_d N_XI11/XI6/NET34_XI11/XI6/MM1_g
+ N_VSS_XI11/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM9 N_XI11/XI6/NET36_XI11/XI6/MM9_d N_WL<19>_XI11/XI6/MM9_g
+ N_BL<9>_XI11/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM6 N_XI11/XI6/NET35_XI11/XI6/MM6_d N_XI11/XI6/NET36_XI11/XI6/MM6_g
+ N_VSS_XI11/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM7 N_XI11/XI6/NET36_XI11/XI6/MM7_d N_XI11/XI6/NET35_XI11/XI6/MM7_g
+ N_VSS_XI11/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM8 N_XI11/XI6/NET35_XI11/XI6/MM8_d N_WL<19>_XI11/XI6/MM8_g
+ N_BLN<9>_XI11/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI6/MM5 N_XI11/XI6/NET34_XI11/XI6/MM5_d N_XI11/XI6/NET33_XI11/XI6/MM5_g
+ N_VDD_XI11/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI6/MM4 N_XI11/XI6/NET33_XI11/XI6/MM4_d N_XI11/XI6/NET34_XI11/XI6/MM4_g
+ N_VDD_XI11/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI6/MM10 N_XI11/XI6/NET35_XI11/XI6/MM10_d N_XI11/XI6/NET36_XI11/XI6/MM10_g
+ N_VDD_XI11/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI6/MM11 N_XI11/XI6/NET36_XI11/XI6/MM11_d N_XI11/XI6/NET35_XI11/XI6/MM11_g
+ N_VDD_XI11/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI7/MM2 N_XI11/XI7/NET34_XI11/XI7/MM2_d N_XI11/XI7/NET33_XI11/XI7/MM2_g
+ N_VSS_XI11/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM3 N_XI11/XI7/NET33_XI11/XI7/MM3_d N_WL<18>_XI11/XI7/MM3_g
+ N_BLN<8>_XI11/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM0 N_XI11/XI7/NET34_XI11/XI7/MM0_d N_WL<18>_XI11/XI7/MM0_g
+ N_BL<8>_XI11/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM1 N_XI11/XI7/NET33_XI11/XI7/MM1_d N_XI11/XI7/NET34_XI11/XI7/MM1_g
+ N_VSS_XI11/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM9 N_XI11/XI7/NET36_XI11/XI7/MM9_d N_WL<19>_XI11/XI7/MM9_g
+ N_BL<8>_XI11/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM6 N_XI11/XI7/NET35_XI11/XI7/MM6_d N_XI11/XI7/NET36_XI11/XI7/MM6_g
+ N_VSS_XI11/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM7 N_XI11/XI7/NET36_XI11/XI7/MM7_d N_XI11/XI7/NET35_XI11/XI7/MM7_g
+ N_VSS_XI11/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM8 N_XI11/XI7/NET35_XI11/XI7/MM8_d N_WL<19>_XI11/XI7/MM8_g
+ N_BLN<8>_XI11/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI7/MM5 N_XI11/XI7/NET34_XI11/XI7/MM5_d N_XI11/XI7/NET33_XI11/XI7/MM5_g
+ N_VDD_XI11/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI7/MM4 N_XI11/XI7/NET33_XI11/XI7/MM4_d N_XI11/XI7/NET34_XI11/XI7/MM4_g
+ N_VDD_XI11/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI7/MM10 N_XI11/XI7/NET35_XI11/XI7/MM10_d N_XI11/XI7/NET36_XI11/XI7/MM10_g
+ N_VDD_XI11/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI7/MM11 N_XI11/XI7/NET36_XI11/XI7/MM11_d N_XI11/XI7/NET35_XI11/XI7/MM11_g
+ N_VDD_XI11/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI8/MM2 N_XI11/XI8/NET34_XI11/XI8/MM2_d N_XI11/XI8/NET33_XI11/XI8/MM2_g
+ N_VSS_XI11/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM3 N_XI11/XI8/NET33_XI11/XI8/MM3_d N_WL<18>_XI11/XI8/MM3_g
+ N_BLN<7>_XI11/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM0 N_XI11/XI8/NET34_XI11/XI8/MM0_d N_WL<18>_XI11/XI8/MM0_g
+ N_BL<7>_XI11/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM1 N_XI11/XI8/NET33_XI11/XI8/MM1_d N_XI11/XI8/NET34_XI11/XI8/MM1_g
+ N_VSS_XI11/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM9 N_XI11/XI8/NET36_XI11/XI8/MM9_d N_WL<19>_XI11/XI8/MM9_g
+ N_BL<7>_XI11/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM6 N_XI11/XI8/NET35_XI11/XI8/MM6_d N_XI11/XI8/NET36_XI11/XI8/MM6_g
+ N_VSS_XI11/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM7 N_XI11/XI8/NET36_XI11/XI8/MM7_d N_XI11/XI8/NET35_XI11/XI8/MM7_g
+ N_VSS_XI11/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM8 N_XI11/XI8/NET35_XI11/XI8/MM8_d N_WL<19>_XI11/XI8/MM8_g
+ N_BLN<7>_XI11/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI8/MM5 N_XI11/XI8/NET34_XI11/XI8/MM5_d N_XI11/XI8/NET33_XI11/XI8/MM5_g
+ N_VDD_XI11/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI8/MM4 N_XI11/XI8/NET33_XI11/XI8/MM4_d N_XI11/XI8/NET34_XI11/XI8/MM4_g
+ N_VDD_XI11/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI8/MM10 N_XI11/XI8/NET35_XI11/XI8/MM10_d N_XI11/XI8/NET36_XI11/XI8/MM10_g
+ N_VDD_XI11/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI8/MM11 N_XI11/XI8/NET36_XI11/XI8/MM11_d N_XI11/XI8/NET35_XI11/XI8/MM11_g
+ N_VDD_XI11/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI9/MM2 N_XI11/XI9/NET34_XI11/XI9/MM2_d N_XI11/XI9/NET33_XI11/XI9/MM2_g
+ N_VSS_XI11/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM3 N_XI11/XI9/NET33_XI11/XI9/MM3_d N_WL<18>_XI11/XI9/MM3_g
+ N_BLN<6>_XI11/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM0 N_XI11/XI9/NET34_XI11/XI9/MM0_d N_WL<18>_XI11/XI9/MM0_g
+ N_BL<6>_XI11/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM1 N_XI11/XI9/NET33_XI11/XI9/MM1_d N_XI11/XI9/NET34_XI11/XI9/MM1_g
+ N_VSS_XI11/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM9 N_XI11/XI9/NET36_XI11/XI9/MM9_d N_WL<19>_XI11/XI9/MM9_g
+ N_BL<6>_XI11/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM6 N_XI11/XI9/NET35_XI11/XI9/MM6_d N_XI11/XI9/NET36_XI11/XI9/MM6_g
+ N_VSS_XI11/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM7 N_XI11/XI9/NET36_XI11/XI9/MM7_d N_XI11/XI9/NET35_XI11/XI9/MM7_g
+ N_VSS_XI11/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM8 N_XI11/XI9/NET35_XI11/XI9/MM8_d N_WL<19>_XI11/XI9/MM8_g
+ N_BLN<6>_XI11/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI9/MM5 N_XI11/XI9/NET34_XI11/XI9/MM5_d N_XI11/XI9/NET33_XI11/XI9/MM5_g
+ N_VDD_XI11/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI9/MM4 N_XI11/XI9/NET33_XI11/XI9/MM4_d N_XI11/XI9/NET34_XI11/XI9/MM4_g
+ N_VDD_XI11/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI9/MM10 N_XI11/XI9/NET35_XI11/XI9/MM10_d N_XI11/XI9/NET36_XI11/XI9/MM10_g
+ N_VDD_XI11/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI9/MM11 N_XI11/XI9/NET36_XI11/XI9/MM11_d N_XI11/XI9/NET35_XI11/XI9/MM11_g
+ N_VDD_XI11/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI10/MM2 N_XI11/XI10/NET34_XI11/XI10/MM2_d
+ N_XI11/XI10/NET33_XI11/XI10/MM2_g N_VSS_XI11/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI10/MM3 N_XI11/XI10/NET33_XI11/XI10/MM3_d N_WL<18>_XI11/XI10/MM3_g
+ N_BLN<5>_XI11/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI10/MM0 N_XI11/XI10/NET34_XI11/XI10/MM0_d N_WL<18>_XI11/XI10/MM0_g
+ N_BL<5>_XI11/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI10/MM1 N_XI11/XI10/NET33_XI11/XI10/MM1_d
+ N_XI11/XI10/NET34_XI11/XI10/MM1_g N_VSS_XI11/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI10/MM9 N_XI11/XI10/NET36_XI11/XI10/MM9_d N_WL<19>_XI11/XI10/MM9_g
+ N_BL<5>_XI11/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI10/MM6 N_XI11/XI10/NET35_XI11/XI10/MM6_d
+ N_XI11/XI10/NET36_XI11/XI10/MM6_g N_VSS_XI11/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI10/MM7 N_XI11/XI10/NET36_XI11/XI10/MM7_d
+ N_XI11/XI10/NET35_XI11/XI10/MM7_g N_VSS_XI11/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI10/MM8 N_XI11/XI10/NET35_XI11/XI10/MM8_d N_WL<19>_XI11/XI10/MM8_g
+ N_BLN<5>_XI11/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI10/MM5 N_XI11/XI10/NET34_XI11/XI10/MM5_d
+ N_XI11/XI10/NET33_XI11/XI10/MM5_g N_VDD_XI11/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI10/MM4 N_XI11/XI10/NET33_XI11/XI10/MM4_d
+ N_XI11/XI10/NET34_XI11/XI10/MM4_g N_VDD_XI11/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI10/MM10 N_XI11/XI10/NET35_XI11/XI10/MM10_d
+ N_XI11/XI10/NET36_XI11/XI10/MM10_g N_VDD_XI11/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI10/MM11 N_XI11/XI10/NET36_XI11/XI10/MM11_d
+ N_XI11/XI10/NET35_XI11/XI10/MM11_g N_VDD_XI11/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI11/MM2 N_XI11/XI11/NET34_XI11/XI11/MM2_d
+ N_XI11/XI11/NET33_XI11/XI11/MM2_g N_VSS_XI11/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI11/MM3 N_XI11/XI11/NET33_XI11/XI11/MM3_d N_WL<18>_XI11/XI11/MM3_g
+ N_BLN<4>_XI11/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI11/MM0 N_XI11/XI11/NET34_XI11/XI11/MM0_d N_WL<18>_XI11/XI11/MM0_g
+ N_BL<4>_XI11/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI11/MM1 N_XI11/XI11/NET33_XI11/XI11/MM1_d
+ N_XI11/XI11/NET34_XI11/XI11/MM1_g N_VSS_XI11/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI11/MM9 N_XI11/XI11/NET36_XI11/XI11/MM9_d N_WL<19>_XI11/XI11/MM9_g
+ N_BL<4>_XI11/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI11/MM6 N_XI11/XI11/NET35_XI11/XI11/MM6_d
+ N_XI11/XI11/NET36_XI11/XI11/MM6_g N_VSS_XI11/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI11/MM7 N_XI11/XI11/NET36_XI11/XI11/MM7_d
+ N_XI11/XI11/NET35_XI11/XI11/MM7_g N_VSS_XI11/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI11/MM8 N_XI11/XI11/NET35_XI11/XI11/MM8_d N_WL<19>_XI11/XI11/MM8_g
+ N_BLN<4>_XI11/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI11/MM5 N_XI11/XI11/NET34_XI11/XI11/MM5_d
+ N_XI11/XI11/NET33_XI11/XI11/MM5_g N_VDD_XI11/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI11/MM4 N_XI11/XI11/NET33_XI11/XI11/MM4_d
+ N_XI11/XI11/NET34_XI11/XI11/MM4_g N_VDD_XI11/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI11/MM10 N_XI11/XI11/NET35_XI11/XI11/MM10_d
+ N_XI11/XI11/NET36_XI11/XI11/MM10_g N_VDD_XI11/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI11/MM11 N_XI11/XI11/NET36_XI11/XI11/MM11_d
+ N_XI11/XI11/NET35_XI11/XI11/MM11_g N_VDD_XI11/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI12/MM2 N_XI11/XI12/NET34_XI11/XI12/MM2_d
+ N_XI11/XI12/NET33_XI11/XI12/MM2_g N_VSS_XI11/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI12/MM3 N_XI11/XI12/NET33_XI11/XI12/MM3_d N_WL<18>_XI11/XI12/MM3_g
+ N_BLN<3>_XI11/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI12/MM0 N_XI11/XI12/NET34_XI11/XI12/MM0_d N_WL<18>_XI11/XI12/MM0_g
+ N_BL<3>_XI11/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI12/MM1 N_XI11/XI12/NET33_XI11/XI12/MM1_d
+ N_XI11/XI12/NET34_XI11/XI12/MM1_g N_VSS_XI11/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI12/MM9 N_XI11/XI12/NET36_XI11/XI12/MM9_d N_WL<19>_XI11/XI12/MM9_g
+ N_BL<3>_XI11/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI12/MM6 N_XI11/XI12/NET35_XI11/XI12/MM6_d
+ N_XI11/XI12/NET36_XI11/XI12/MM6_g N_VSS_XI11/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI12/MM7 N_XI11/XI12/NET36_XI11/XI12/MM7_d
+ N_XI11/XI12/NET35_XI11/XI12/MM7_g N_VSS_XI11/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI12/MM8 N_XI11/XI12/NET35_XI11/XI12/MM8_d N_WL<19>_XI11/XI12/MM8_g
+ N_BLN<3>_XI11/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI12/MM5 N_XI11/XI12/NET34_XI11/XI12/MM5_d
+ N_XI11/XI12/NET33_XI11/XI12/MM5_g N_VDD_XI11/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI12/MM4 N_XI11/XI12/NET33_XI11/XI12/MM4_d
+ N_XI11/XI12/NET34_XI11/XI12/MM4_g N_VDD_XI11/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI12/MM10 N_XI11/XI12/NET35_XI11/XI12/MM10_d
+ N_XI11/XI12/NET36_XI11/XI12/MM10_g N_VDD_XI11/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI12/MM11 N_XI11/XI12/NET36_XI11/XI12/MM11_d
+ N_XI11/XI12/NET35_XI11/XI12/MM11_g N_VDD_XI11/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI13/MM2 N_XI11/XI13/NET34_XI11/XI13/MM2_d
+ N_XI11/XI13/NET33_XI11/XI13/MM2_g N_VSS_XI11/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI13/MM3 N_XI11/XI13/NET33_XI11/XI13/MM3_d N_WL<18>_XI11/XI13/MM3_g
+ N_BLN<2>_XI11/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI13/MM0 N_XI11/XI13/NET34_XI11/XI13/MM0_d N_WL<18>_XI11/XI13/MM0_g
+ N_BL<2>_XI11/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI13/MM1 N_XI11/XI13/NET33_XI11/XI13/MM1_d
+ N_XI11/XI13/NET34_XI11/XI13/MM1_g N_VSS_XI11/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI13/MM9 N_XI11/XI13/NET36_XI11/XI13/MM9_d N_WL<19>_XI11/XI13/MM9_g
+ N_BL<2>_XI11/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI13/MM6 N_XI11/XI13/NET35_XI11/XI13/MM6_d
+ N_XI11/XI13/NET36_XI11/XI13/MM6_g N_VSS_XI11/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI13/MM7 N_XI11/XI13/NET36_XI11/XI13/MM7_d
+ N_XI11/XI13/NET35_XI11/XI13/MM7_g N_VSS_XI11/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI13/MM8 N_XI11/XI13/NET35_XI11/XI13/MM8_d N_WL<19>_XI11/XI13/MM8_g
+ N_BLN<2>_XI11/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI13/MM5 N_XI11/XI13/NET34_XI11/XI13/MM5_d
+ N_XI11/XI13/NET33_XI11/XI13/MM5_g N_VDD_XI11/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI13/MM4 N_XI11/XI13/NET33_XI11/XI13/MM4_d
+ N_XI11/XI13/NET34_XI11/XI13/MM4_g N_VDD_XI11/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI13/MM10 N_XI11/XI13/NET35_XI11/XI13/MM10_d
+ N_XI11/XI13/NET36_XI11/XI13/MM10_g N_VDD_XI11/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI13/MM11 N_XI11/XI13/NET36_XI11/XI13/MM11_d
+ N_XI11/XI13/NET35_XI11/XI13/MM11_g N_VDD_XI11/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI14/MM2 N_XI11/XI14/NET34_XI11/XI14/MM2_d
+ N_XI11/XI14/NET33_XI11/XI14/MM2_g N_VSS_XI11/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI14/MM3 N_XI11/XI14/NET33_XI11/XI14/MM3_d N_WL<18>_XI11/XI14/MM3_g
+ N_BLN<1>_XI11/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI14/MM0 N_XI11/XI14/NET34_XI11/XI14/MM0_d N_WL<18>_XI11/XI14/MM0_g
+ N_BL<1>_XI11/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI14/MM1 N_XI11/XI14/NET33_XI11/XI14/MM1_d
+ N_XI11/XI14/NET34_XI11/XI14/MM1_g N_VSS_XI11/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI14/MM9 N_XI11/XI14/NET36_XI11/XI14/MM9_d N_WL<19>_XI11/XI14/MM9_g
+ N_BL<1>_XI11/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI14/MM6 N_XI11/XI14/NET35_XI11/XI14/MM6_d
+ N_XI11/XI14/NET36_XI11/XI14/MM6_g N_VSS_XI11/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI14/MM7 N_XI11/XI14/NET36_XI11/XI14/MM7_d
+ N_XI11/XI14/NET35_XI11/XI14/MM7_g N_VSS_XI11/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI14/MM8 N_XI11/XI14/NET35_XI11/XI14/MM8_d N_WL<19>_XI11/XI14/MM8_g
+ N_BLN<1>_XI11/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI14/MM5 N_XI11/XI14/NET34_XI11/XI14/MM5_d
+ N_XI11/XI14/NET33_XI11/XI14/MM5_g N_VDD_XI11/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI14/MM4 N_XI11/XI14/NET33_XI11/XI14/MM4_d
+ N_XI11/XI14/NET34_XI11/XI14/MM4_g N_VDD_XI11/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI14/MM10 N_XI11/XI14/NET35_XI11/XI14/MM10_d
+ N_XI11/XI14/NET36_XI11/XI14/MM10_g N_VDD_XI11/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI14/MM11 N_XI11/XI14/NET36_XI11/XI14/MM11_d
+ N_XI11/XI14/NET35_XI11/XI14/MM11_g N_VDD_XI11/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI15/MM2 N_XI11/XI15/NET34_XI11/XI15/MM2_d
+ N_XI11/XI15/NET33_XI11/XI15/MM2_g N_VSS_XI11/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI15/MM3 N_XI11/XI15/NET33_XI11/XI15/MM3_d N_WL<18>_XI11/XI15/MM3_g
+ N_BLN<0>_XI11/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI15/MM0 N_XI11/XI15/NET34_XI11/XI15/MM0_d N_WL<18>_XI11/XI15/MM0_g
+ N_BL<0>_XI11/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI15/MM1 N_XI11/XI15/NET33_XI11/XI15/MM1_d
+ N_XI11/XI15/NET34_XI11/XI15/MM1_g N_VSS_XI11/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI15/MM9 N_XI11/XI15/NET36_XI11/XI15/MM9_d N_WL<19>_XI11/XI15/MM9_g
+ N_BL<0>_XI11/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI15/MM6 N_XI11/XI15/NET35_XI11/XI15/MM6_d
+ N_XI11/XI15/NET36_XI11/XI15/MM6_g N_VSS_XI11/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI15/MM7 N_XI11/XI15/NET36_XI11/XI15/MM7_d
+ N_XI11/XI15/NET35_XI11/XI15/MM7_g N_VSS_XI11/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/XI15/MM8 N_XI11/XI15/NET35_XI11/XI15/MM8_d N_WL<19>_XI11/XI15/MM8_g
+ N_BLN<0>_XI11/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI11/XI15/MM5 N_XI11/XI15/NET34_XI11/XI15/MM5_d
+ N_XI11/XI15/NET33_XI11/XI15/MM5_g N_VDD_XI11/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI15/MM4 N_XI11/XI15/NET33_XI11/XI15/MM4_d
+ N_XI11/XI15/NET34_XI11/XI15/MM4_g N_VDD_XI11/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI15/MM10 N_XI11/XI15/NET35_XI11/XI15/MM10_d
+ N_XI11/XI15/NET36_XI11/XI15/MM10_g N_VDD_XI11/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/XI15/MM11 N_XI11/XI15/NET36_XI11/XI15/MM11_d
+ N_XI11/XI15/NET35_XI11/XI15/MM11_g N_VDD_XI11/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI0/MM2 N_XI12/XI0/NET34_XI12/XI0/MM2_d N_XI12/XI0/NET33_XI12/XI0/MM2_g
+ N_VSS_XI12/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI0/MM3 N_XI12/XI0/NET33_XI12/XI0/MM3_d N_WL<20>_XI12/XI0/MM3_g
+ N_BLN<15>_XI12/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI0/MM0 N_XI12/XI0/NET34_XI12/XI0/MM0_d N_WL<20>_XI12/XI0/MM0_g
+ N_BL<15>_XI12/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI0/MM1 N_XI12/XI0/NET33_XI12/XI0/MM1_d N_XI12/XI0/NET34_XI12/XI0/MM1_g
+ N_VSS_XI12/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI0/MM9 N_XI12/XI0/NET36_XI12/XI0/MM9_d N_WL<21>_XI12/XI0/MM9_g
+ N_BL<15>_XI12/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI0/MM6 N_XI12/XI0/NET35_XI12/XI0/MM6_d N_XI12/XI0/NET36_XI12/XI0/MM6_g
+ N_VSS_XI12/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI0/MM7 N_XI12/XI0/NET36_XI12/XI0/MM7_d N_XI12/XI0/NET35_XI12/XI0/MM7_g
+ N_VSS_XI12/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI0/MM8 N_XI12/XI0/NET35_XI12/XI0/MM8_d N_WL<21>_XI12/XI0/MM8_g
+ N_BLN<15>_XI12/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI0/MM5 N_XI12/XI0/NET34_XI12/XI0/MM5_d N_XI12/XI0/NET33_XI12/XI0/MM5_g
+ N_VDD_XI12/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI0/MM4 N_XI12/XI0/NET33_XI12/XI0/MM4_d N_XI12/XI0/NET34_XI12/XI0/MM4_g
+ N_VDD_XI12/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI0/MM10 N_XI12/XI0/NET35_XI12/XI0/MM10_d N_XI12/XI0/NET36_XI12/XI0/MM10_g
+ N_VDD_XI12/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI0/MM11 N_XI12/XI0/NET36_XI12/XI0/MM11_d N_XI12/XI0/NET35_XI12/XI0/MM11_g
+ N_VDD_XI12/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI1/MM2 N_XI12/XI1/NET34_XI12/XI1/MM2_d N_XI12/XI1/NET33_XI12/XI1/MM2_g
+ N_VSS_XI12/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI1/MM3 N_XI12/XI1/NET33_XI12/XI1/MM3_d N_WL<20>_XI12/XI1/MM3_g
+ N_BLN<14>_XI12/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI1/MM0 N_XI12/XI1/NET34_XI12/XI1/MM0_d N_WL<20>_XI12/XI1/MM0_g
+ N_BL<14>_XI12/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI1/MM1 N_XI12/XI1/NET33_XI12/XI1/MM1_d N_XI12/XI1/NET34_XI12/XI1/MM1_g
+ N_VSS_XI12/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI1/MM9 N_XI12/XI1/NET36_XI12/XI1/MM9_d N_WL<21>_XI12/XI1/MM9_g
+ N_BL<14>_XI12/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI1/MM6 N_XI12/XI1/NET35_XI12/XI1/MM6_d N_XI12/XI1/NET36_XI12/XI1/MM6_g
+ N_VSS_XI12/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI1/MM7 N_XI12/XI1/NET36_XI12/XI1/MM7_d N_XI12/XI1/NET35_XI12/XI1/MM7_g
+ N_VSS_XI12/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI1/MM8 N_XI12/XI1/NET35_XI12/XI1/MM8_d N_WL<21>_XI12/XI1/MM8_g
+ N_BLN<14>_XI12/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI1/MM5 N_XI12/XI1/NET34_XI12/XI1/MM5_d N_XI12/XI1/NET33_XI12/XI1/MM5_g
+ N_VDD_XI12/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI1/MM4 N_XI12/XI1/NET33_XI12/XI1/MM4_d N_XI12/XI1/NET34_XI12/XI1/MM4_g
+ N_VDD_XI12/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI1/MM10 N_XI12/XI1/NET35_XI12/XI1/MM10_d N_XI12/XI1/NET36_XI12/XI1/MM10_g
+ N_VDD_XI12/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI1/MM11 N_XI12/XI1/NET36_XI12/XI1/MM11_d N_XI12/XI1/NET35_XI12/XI1/MM11_g
+ N_VDD_XI12/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI2/MM2 N_XI12/XI2/NET34_XI12/XI2/MM2_d N_XI12/XI2/NET33_XI12/XI2/MM2_g
+ N_VSS_XI12/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI2/MM3 N_XI12/XI2/NET33_XI12/XI2/MM3_d N_WL<20>_XI12/XI2/MM3_g
+ N_BLN<13>_XI12/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI2/MM0 N_XI12/XI2/NET34_XI12/XI2/MM0_d N_WL<20>_XI12/XI2/MM0_g
+ N_BL<13>_XI12/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI2/MM1 N_XI12/XI2/NET33_XI12/XI2/MM1_d N_XI12/XI2/NET34_XI12/XI2/MM1_g
+ N_VSS_XI12/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI2/MM9 N_XI12/XI2/NET36_XI12/XI2/MM9_d N_WL<21>_XI12/XI2/MM9_g
+ N_BL<13>_XI12/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI2/MM6 N_XI12/XI2/NET35_XI12/XI2/MM6_d N_XI12/XI2/NET36_XI12/XI2/MM6_g
+ N_VSS_XI12/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI2/MM7 N_XI12/XI2/NET36_XI12/XI2/MM7_d N_XI12/XI2/NET35_XI12/XI2/MM7_g
+ N_VSS_XI12/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI2/MM8 N_XI12/XI2/NET35_XI12/XI2/MM8_d N_WL<21>_XI12/XI2/MM8_g
+ N_BLN<13>_XI12/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI2/MM5 N_XI12/XI2/NET34_XI12/XI2/MM5_d N_XI12/XI2/NET33_XI12/XI2/MM5_g
+ N_VDD_XI12/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI2/MM4 N_XI12/XI2/NET33_XI12/XI2/MM4_d N_XI12/XI2/NET34_XI12/XI2/MM4_g
+ N_VDD_XI12/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI2/MM10 N_XI12/XI2/NET35_XI12/XI2/MM10_d N_XI12/XI2/NET36_XI12/XI2/MM10_g
+ N_VDD_XI12/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI2/MM11 N_XI12/XI2/NET36_XI12/XI2/MM11_d N_XI12/XI2/NET35_XI12/XI2/MM11_g
+ N_VDD_XI12/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI3/MM2 N_XI12/XI3/NET34_XI12/XI3/MM2_d N_XI12/XI3/NET33_XI12/XI3/MM2_g
+ N_VSS_XI12/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI3/MM3 N_XI12/XI3/NET33_XI12/XI3/MM3_d N_WL<20>_XI12/XI3/MM3_g
+ N_BLN<12>_XI12/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI3/MM0 N_XI12/XI3/NET34_XI12/XI3/MM0_d N_WL<20>_XI12/XI3/MM0_g
+ N_BL<12>_XI12/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI3/MM1 N_XI12/XI3/NET33_XI12/XI3/MM1_d N_XI12/XI3/NET34_XI12/XI3/MM1_g
+ N_VSS_XI12/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI3/MM9 N_XI12/XI3/NET36_XI12/XI3/MM9_d N_WL<21>_XI12/XI3/MM9_g
+ N_BL<12>_XI12/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI3/MM6 N_XI12/XI3/NET35_XI12/XI3/MM6_d N_XI12/XI3/NET36_XI12/XI3/MM6_g
+ N_VSS_XI12/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI3/MM7 N_XI12/XI3/NET36_XI12/XI3/MM7_d N_XI12/XI3/NET35_XI12/XI3/MM7_g
+ N_VSS_XI12/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI3/MM8 N_XI12/XI3/NET35_XI12/XI3/MM8_d N_WL<21>_XI12/XI3/MM8_g
+ N_BLN<12>_XI12/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI3/MM5 N_XI12/XI3/NET34_XI12/XI3/MM5_d N_XI12/XI3/NET33_XI12/XI3/MM5_g
+ N_VDD_XI12/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI3/MM4 N_XI12/XI3/NET33_XI12/XI3/MM4_d N_XI12/XI3/NET34_XI12/XI3/MM4_g
+ N_VDD_XI12/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI3/MM10 N_XI12/XI3/NET35_XI12/XI3/MM10_d N_XI12/XI3/NET36_XI12/XI3/MM10_g
+ N_VDD_XI12/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI3/MM11 N_XI12/XI3/NET36_XI12/XI3/MM11_d N_XI12/XI3/NET35_XI12/XI3/MM11_g
+ N_VDD_XI12/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI4/MM2 N_XI12/XI4/NET34_XI12/XI4/MM2_d N_XI12/XI4/NET33_XI12/XI4/MM2_g
+ N_VSS_XI12/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI4/MM3 N_XI12/XI4/NET33_XI12/XI4/MM3_d N_WL<20>_XI12/XI4/MM3_g
+ N_BLN<11>_XI12/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI4/MM0 N_XI12/XI4/NET34_XI12/XI4/MM0_d N_WL<20>_XI12/XI4/MM0_g
+ N_BL<11>_XI12/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI4/MM1 N_XI12/XI4/NET33_XI12/XI4/MM1_d N_XI12/XI4/NET34_XI12/XI4/MM1_g
+ N_VSS_XI12/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI4/MM9 N_XI12/XI4/NET36_XI12/XI4/MM9_d N_WL<21>_XI12/XI4/MM9_g
+ N_BL<11>_XI12/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI4/MM6 N_XI12/XI4/NET35_XI12/XI4/MM6_d N_XI12/XI4/NET36_XI12/XI4/MM6_g
+ N_VSS_XI12/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI4/MM7 N_XI12/XI4/NET36_XI12/XI4/MM7_d N_XI12/XI4/NET35_XI12/XI4/MM7_g
+ N_VSS_XI12/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI4/MM8 N_XI12/XI4/NET35_XI12/XI4/MM8_d N_WL<21>_XI12/XI4/MM8_g
+ N_BLN<11>_XI12/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI4/MM5 N_XI12/XI4/NET34_XI12/XI4/MM5_d N_XI12/XI4/NET33_XI12/XI4/MM5_g
+ N_VDD_XI12/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI4/MM4 N_XI12/XI4/NET33_XI12/XI4/MM4_d N_XI12/XI4/NET34_XI12/XI4/MM4_g
+ N_VDD_XI12/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI4/MM10 N_XI12/XI4/NET35_XI12/XI4/MM10_d N_XI12/XI4/NET36_XI12/XI4/MM10_g
+ N_VDD_XI12/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI4/MM11 N_XI12/XI4/NET36_XI12/XI4/MM11_d N_XI12/XI4/NET35_XI12/XI4/MM11_g
+ N_VDD_XI12/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI5/MM2 N_XI12/XI5/NET34_XI12/XI5/MM2_d N_XI12/XI5/NET33_XI12/XI5/MM2_g
+ N_VSS_XI12/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI5/MM3 N_XI12/XI5/NET33_XI12/XI5/MM3_d N_WL<20>_XI12/XI5/MM3_g
+ N_BLN<10>_XI12/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI5/MM0 N_XI12/XI5/NET34_XI12/XI5/MM0_d N_WL<20>_XI12/XI5/MM0_g
+ N_BL<10>_XI12/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI5/MM1 N_XI12/XI5/NET33_XI12/XI5/MM1_d N_XI12/XI5/NET34_XI12/XI5/MM1_g
+ N_VSS_XI12/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI5/MM9 N_XI12/XI5/NET36_XI12/XI5/MM9_d N_WL<21>_XI12/XI5/MM9_g
+ N_BL<10>_XI12/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI5/MM6 N_XI12/XI5/NET35_XI12/XI5/MM6_d N_XI12/XI5/NET36_XI12/XI5/MM6_g
+ N_VSS_XI12/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI5/MM7 N_XI12/XI5/NET36_XI12/XI5/MM7_d N_XI12/XI5/NET35_XI12/XI5/MM7_g
+ N_VSS_XI12/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI5/MM8 N_XI12/XI5/NET35_XI12/XI5/MM8_d N_WL<21>_XI12/XI5/MM8_g
+ N_BLN<10>_XI12/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI5/MM5 N_XI12/XI5/NET34_XI12/XI5/MM5_d N_XI12/XI5/NET33_XI12/XI5/MM5_g
+ N_VDD_XI12/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI5/MM4 N_XI12/XI5/NET33_XI12/XI5/MM4_d N_XI12/XI5/NET34_XI12/XI5/MM4_g
+ N_VDD_XI12/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI5/MM10 N_XI12/XI5/NET35_XI12/XI5/MM10_d N_XI12/XI5/NET36_XI12/XI5/MM10_g
+ N_VDD_XI12/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI5/MM11 N_XI12/XI5/NET36_XI12/XI5/MM11_d N_XI12/XI5/NET35_XI12/XI5/MM11_g
+ N_VDD_XI12/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI6/MM2 N_XI12/XI6/NET34_XI12/XI6/MM2_d N_XI12/XI6/NET33_XI12/XI6/MM2_g
+ N_VSS_XI12/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM3 N_XI12/XI6/NET33_XI12/XI6/MM3_d N_WL<20>_XI12/XI6/MM3_g
+ N_BLN<9>_XI12/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM0 N_XI12/XI6/NET34_XI12/XI6/MM0_d N_WL<20>_XI12/XI6/MM0_g
+ N_BL<9>_XI12/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM1 N_XI12/XI6/NET33_XI12/XI6/MM1_d N_XI12/XI6/NET34_XI12/XI6/MM1_g
+ N_VSS_XI12/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM9 N_XI12/XI6/NET36_XI12/XI6/MM9_d N_WL<21>_XI12/XI6/MM9_g
+ N_BL<9>_XI12/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM6 N_XI12/XI6/NET35_XI12/XI6/MM6_d N_XI12/XI6/NET36_XI12/XI6/MM6_g
+ N_VSS_XI12/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM7 N_XI12/XI6/NET36_XI12/XI6/MM7_d N_XI12/XI6/NET35_XI12/XI6/MM7_g
+ N_VSS_XI12/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM8 N_XI12/XI6/NET35_XI12/XI6/MM8_d N_WL<21>_XI12/XI6/MM8_g
+ N_BLN<9>_XI12/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI6/MM5 N_XI12/XI6/NET34_XI12/XI6/MM5_d N_XI12/XI6/NET33_XI12/XI6/MM5_g
+ N_VDD_XI12/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI6/MM4 N_XI12/XI6/NET33_XI12/XI6/MM4_d N_XI12/XI6/NET34_XI12/XI6/MM4_g
+ N_VDD_XI12/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI6/MM10 N_XI12/XI6/NET35_XI12/XI6/MM10_d N_XI12/XI6/NET36_XI12/XI6/MM10_g
+ N_VDD_XI12/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI6/MM11 N_XI12/XI6/NET36_XI12/XI6/MM11_d N_XI12/XI6/NET35_XI12/XI6/MM11_g
+ N_VDD_XI12/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI7/MM2 N_XI12/XI7/NET34_XI12/XI7/MM2_d N_XI12/XI7/NET33_XI12/XI7/MM2_g
+ N_VSS_XI12/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM3 N_XI12/XI7/NET33_XI12/XI7/MM3_d N_WL<20>_XI12/XI7/MM3_g
+ N_BLN<8>_XI12/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM0 N_XI12/XI7/NET34_XI12/XI7/MM0_d N_WL<20>_XI12/XI7/MM0_g
+ N_BL<8>_XI12/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM1 N_XI12/XI7/NET33_XI12/XI7/MM1_d N_XI12/XI7/NET34_XI12/XI7/MM1_g
+ N_VSS_XI12/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM9 N_XI12/XI7/NET36_XI12/XI7/MM9_d N_WL<21>_XI12/XI7/MM9_g
+ N_BL<8>_XI12/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM6 N_XI12/XI7/NET35_XI12/XI7/MM6_d N_XI12/XI7/NET36_XI12/XI7/MM6_g
+ N_VSS_XI12/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM7 N_XI12/XI7/NET36_XI12/XI7/MM7_d N_XI12/XI7/NET35_XI12/XI7/MM7_g
+ N_VSS_XI12/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM8 N_XI12/XI7/NET35_XI12/XI7/MM8_d N_WL<21>_XI12/XI7/MM8_g
+ N_BLN<8>_XI12/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI7/MM5 N_XI12/XI7/NET34_XI12/XI7/MM5_d N_XI12/XI7/NET33_XI12/XI7/MM5_g
+ N_VDD_XI12/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI7/MM4 N_XI12/XI7/NET33_XI12/XI7/MM4_d N_XI12/XI7/NET34_XI12/XI7/MM4_g
+ N_VDD_XI12/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI7/MM10 N_XI12/XI7/NET35_XI12/XI7/MM10_d N_XI12/XI7/NET36_XI12/XI7/MM10_g
+ N_VDD_XI12/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI7/MM11 N_XI12/XI7/NET36_XI12/XI7/MM11_d N_XI12/XI7/NET35_XI12/XI7/MM11_g
+ N_VDD_XI12/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI8/MM2 N_XI12/XI8/NET34_XI12/XI8/MM2_d N_XI12/XI8/NET33_XI12/XI8/MM2_g
+ N_VSS_XI12/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM3 N_XI12/XI8/NET33_XI12/XI8/MM3_d N_WL<20>_XI12/XI8/MM3_g
+ N_BLN<7>_XI12/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM0 N_XI12/XI8/NET34_XI12/XI8/MM0_d N_WL<20>_XI12/XI8/MM0_g
+ N_BL<7>_XI12/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM1 N_XI12/XI8/NET33_XI12/XI8/MM1_d N_XI12/XI8/NET34_XI12/XI8/MM1_g
+ N_VSS_XI12/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM9 N_XI12/XI8/NET36_XI12/XI8/MM9_d N_WL<21>_XI12/XI8/MM9_g
+ N_BL<7>_XI12/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM6 N_XI12/XI8/NET35_XI12/XI8/MM6_d N_XI12/XI8/NET36_XI12/XI8/MM6_g
+ N_VSS_XI12/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM7 N_XI12/XI8/NET36_XI12/XI8/MM7_d N_XI12/XI8/NET35_XI12/XI8/MM7_g
+ N_VSS_XI12/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM8 N_XI12/XI8/NET35_XI12/XI8/MM8_d N_WL<21>_XI12/XI8/MM8_g
+ N_BLN<7>_XI12/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI8/MM5 N_XI12/XI8/NET34_XI12/XI8/MM5_d N_XI12/XI8/NET33_XI12/XI8/MM5_g
+ N_VDD_XI12/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI8/MM4 N_XI12/XI8/NET33_XI12/XI8/MM4_d N_XI12/XI8/NET34_XI12/XI8/MM4_g
+ N_VDD_XI12/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI8/MM10 N_XI12/XI8/NET35_XI12/XI8/MM10_d N_XI12/XI8/NET36_XI12/XI8/MM10_g
+ N_VDD_XI12/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI8/MM11 N_XI12/XI8/NET36_XI12/XI8/MM11_d N_XI12/XI8/NET35_XI12/XI8/MM11_g
+ N_VDD_XI12/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI9/MM2 N_XI12/XI9/NET34_XI12/XI9/MM2_d N_XI12/XI9/NET33_XI12/XI9/MM2_g
+ N_VSS_XI12/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM3 N_XI12/XI9/NET33_XI12/XI9/MM3_d N_WL<20>_XI12/XI9/MM3_g
+ N_BLN<6>_XI12/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM0 N_XI12/XI9/NET34_XI12/XI9/MM0_d N_WL<20>_XI12/XI9/MM0_g
+ N_BL<6>_XI12/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM1 N_XI12/XI9/NET33_XI12/XI9/MM1_d N_XI12/XI9/NET34_XI12/XI9/MM1_g
+ N_VSS_XI12/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM9 N_XI12/XI9/NET36_XI12/XI9/MM9_d N_WL<21>_XI12/XI9/MM9_g
+ N_BL<6>_XI12/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM6 N_XI12/XI9/NET35_XI12/XI9/MM6_d N_XI12/XI9/NET36_XI12/XI9/MM6_g
+ N_VSS_XI12/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM7 N_XI12/XI9/NET36_XI12/XI9/MM7_d N_XI12/XI9/NET35_XI12/XI9/MM7_g
+ N_VSS_XI12/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM8 N_XI12/XI9/NET35_XI12/XI9/MM8_d N_WL<21>_XI12/XI9/MM8_g
+ N_BLN<6>_XI12/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI9/MM5 N_XI12/XI9/NET34_XI12/XI9/MM5_d N_XI12/XI9/NET33_XI12/XI9/MM5_g
+ N_VDD_XI12/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI9/MM4 N_XI12/XI9/NET33_XI12/XI9/MM4_d N_XI12/XI9/NET34_XI12/XI9/MM4_g
+ N_VDD_XI12/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI9/MM10 N_XI12/XI9/NET35_XI12/XI9/MM10_d N_XI12/XI9/NET36_XI12/XI9/MM10_g
+ N_VDD_XI12/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI9/MM11 N_XI12/XI9/NET36_XI12/XI9/MM11_d N_XI12/XI9/NET35_XI12/XI9/MM11_g
+ N_VDD_XI12/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI10/MM2 N_XI12/XI10/NET34_XI12/XI10/MM2_d
+ N_XI12/XI10/NET33_XI12/XI10/MM2_g N_VSS_XI12/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI10/MM3 N_XI12/XI10/NET33_XI12/XI10/MM3_d N_WL<20>_XI12/XI10/MM3_g
+ N_BLN<5>_XI12/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI10/MM0 N_XI12/XI10/NET34_XI12/XI10/MM0_d N_WL<20>_XI12/XI10/MM0_g
+ N_BL<5>_XI12/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI10/MM1 N_XI12/XI10/NET33_XI12/XI10/MM1_d
+ N_XI12/XI10/NET34_XI12/XI10/MM1_g N_VSS_XI12/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI10/MM9 N_XI12/XI10/NET36_XI12/XI10/MM9_d N_WL<21>_XI12/XI10/MM9_g
+ N_BL<5>_XI12/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI10/MM6 N_XI12/XI10/NET35_XI12/XI10/MM6_d
+ N_XI12/XI10/NET36_XI12/XI10/MM6_g N_VSS_XI12/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI10/MM7 N_XI12/XI10/NET36_XI12/XI10/MM7_d
+ N_XI12/XI10/NET35_XI12/XI10/MM7_g N_VSS_XI12/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI10/MM8 N_XI12/XI10/NET35_XI12/XI10/MM8_d N_WL<21>_XI12/XI10/MM8_g
+ N_BLN<5>_XI12/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI10/MM5 N_XI12/XI10/NET34_XI12/XI10/MM5_d
+ N_XI12/XI10/NET33_XI12/XI10/MM5_g N_VDD_XI12/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI10/MM4 N_XI12/XI10/NET33_XI12/XI10/MM4_d
+ N_XI12/XI10/NET34_XI12/XI10/MM4_g N_VDD_XI12/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI10/MM10 N_XI12/XI10/NET35_XI12/XI10/MM10_d
+ N_XI12/XI10/NET36_XI12/XI10/MM10_g N_VDD_XI12/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI10/MM11 N_XI12/XI10/NET36_XI12/XI10/MM11_d
+ N_XI12/XI10/NET35_XI12/XI10/MM11_g N_VDD_XI12/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI11/MM2 N_XI12/XI11/NET34_XI12/XI11/MM2_d
+ N_XI12/XI11/NET33_XI12/XI11/MM2_g N_VSS_XI12/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI11/MM3 N_XI12/XI11/NET33_XI12/XI11/MM3_d N_WL<20>_XI12/XI11/MM3_g
+ N_BLN<4>_XI12/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI11/MM0 N_XI12/XI11/NET34_XI12/XI11/MM0_d N_WL<20>_XI12/XI11/MM0_g
+ N_BL<4>_XI12/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI11/MM1 N_XI12/XI11/NET33_XI12/XI11/MM1_d
+ N_XI12/XI11/NET34_XI12/XI11/MM1_g N_VSS_XI12/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI11/MM9 N_XI12/XI11/NET36_XI12/XI11/MM9_d N_WL<21>_XI12/XI11/MM9_g
+ N_BL<4>_XI12/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI11/MM6 N_XI12/XI11/NET35_XI12/XI11/MM6_d
+ N_XI12/XI11/NET36_XI12/XI11/MM6_g N_VSS_XI12/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI11/MM7 N_XI12/XI11/NET36_XI12/XI11/MM7_d
+ N_XI12/XI11/NET35_XI12/XI11/MM7_g N_VSS_XI12/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI11/MM8 N_XI12/XI11/NET35_XI12/XI11/MM8_d N_WL<21>_XI12/XI11/MM8_g
+ N_BLN<4>_XI12/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI11/MM5 N_XI12/XI11/NET34_XI12/XI11/MM5_d
+ N_XI12/XI11/NET33_XI12/XI11/MM5_g N_VDD_XI12/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI11/MM4 N_XI12/XI11/NET33_XI12/XI11/MM4_d
+ N_XI12/XI11/NET34_XI12/XI11/MM4_g N_VDD_XI12/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI11/MM10 N_XI12/XI11/NET35_XI12/XI11/MM10_d
+ N_XI12/XI11/NET36_XI12/XI11/MM10_g N_VDD_XI12/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI11/MM11 N_XI12/XI11/NET36_XI12/XI11/MM11_d
+ N_XI12/XI11/NET35_XI12/XI11/MM11_g N_VDD_XI12/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI12/MM2 N_XI12/XI12/NET34_XI12/XI12/MM2_d
+ N_XI12/XI12/NET33_XI12/XI12/MM2_g N_VSS_XI12/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI12/MM3 N_XI12/XI12/NET33_XI12/XI12/MM3_d N_WL<20>_XI12/XI12/MM3_g
+ N_BLN<3>_XI12/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI12/MM0 N_XI12/XI12/NET34_XI12/XI12/MM0_d N_WL<20>_XI12/XI12/MM0_g
+ N_BL<3>_XI12/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI12/MM1 N_XI12/XI12/NET33_XI12/XI12/MM1_d
+ N_XI12/XI12/NET34_XI12/XI12/MM1_g N_VSS_XI12/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI12/MM9 N_XI12/XI12/NET36_XI12/XI12/MM9_d N_WL<21>_XI12/XI12/MM9_g
+ N_BL<3>_XI12/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI12/MM6 N_XI12/XI12/NET35_XI12/XI12/MM6_d
+ N_XI12/XI12/NET36_XI12/XI12/MM6_g N_VSS_XI12/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI12/MM7 N_XI12/XI12/NET36_XI12/XI12/MM7_d
+ N_XI12/XI12/NET35_XI12/XI12/MM7_g N_VSS_XI12/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI12/MM8 N_XI12/XI12/NET35_XI12/XI12/MM8_d N_WL<21>_XI12/XI12/MM8_g
+ N_BLN<3>_XI12/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI12/MM5 N_XI12/XI12/NET34_XI12/XI12/MM5_d
+ N_XI12/XI12/NET33_XI12/XI12/MM5_g N_VDD_XI12/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI12/MM4 N_XI12/XI12/NET33_XI12/XI12/MM4_d
+ N_XI12/XI12/NET34_XI12/XI12/MM4_g N_VDD_XI12/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI12/MM10 N_XI12/XI12/NET35_XI12/XI12/MM10_d
+ N_XI12/XI12/NET36_XI12/XI12/MM10_g N_VDD_XI12/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI12/MM11 N_XI12/XI12/NET36_XI12/XI12/MM11_d
+ N_XI12/XI12/NET35_XI12/XI12/MM11_g N_VDD_XI12/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI13/MM2 N_XI12/XI13/NET34_XI12/XI13/MM2_d
+ N_XI12/XI13/NET33_XI12/XI13/MM2_g N_VSS_XI12/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI13/MM3 N_XI12/XI13/NET33_XI12/XI13/MM3_d N_WL<20>_XI12/XI13/MM3_g
+ N_BLN<2>_XI12/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI13/MM0 N_XI12/XI13/NET34_XI12/XI13/MM0_d N_WL<20>_XI12/XI13/MM0_g
+ N_BL<2>_XI12/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI13/MM1 N_XI12/XI13/NET33_XI12/XI13/MM1_d
+ N_XI12/XI13/NET34_XI12/XI13/MM1_g N_VSS_XI12/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI13/MM9 N_XI12/XI13/NET36_XI12/XI13/MM9_d N_WL<21>_XI12/XI13/MM9_g
+ N_BL<2>_XI12/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI13/MM6 N_XI12/XI13/NET35_XI12/XI13/MM6_d
+ N_XI12/XI13/NET36_XI12/XI13/MM6_g N_VSS_XI12/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI13/MM7 N_XI12/XI13/NET36_XI12/XI13/MM7_d
+ N_XI12/XI13/NET35_XI12/XI13/MM7_g N_VSS_XI12/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI13/MM8 N_XI12/XI13/NET35_XI12/XI13/MM8_d N_WL<21>_XI12/XI13/MM8_g
+ N_BLN<2>_XI12/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI13/MM5 N_XI12/XI13/NET34_XI12/XI13/MM5_d
+ N_XI12/XI13/NET33_XI12/XI13/MM5_g N_VDD_XI12/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI13/MM4 N_XI12/XI13/NET33_XI12/XI13/MM4_d
+ N_XI12/XI13/NET34_XI12/XI13/MM4_g N_VDD_XI12/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI13/MM10 N_XI12/XI13/NET35_XI12/XI13/MM10_d
+ N_XI12/XI13/NET36_XI12/XI13/MM10_g N_VDD_XI12/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI13/MM11 N_XI12/XI13/NET36_XI12/XI13/MM11_d
+ N_XI12/XI13/NET35_XI12/XI13/MM11_g N_VDD_XI12/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI14/MM2 N_XI12/XI14/NET34_XI12/XI14/MM2_d
+ N_XI12/XI14/NET33_XI12/XI14/MM2_g N_VSS_XI12/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI14/MM3 N_XI12/XI14/NET33_XI12/XI14/MM3_d N_WL<20>_XI12/XI14/MM3_g
+ N_BLN<1>_XI12/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI14/MM0 N_XI12/XI14/NET34_XI12/XI14/MM0_d N_WL<20>_XI12/XI14/MM0_g
+ N_BL<1>_XI12/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI14/MM1 N_XI12/XI14/NET33_XI12/XI14/MM1_d
+ N_XI12/XI14/NET34_XI12/XI14/MM1_g N_VSS_XI12/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI14/MM9 N_XI12/XI14/NET36_XI12/XI14/MM9_d N_WL<21>_XI12/XI14/MM9_g
+ N_BL<1>_XI12/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI14/MM6 N_XI12/XI14/NET35_XI12/XI14/MM6_d
+ N_XI12/XI14/NET36_XI12/XI14/MM6_g N_VSS_XI12/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI14/MM7 N_XI12/XI14/NET36_XI12/XI14/MM7_d
+ N_XI12/XI14/NET35_XI12/XI14/MM7_g N_VSS_XI12/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI14/MM8 N_XI12/XI14/NET35_XI12/XI14/MM8_d N_WL<21>_XI12/XI14/MM8_g
+ N_BLN<1>_XI12/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI14/MM5 N_XI12/XI14/NET34_XI12/XI14/MM5_d
+ N_XI12/XI14/NET33_XI12/XI14/MM5_g N_VDD_XI12/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI14/MM4 N_XI12/XI14/NET33_XI12/XI14/MM4_d
+ N_XI12/XI14/NET34_XI12/XI14/MM4_g N_VDD_XI12/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI14/MM10 N_XI12/XI14/NET35_XI12/XI14/MM10_d
+ N_XI12/XI14/NET36_XI12/XI14/MM10_g N_VDD_XI12/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI14/MM11 N_XI12/XI14/NET36_XI12/XI14/MM11_d
+ N_XI12/XI14/NET35_XI12/XI14/MM11_g N_VDD_XI12/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI15/MM2 N_XI12/XI15/NET34_XI12/XI15/MM2_d
+ N_XI12/XI15/NET33_XI12/XI15/MM2_g N_VSS_XI12/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI15/MM3 N_XI12/XI15/NET33_XI12/XI15/MM3_d N_WL<20>_XI12/XI15/MM3_g
+ N_BLN<0>_XI12/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI15/MM0 N_XI12/XI15/NET34_XI12/XI15/MM0_d N_WL<20>_XI12/XI15/MM0_g
+ N_BL<0>_XI12/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI15/MM1 N_XI12/XI15/NET33_XI12/XI15/MM1_d
+ N_XI12/XI15/NET34_XI12/XI15/MM1_g N_VSS_XI12/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI15/MM9 N_XI12/XI15/NET36_XI12/XI15/MM9_d N_WL<21>_XI12/XI15/MM9_g
+ N_BL<0>_XI12/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI15/MM6 N_XI12/XI15/NET35_XI12/XI15/MM6_d
+ N_XI12/XI15/NET36_XI12/XI15/MM6_g N_VSS_XI12/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI15/MM7 N_XI12/XI15/NET36_XI12/XI15/MM7_d
+ N_XI12/XI15/NET35_XI12/XI15/MM7_g N_VSS_XI12/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/XI15/MM8 N_XI12/XI15/NET35_XI12/XI15/MM8_d N_WL<21>_XI12/XI15/MM8_g
+ N_BLN<0>_XI12/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI12/XI15/MM5 N_XI12/XI15/NET34_XI12/XI15/MM5_d
+ N_XI12/XI15/NET33_XI12/XI15/MM5_g N_VDD_XI12/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI15/MM4 N_XI12/XI15/NET33_XI12/XI15/MM4_d
+ N_XI12/XI15/NET34_XI12/XI15/MM4_g N_VDD_XI12/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI15/MM10 N_XI12/XI15/NET35_XI12/XI15/MM10_d
+ N_XI12/XI15/NET36_XI12/XI15/MM10_g N_VDD_XI12/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/XI15/MM11 N_XI12/XI15/NET36_XI12/XI15/MM11_d
+ N_XI12/XI15/NET35_XI12/XI15/MM11_g N_VDD_XI12/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI0/MM2 N_XI13/XI0/NET34_XI13/XI0/MM2_d N_XI13/XI0/NET33_XI13/XI0/MM2_g
+ N_VSS_XI13/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI0/MM3 N_XI13/XI0/NET33_XI13/XI0/MM3_d N_WL<22>_XI13/XI0/MM3_g
+ N_BLN<15>_XI13/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI0/MM0 N_XI13/XI0/NET34_XI13/XI0/MM0_d N_WL<22>_XI13/XI0/MM0_g
+ N_BL<15>_XI13/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI0/MM1 N_XI13/XI0/NET33_XI13/XI0/MM1_d N_XI13/XI0/NET34_XI13/XI0/MM1_g
+ N_VSS_XI13/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI0/MM9 N_XI13/XI0/NET36_XI13/XI0/MM9_d N_WL<23>_XI13/XI0/MM9_g
+ N_BL<15>_XI13/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI0/MM6 N_XI13/XI0/NET35_XI13/XI0/MM6_d N_XI13/XI0/NET36_XI13/XI0/MM6_g
+ N_VSS_XI13/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI0/MM7 N_XI13/XI0/NET36_XI13/XI0/MM7_d N_XI13/XI0/NET35_XI13/XI0/MM7_g
+ N_VSS_XI13/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI0/MM8 N_XI13/XI0/NET35_XI13/XI0/MM8_d N_WL<23>_XI13/XI0/MM8_g
+ N_BLN<15>_XI13/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI0/MM5 N_XI13/XI0/NET34_XI13/XI0/MM5_d N_XI13/XI0/NET33_XI13/XI0/MM5_g
+ N_VDD_XI13/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI0/MM4 N_XI13/XI0/NET33_XI13/XI0/MM4_d N_XI13/XI0/NET34_XI13/XI0/MM4_g
+ N_VDD_XI13/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI0/MM10 N_XI13/XI0/NET35_XI13/XI0/MM10_d N_XI13/XI0/NET36_XI13/XI0/MM10_g
+ N_VDD_XI13/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI0/MM11 N_XI13/XI0/NET36_XI13/XI0/MM11_d N_XI13/XI0/NET35_XI13/XI0/MM11_g
+ N_VDD_XI13/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI1/MM2 N_XI13/XI1/NET34_XI13/XI1/MM2_d N_XI13/XI1/NET33_XI13/XI1/MM2_g
+ N_VSS_XI13/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI1/MM3 N_XI13/XI1/NET33_XI13/XI1/MM3_d N_WL<22>_XI13/XI1/MM3_g
+ N_BLN<14>_XI13/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI1/MM0 N_XI13/XI1/NET34_XI13/XI1/MM0_d N_WL<22>_XI13/XI1/MM0_g
+ N_BL<14>_XI13/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI1/MM1 N_XI13/XI1/NET33_XI13/XI1/MM1_d N_XI13/XI1/NET34_XI13/XI1/MM1_g
+ N_VSS_XI13/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI1/MM9 N_XI13/XI1/NET36_XI13/XI1/MM9_d N_WL<23>_XI13/XI1/MM9_g
+ N_BL<14>_XI13/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI1/MM6 N_XI13/XI1/NET35_XI13/XI1/MM6_d N_XI13/XI1/NET36_XI13/XI1/MM6_g
+ N_VSS_XI13/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI1/MM7 N_XI13/XI1/NET36_XI13/XI1/MM7_d N_XI13/XI1/NET35_XI13/XI1/MM7_g
+ N_VSS_XI13/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI1/MM8 N_XI13/XI1/NET35_XI13/XI1/MM8_d N_WL<23>_XI13/XI1/MM8_g
+ N_BLN<14>_XI13/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI1/MM5 N_XI13/XI1/NET34_XI13/XI1/MM5_d N_XI13/XI1/NET33_XI13/XI1/MM5_g
+ N_VDD_XI13/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI1/MM4 N_XI13/XI1/NET33_XI13/XI1/MM4_d N_XI13/XI1/NET34_XI13/XI1/MM4_g
+ N_VDD_XI13/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI1/MM10 N_XI13/XI1/NET35_XI13/XI1/MM10_d N_XI13/XI1/NET36_XI13/XI1/MM10_g
+ N_VDD_XI13/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI1/MM11 N_XI13/XI1/NET36_XI13/XI1/MM11_d N_XI13/XI1/NET35_XI13/XI1/MM11_g
+ N_VDD_XI13/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI2/MM2 N_XI13/XI2/NET34_XI13/XI2/MM2_d N_XI13/XI2/NET33_XI13/XI2/MM2_g
+ N_VSS_XI13/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI2/MM3 N_XI13/XI2/NET33_XI13/XI2/MM3_d N_WL<22>_XI13/XI2/MM3_g
+ N_BLN<13>_XI13/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI2/MM0 N_XI13/XI2/NET34_XI13/XI2/MM0_d N_WL<22>_XI13/XI2/MM0_g
+ N_BL<13>_XI13/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI2/MM1 N_XI13/XI2/NET33_XI13/XI2/MM1_d N_XI13/XI2/NET34_XI13/XI2/MM1_g
+ N_VSS_XI13/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI2/MM9 N_XI13/XI2/NET36_XI13/XI2/MM9_d N_WL<23>_XI13/XI2/MM9_g
+ N_BL<13>_XI13/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI2/MM6 N_XI13/XI2/NET35_XI13/XI2/MM6_d N_XI13/XI2/NET36_XI13/XI2/MM6_g
+ N_VSS_XI13/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI2/MM7 N_XI13/XI2/NET36_XI13/XI2/MM7_d N_XI13/XI2/NET35_XI13/XI2/MM7_g
+ N_VSS_XI13/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI2/MM8 N_XI13/XI2/NET35_XI13/XI2/MM8_d N_WL<23>_XI13/XI2/MM8_g
+ N_BLN<13>_XI13/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI2/MM5 N_XI13/XI2/NET34_XI13/XI2/MM5_d N_XI13/XI2/NET33_XI13/XI2/MM5_g
+ N_VDD_XI13/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI2/MM4 N_XI13/XI2/NET33_XI13/XI2/MM4_d N_XI13/XI2/NET34_XI13/XI2/MM4_g
+ N_VDD_XI13/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI2/MM10 N_XI13/XI2/NET35_XI13/XI2/MM10_d N_XI13/XI2/NET36_XI13/XI2/MM10_g
+ N_VDD_XI13/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI2/MM11 N_XI13/XI2/NET36_XI13/XI2/MM11_d N_XI13/XI2/NET35_XI13/XI2/MM11_g
+ N_VDD_XI13/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI3/MM2 N_XI13/XI3/NET34_XI13/XI3/MM2_d N_XI13/XI3/NET33_XI13/XI3/MM2_g
+ N_VSS_XI13/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI3/MM3 N_XI13/XI3/NET33_XI13/XI3/MM3_d N_WL<22>_XI13/XI3/MM3_g
+ N_BLN<12>_XI13/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI3/MM0 N_XI13/XI3/NET34_XI13/XI3/MM0_d N_WL<22>_XI13/XI3/MM0_g
+ N_BL<12>_XI13/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI3/MM1 N_XI13/XI3/NET33_XI13/XI3/MM1_d N_XI13/XI3/NET34_XI13/XI3/MM1_g
+ N_VSS_XI13/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI3/MM9 N_XI13/XI3/NET36_XI13/XI3/MM9_d N_WL<23>_XI13/XI3/MM9_g
+ N_BL<12>_XI13/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI3/MM6 N_XI13/XI3/NET35_XI13/XI3/MM6_d N_XI13/XI3/NET36_XI13/XI3/MM6_g
+ N_VSS_XI13/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI3/MM7 N_XI13/XI3/NET36_XI13/XI3/MM7_d N_XI13/XI3/NET35_XI13/XI3/MM7_g
+ N_VSS_XI13/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI3/MM8 N_XI13/XI3/NET35_XI13/XI3/MM8_d N_WL<23>_XI13/XI3/MM8_g
+ N_BLN<12>_XI13/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI3/MM5 N_XI13/XI3/NET34_XI13/XI3/MM5_d N_XI13/XI3/NET33_XI13/XI3/MM5_g
+ N_VDD_XI13/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI3/MM4 N_XI13/XI3/NET33_XI13/XI3/MM4_d N_XI13/XI3/NET34_XI13/XI3/MM4_g
+ N_VDD_XI13/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI3/MM10 N_XI13/XI3/NET35_XI13/XI3/MM10_d N_XI13/XI3/NET36_XI13/XI3/MM10_g
+ N_VDD_XI13/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI3/MM11 N_XI13/XI3/NET36_XI13/XI3/MM11_d N_XI13/XI3/NET35_XI13/XI3/MM11_g
+ N_VDD_XI13/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI4/MM2 N_XI13/XI4/NET34_XI13/XI4/MM2_d N_XI13/XI4/NET33_XI13/XI4/MM2_g
+ N_VSS_XI13/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI4/MM3 N_XI13/XI4/NET33_XI13/XI4/MM3_d N_WL<22>_XI13/XI4/MM3_g
+ N_BLN<11>_XI13/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI4/MM0 N_XI13/XI4/NET34_XI13/XI4/MM0_d N_WL<22>_XI13/XI4/MM0_g
+ N_BL<11>_XI13/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI4/MM1 N_XI13/XI4/NET33_XI13/XI4/MM1_d N_XI13/XI4/NET34_XI13/XI4/MM1_g
+ N_VSS_XI13/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI4/MM9 N_XI13/XI4/NET36_XI13/XI4/MM9_d N_WL<23>_XI13/XI4/MM9_g
+ N_BL<11>_XI13/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI4/MM6 N_XI13/XI4/NET35_XI13/XI4/MM6_d N_XI13/XI4/NET36_XI13/XI4/MM6_g
+ N_VSS_XI13/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI4/MM7 N_XI13/XI4/NET36_XI13/XI4/MM7_d N_XI13/XI4/NET35_XI13/XI4/MM7_g
+ N_VSS_XI13/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI4/MM8 N_XI13/XI4/NET35_XI13/XI4/MM8_d N_WL<23>_XI13/XI4/MM8_g
+ N_BLN<11>_XI13/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI4/MM5 N_XI13/XI4/NET34_XI13/XI4/MM5_d N_XI13/XI4/NET33_XI13/XI4/MM5_g
+ N_VDD_XI13/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI4/MM4 N_XI13/XI4/NET33_XI13/XI4/MM4_d N_XI13/XI4/NET34_XI13/XI4/MM4_g
+ N_VDD_XI13/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI4/MM10 N_XI13/XI4/NET35_XI13/XI4/MM10_d N_XI13/XI4/NET36_XI13/XI4/MM10_g
+ N_VDD_XI13/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI4/MM11 N_XI13/XI4/NET36_XI13/XI4/MM11_d N_XI13/XI4/NET35_XI13/XI4/MM11_g
+ N_VDD_XI13/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI5/MM2 N_XI13/XI5/NET34_XI13/XI5/MM2_d N_XI13/XI5/NET33_XI13/XI5/MM2_g
+ N_VSS_XI13/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI5/MM3 N_XI13/XI5/NET33_XI13/XI5/MM3_d N_WL<22>_XI13/XI5/MM3_g
+ N_BLN<10>_XI13/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI5/MM0 N_XI13/XI5/NET34_XI13/XI5/MM0_d N_WL<22>_XI13/XI5/MM0_g
+ N_BL<10>_XI13/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI5/MM1 N_XI13/XI5/NET33_XI13/XI5/MM1_d N_XI13/XI5/NET34_XI13/XI5/MM1_g
+ N_VSS_XI13/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI5/MM9 N_XI13/XI5/NET36_XI13/XI5/MM9_d N_WL<23>_XI13/XI5/MM9_g
+ N_BL<10>_XI13/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI5/MM6 N_XI13/XI5/NET35_XI13/XI5/MM6_d N_XI13/XI5/NET36_XI13/XI5/MM6_g
+ N_VSS_XI13/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI5/MM7 N_XI13/XI5/NET36_XI13/XI5/MM7_d N_XI13/XI5/NET35_XI13/XI5/MM7_g
+ N_VSS_XI13/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI5/MM8 N_XI13/XI5/NET35_XI13/XI5/MM8_d N_WL<23>_XI13/XI5/MM8_g
+ N_BLN<10>_XI13/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI5/MM5 N_XI13/XI5/NET34_XI13/XI5/MM5_d N_XI13/XI5/NET33_XI13/XI5/MM5_g
+ N_VDD_XI13/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI5/MM4 N_XI13/XI5/NET33_XI13/XI5/MM4_d N_XI13/XI5/NET34_XI13/XI5/MM4_g
+ N_VDD_XI13/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI5/MM10 N_XI13/XI5/NET35_XI13/XI5/MM10_d N_XI13/XI5/NET36_XI13/XI5/MM10_g
+ N_VDD_XI13/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI5/MM11 N_XI13/XI5/NET36_XI13/XI5/MM11_d N_XI13/XI5/NET35_XI13/XI5/MM11_g
+ N_VDD_XI13/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI6/MM2 N_XI13/XI6/NET34_XI13/XI6/MM2_d N_XI13/XI6/NET33_XI13/XI6/MM2_g
+ N_VSS_XI13/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM3 N_XI13/XI6/NET33_XI13/XI6/MM3_d N_WL<22>_XI13/XI6/MM3_g
+ N_BLN<9>_XI13/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM0 N_XI13/XI6/NET34_XI13/XI6/MM0_d N_WL<22>_XI13/XI6/MM0_g
+ N_BL<9>_XI13/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM1 N_XI13/XI6/NET33_XI13/XI6/MM1_d N_XI13/XI6/NET34_XI13/XI6/MM1_g
+ N_VSS_XI13/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM9 N_XI13/XI6/NET36_XI13/XI6/MM9_d N_WL<23>_XI13/XI6/MM9_g
+ N_BL<9>_XI13/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM6 N_XI13/XI6/NET35_XI13/XI6/MM6_d N_XI13/XI6/NET36_XI13/XI6/MM6_g
+ N_VSS_XI13/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM7 N_XI13/XI6/NET36_XI13/XI6/MM7_d N_XI13/XI6/NET35_XI13/XI6/MM7_g
+ N_VSS_XI13/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM8 N_XI13/XI6/NET35_XI13/XI6/MM8_d N_WL<23>_XI13/XI6/MM8_g
+ N_BLN<9>_XI13/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI6/MM5 N_XI13/XI6/NET34_XI13/XI6/MM5_d N_XI13/XI6/NET33_XI13/XI6/MM5_g
+ N_VDD_XI13/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI6/MM4 N_XI13/XI6/NET33_XI13/XI6/MM4_d N_XI13/XI6/NET34_XI13/XI6/MM4_g
+ N_VDD_XI13/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI6/MM10 N_XI13/XI6/NET35_XI13/XI6/MM10_d N_XI13/XI6/NET36_XI13/XI6/MM10_g
+ N_VDD_XI13/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI6/MM11 N_XI13/XI6/NET36_XI13/XI6/MM11_d N_XI13/XI6/NET35_XI13/XI6/MM11_g
+ N_VDD_XI13/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI7/MM2 N_XI13/XI7/NET34_XI13/XI7/MM2_d N_XI13/XI7/NET33_XI13/XI7/MM2_g
+ N_VSS_XI13/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM3 N_XI13/XI7/NET33_XI13/XI7/MM3_d N_WL<22>_XI13/XI7/MM3_g
+ N_BLN<8>_XI13/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM0 N_XI13/XI7/NET34_XI13/XI7/MM0_d N_WL<22>_XI13/XI7/MM0_g
+ N_BL<8>_XI13/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM1 N_XI13/XI7/NET33_XI13/XI7/MM1_d N_XI13/XI7/NET34_XI13/XI7/MM1_g
+ N_VSS_XI13/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM9 N_XI13/XI7/NET36_XI13/XI7/MM9_d N_WL<23>_XI13/XI7/MM9_g
+ N_BL<8>_XI13/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM6 N_XI13/XI7/NET35_XI13/XI7/MM6_d N_XI13/XI7/NET36_XI13/XI7/MM6_g
+ N_VSS_XI13/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM7 N_XI13/XI7/NET36_XI13/XI7/MM7_d N_XI13/XI7/NET35_XI13/XI7/MM7_g
+ N_VSS_XI13/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM8 N_XI13/XI7/NET35_XI13/XI7/MM8_d N_WL<23>_XI13/XI7/MM8_g
+ N_BLN<8>_XI13/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI7/MM5 N_XI13/XI7/NET34_XI13/XI7/MM5_d N_XI13/XI7/NET33_XI13/XI7/MM5_g
+ N_VDD_XI13/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI7/MM4 N_XI13/XI7/NET33_XI13/XI7/MM4_d N_XI13/XI7/NET34_XI13/XI7/MM4_g
+ N_VDD_XI13/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI7/MM10 N_XI13/XI7/NET35_XI13/XI7/MM10_d N_XI13/XI7/NET36_XI13/XI7/MM10_g
+ N_VDD_XI13/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI7/MM11 N_XI13/XI7/NET36_XI13/XI7/MM11_d N_XI13/XI7/NET35_XI13/XI7/MM11_g
+ N_VDD_XI13/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI8/MM2 N_XI13/XI8/NET34_XI13/XI8/MM2_d N_XI13/XI8/NET33_XI13/XI8/MM2_g
+ N_VSS_XI13/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM3 N_XI13/XI8/NET33_XI13/XI8/MM3_d N_WL<22>_XI13/XI8/MM3_g
+ N_BLN<7>_XI13/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM0 N_XI13/XI8/NET34_XI13/XI8/MM0_d N_WL<22>_XI13/XI8/MM0_g
+ N_BL<7>_XI13/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM1 N_XI13/XI8/NET33_XI13/XI8/MM1_d N_XI13/XI8/NET34_XI13/XI8/MM1_g
+ N_VSS_XI13/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM9 N_XI13/XI8/NET36_XI13/XI8/MM9_d N_WL<23>_XI13/XI8/MM9_g
+ N_BL<7>_XI13/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM6 N_XI13/XI8/NET35_XI13/XI8/MM6_d N_XI13/XI8/NET36_XI13/XI8/MM6_g
+ N_VSS_XI13/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM7 N_XI13/XI8/NET36_XI13/XI8/MM7_d N_XI13/XI8/NET35_XI13/XI8/MM7_g
+ N_VSS_XI13/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM8 N_XI13/XI8/NET35_XI13/XI8/MM8_d N_WL<23>_XI13/XI8/MM8_g
+ N_BLN<7>_XI13/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI8/MM5 N_XI13/XI8/NET34_XI13/XI8/MM5_d N_XI13/XI8/NET33_XI13/XI8/MM5_g
+ N_VDD_XI13/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI8/MM4 N_XI13/XI8/NET33_XI13/XI8/MM4_d N_XI13/XI8/NET34_XI13/XI8/MM4_g
+ N_VDD_XI13/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI8/MM10 N_XI13/XI8/NET35_XI13/XI8/MM10_d N_XI13/XI8/NET36_XI13/XI8/MM10_g
+ N_VDD_XI13/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI8/MM11 N_XI13/XI8/NET36_XI13/XI8/MM11_d N_XI13/XI8/NET35_XI13/XI8/MM11_g
+ N_VDD_XI13/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI9/MM2 N_XI13/XI9/NET34_XI13/XI9/MM2_d N_XI13/XI9/NET33_XI13/XI9/MM2_g
+ N_VSS_XI13/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM3 N_XI13/XI9/NET33_XI13/XI9/MM3_d N_WL<22>_XI13/XI9/MM3_g
+ N_BLN<6>_XI13/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM0 N_XI13/XI9/NET34_XI13/XI9/MM0_d N_WL<22>_XI13/XI9/MM0_g
+ N_BL<6>_XI13/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM1 N_XI13/XI9/NET33_XI13/XI9/MM1_d N_XI13/XI9/NET34_XI13/XI9/MM1_g
+ N_VSS_XI13/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM9 N_XI13/XI9/NET36_XI13/XI9/MM9_d N_WL<23>_XI13/XI9/MM9_g
+ N_BL<6>_XI13/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM6 N_XI13/XI9/NET35_XI13/XI9/MM6_d N_XI13/XI9/NET36_XI13/XI9/MM6_g
+ N_VSS_XI13/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM7 N_XI13/XI9/NET36_XI13/XI9/MM7_d N_XI13/XI9/NET35_XI13/XI9/MM7_g
+ N_VSS_XI13/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM8 N_XI13/XI9/NET35_XI13/XI9/MM8_d N_WL<23>_XI13/XI9/MM8_g
+ N_BLN<6>_XI13/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI9/MM5 N_XI13/XI9/NET34_XI13/XI9/MM5_d N_XI13/XI9/NET33_XI13/XI9/MM5_g
+ N_VDD_XI13/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI9/MM4 N_XI13/XI9/NET33_XI13/XI9/MM4_d N_XI13/XI9/NET34_XI13/XI9/MM4_g
+ N_VDD_XI13/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI9/MM10 N_XI13/XI9/NET35_XI13/XI9/MM10_d N_XI13/XI9/NET36_XI13/XI9/MM10_g
+ N_VDD_XI13/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI9/MM11 N_XI13/XI9/NET36_XI13/XI9/MM11_d N_XI13/XI9/NET35_XI13/XI9/MM11_g
+ N_VDD_XI13/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI10/MM2 N_XI13/XI10/NET34_XI13/XI10/MM2_d
+ N_XI13/XI10/NET33_XI13/XI10/MM2_g N_VSS_XI13/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI10/MM3 N_XI13/XI10/NET33_XI13/XI10/MM3_d N_WL<22>_XI13/XI10/MM3_g
+ N_BLN<5>_XI13/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI10/MM0 N_XI13/XI10/NET34_XI13/XI10/MM0_d N_WL<22>_XI13/XI10/MM0_g
+ N_BL<5>_XI13/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI10/MM1 N_XI13/XI10/NET33_XI13/XI10/MM1_d
+ N_XI13/XI10/NET34_XI13/XI10/MM1_g N_VSS_XI13/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI10/MM9 N_XI13/XI10/NET36_XI13/XI10/MM9_d N_WL<23>_XI13/XI10/MM9_g
+ N_BL<5>_XI13/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI10/MM6 N_XI13/XI10/NET35_XI13/XI10/MM6_d
+ N_XI13/XI10/NET36_XI13/XI10/MM6_g N_VSS_XI13/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI10/MM7 N_XI13/XI10/NET36_XI13/XI10/MM7_d
+ N_XI13/XI10/NET35_XI13/XI10/MM7_g N_VSS_XI13/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI10/MM8 N_XI13/XI10/NET35_XI13/XI10/MM8_d N_WL<23>_XI13/XI10/MM8_g
+ N_BLN<5>_XI13/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI10/MM5 N_XI13/XI10/NET34_XI13/XI10/MM5_d
+ N_XI13/XI10/NET33_XI13/XI10/MM5_g N_VDD_XI13/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI10/MM4 N_XI13/XI10/NET33_XI13/XI10/MM4_d
+ N_XI13/XI10/NET34_XI13/XI10/MM4_g N_VDD_XI13/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI10/MM10 N_XI13/XI10/NET35_XI13/XI10/MM10_d
+ N_XI13/XI10/NET36_XI13/XI10/MM10_g N_VDD_XI13/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI10/MM11 N_XI13/XI10/NET36_XI13/XI10/MM11_d
+ N_XI13/XI10/NET35_XI13/XI10/MM11_g N_VDD_XI13/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI11/MM2 N_XI13/XI11/NET34_XI13/XI11/MM2_d
+ N_XI13/XI11/NET33_XI13/XI11/MM2_g N_VSS_XI13/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI11/MM3 N_XI13/XI11/NET33_XI13/XI11/MM3_d N_WL<22>_XI13/XI11/MM3_g
+ N_BLN<4>_XI13/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI11/MM0 N_XI13/XI11/NET34_XI13/XI11/MM0_d N_WL<22>_XI13/XI11/MM0_g
+ N_BL<4>_XI13/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI11/MM1 N_XI13/XI11/NET33_XI13/XI11/MM1_d
+ N_XI13/XI11/NET34_XI13/XI11/MM1_g N_VSS_XI13/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI11/MM9 N_XI13/XI11/NET36_XI13/XI11/MM9_d N_WL<23>_XI13/XI11/MM9_g
+ N_BL<4>_XI13/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI11/MM6 N_XI13/XI11/NET35_XI13/XI11/MM6_d
+ N_XI13/XI11/NET36_XI13/XI11/MM6_g N_VSS_XI13/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI11/MM7 N_XI13/XI11/NET36_XI13/XI11/MM7_d
+ N_XI13/XI11/NET35_XI13/XI11/MM7_g N_VSS_XI13/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI11/MM8 N_XI13/XI11/NET35_XI13/XI11/MM8_d N_WL<23>_XI13/XI11/MM8_g
+ N_BLN<4>_XI13/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI11/MM5 N_XI13/XI11/NET34_XI13/XI11/MM5_d
+ N_XI13/XI11/NET33_XI13/XI11/MM5_g N_VDD_XI13/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI11/MM4 N_XI13/XI11/NET33_XI13/XI11/MM4_d
+ N_XI13/XI11/NET34_XI13/XI11/MM4_g N_VDD_XI13/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI11/MM10 N_XI13/XI11/NET35_XI13/XI11/MM10_d
+ N_XI13/XI11/NET36_XI13/XI11/MM10_g N_VDD_XI13/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI11/MM11 N_XI13/XI11/NET36_XI13/XI11/MM11_d
+ N_XI13/XI11/NET35_XI13/XI11/MM11_g N_VDD_XI13/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI12/MM2 N_XI13/XI12/NET34_XI13/XI12/MM2_d
+ N_XI13/XI12/NET33_XI13/XI12/MM2_g N_VSS_XI13/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI12/MM3 N_XI13/XI12/NET33_XI13/XI12/MM3_d N_WL<22>_XI13/XI12/MM3_g
+ N_BLN<3>_XI13/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI12/MM0 N_XI13/XI12/NET34_XI13/XI12/MM0_d N_WL<22>_XI13/XI12/MM0_g
+ N_BL<3>_XI13/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI12/MM1 N_XI13/XI12/NET33_XI13/XI12/MM1_d
+ N_XI13/XI12/NET34_XI13/XI12/MM1_g N_VSS_XI13/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI12/MM9 N_XI13/XI12/NET36_XI13/XI12/MM9_d N_WL<23>_XI13/XI12/MM9_g
+ N_BL<3>_XI13/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI12/MM6 N_XI13/XI12/NET35_XI13/XI12/MM6_d
+ N_XI13/XI12/NET36_XI13/XI12/MM6_g N_VSS_XI13/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI12/MM7 N_XI13/XI12/NET36_XI13/XI12/MM7_d
+ N_XI13/XI12/NET35_XI13/XI12/MM7_g N_VSS_XI13/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI12/MM8 N_XI13/XI12/NET35_XI13/XI12/MM8_d N_WL<23>_XI13/XI12/MM8_g
+ N_BLN<3>_XI13/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI12/MM5 N_XI13/XI12/NET34_XI13/XI12/MM5_d
+ N_XI13/XI12/NET33_XI13/XI12/MM5_g N_VDD_XI13/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI12/MM4 N_XI13/XI12/NET33_XI13/XI12/MM4_d
+ N_XI13/XI12/NET34_XI13/XI12/MM4_g N_VDD_XI13/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI12/MM10 N_XI13/XI12/NET35_XI13/XI12/MM10_d
+ N_XI13/XI12/NET36_XI13/XI12/MM10_g N_VDD_XI13/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI12/MM11 N_XI13/XI12/NET36_XI13/XI12/MM11_d
+ N_XI13/XI12/NET35_XI13/XI12/MM11_g N_VDD_XI13/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI13/MM2 N_XI13/XI13/NET34_XI13/XI13/MM2_d
+ N_XI13/XI13/NET33_XI13/XI13/MM2_g N_VSS_XI13/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI13/MM3 N_XI13/XI13/NET33_XI13/XI13/MM3_d N_WL<22>_XI13/XI13/MM3_g
+ N_BLN<2>_XI13/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI13/MM0 N_XI13/XI13/NET34_XI13/XI13/MM0_d N_WL<22>_XI13/XI13/MM0_g
+ N_BL<2>_XI13/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI13/MM1 N_XI13/XI13/NET33_XI13/XI13/MM1_d
+ N_XI13/XI13/NET34_XI13/XI13/MM1_g N_VSS_XI13/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI13/MM9 N_XI13/XI13/NET36_XI13/XI13/MM9_d N_WL<23>_XI13/XI13/MM9_g
+ N_BL<2>_XI13/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI13/MM6 N_XI13/XI13/NET35_XI13/XI13/MM6_d
+ N_XI13/XI13/NET36_XI13/XI13/MM6_g N_VSS_XI13/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI13/MM7 N_XI13/XI13/NET36_XI13/XI13/MM7_d
+ N_XI13/XI13/NET35_XI13/XI13/MM7_g N_VSS_XI13/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI13/MM8 N_XI13/XI13/NET35_XI13/XI13/MM8_d N_WL<23>_XI13/XI13/MM8_g
+ N_BLN<2>_XI13/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI13/MM5 N_XI13/XI13/NET34_XI13/XI13/MM5_d
+ N_XI13/XI13/NET33_XI13/XI13/MM5_g N_VDD_XI13/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI13/MM4 N_XI13/XI13/NET33_XI13/XI13/MM4_d
+ N_XI13/XI13/NET34_XI13/XI13/MM4_g N_VDD_XI13/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI13/MM10 N_XI13/XI13/NET35_XI13/XI13/MM10_d
+ N_XI13/XI13/NET36_XI13/XI13/MM10_g N_VDD_XI13/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI13/MM11 N_XI13/XI13/NET36_XI13/XI13/MM11_d
+ N_XI13/XI13/NET35_XI13/XI13/MM11_g N_VDD_XI13/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI14/MM2 N_XI13/XI14/NET34_XI13/XI14/MM2_d
+ N_XI13/XI14/NET33_XI13/XI14/MM2_g N_VSS_XI13/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI14/MM3 N_XI13/XI14/NET33_XI13/XI14/MM3_d N_WL<22>_XI13/XI14/MM3_g
+ N_BLN<1>_XI13/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI14/MM0 N_XI13/XI14/NET34_XI13/XI14/MM0_d N_WL<22>_XI13/XI14/MM0_g
+ N_BL<1>_XI13/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI14/MM1 N_XI13/XI14/NET33_XI13/XI14/MM1_d
+ N_XI13/XI14/NET34_XI13/XI14/MM1_g N_VSS_XI13/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI14/MM9 N_XI13/XI14/NET36_XI13/XI14/MM9_d N_WL<23>_XI13/XI14/MM9_g
+ N_BL<1>_XI13/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI14/MM6 N_XI13/XI14/NET35_XI13/XI14/MM6_d
+ N_XI13/XI14/NET36_XI13/XI14/MM6_g N_VSS_XI13/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI14/MM7 N_XI13/XI14/NET36_XI13/XI14/MM7_d
+ N_XI13/XI14/NET35_XI13/XI14/MM7_g N_VSS_XI13/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI14/MM8 N_XI13/XI14/NET35_XI13/XI14/MM8_d N_WL<23>_XI13/XI14/MM8_g
+ N_BLN<1>_XI13/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI14/MM5 N_XI13/XI14/NET34_XI13/XI14/MM5_d
+ N_XI13/XI14/NET33_XI13/XI14/MM5_g N_VDD_XI13/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI14/MM4 N_XI13/XI14/NET33_XI13/XI14/MM4_d
+ N_XI13/XI14/NET34_XI13/XI14/MM4_g N_VDD_XI13/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI14/MM10 N_XI13/XI14/NET35_XI13/XI14/MM10_d
+ N_XI13/XI14/NET36_XI13/XI14/MM10_g N_VDD_XI13/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI14/MM11 N_XI13/XI14/NET36_XI13/XI14/MM11_d
+ N_XI13/XI14/NET35_XI13/XI14/MM11_g N_VDD_XI13/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI15/MM2 N_XI13/XI15/NET34_XI13/XI15/MM2_d
+ N_XI13/XI15/NET33_XI13/XI15/MM2_g N_VSS_XI13/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI15/MM3 N_XI13/XI15/NET33_XI13/XI15/MM3_d N_WL<22>_XI13/XI15/MM3_g
+ N_BLN<0>_XI13/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI15/MM0 N_XI13/XI15/NET34_XI13/XI15/MM0_d N_WL<22>_XI13/XI15/MM0_g
+ N_BL<0>_XI13/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI15/MM1 N_XI13/XI15/NET33_XI13/XI15/MM1_d
+ N_XI13/XI15/NET34_XI13/XI15/MM1_g N_VSS_XI13/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI15/MM9 N_XI13/XI15/NET36_XI13/XI15/MM9_d N_WL<23>_XI13/XI15/MM9_g
+ N_BL<0>_XI13/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI15/MM6 N_XI13/XI15/NET35_XI13/XI15/MM6_d
+ N_XI13/XI15/NET36_XI13/XI15/MM6_g N_VSS_XI13/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI15/MM7 N_XI13/XI15/NET36_XI13/XI15/MM7_d
+ N_XI13/XI15/NET35_XI13/XI15/MM7_g N_VSS_XI13/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/XI15/MM8 N_XI13/XI15/NET35_XI13/XI15/MM8_d N_WL<23>_XI13/XI15/MM8_g
+ N_BLN<0>_XI13/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI13/XI15/MM5 N_XI13/XI15/NET34_XI13/XI15/MM5_d
+ N_XI13/XI15/NET33_XI13/XI15/MM5_g N_VDD_XI13/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI15/MM4 N_XI13/XI15/NET33_XI13/XI15/MM4_d
+ N_XI13/XI15/NET34_XI13/XI15/MM4_g N_VDD_XI13/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI15/MM10 N_XI13/XI15/NET35_XI13/XI15/MM10_d
+ N_XI13/XI15/NET36_XI13/XI15/MM10_g N_VDD_XI13/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/XI15/MM11 N_XI13/XI15/NET36_XI13/XI15/MM11_d
+ N_XI13/XI15/NET35_XI13/XI15/MM11_g N_VDD_XI13/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI0/MM2 N_XI14/XI0/NET34_XI14/XI0/MM2_d N_XI14/XI0/NET33_XI14/XI0/MM2_g
+ N_VSS_XI14/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI0/MM3 N_XI14/XI0/NET33_XI14/XI0/MM3_d N_WL<24>_XI14/XI0/MM3_g
+ N_BLN<15>_XI14/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI0/MM0 N_XI14/XI0/NET34_XI14/XI0/MM0_d N_WL<24>_XI14/XI0/MM0_g
+ N_BL<15>_XI14/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI0/MM1 N_XI14/XI0/NET33_XI14/XI0/MM1_d N_XI14/XI0/NET34_XI14/XI0/MM1_g
+ N_VSS_XI14/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI0/MM9 N_XI14/XI0/NET36_XI14/XI0/MM9_d N_WL<25>_XI14/XI0/MM9_g
+ N_BL<15>_XI14/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI0/MM6 N_XI14/XI0/NET35_XI14/XI0/MM6_d N_XI14/XI0/NET36_XI14/XI0/MM6_g
+ N_VSS_XI14/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI0/MM7 N_XI14/XI0/NET36_XI14/XI0/MM7_d N_XI14/XI0/NET35_XI14/XI0/MM7_g
+ N_VSS_XI14/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI0/MM8 N_XI14/XI0/NET35_XI14/XI0/MM8_d N_WL<25>_XI14/XI0/MM8_g
+ N_BLN<15>_XI14/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI0/MM5 N_XI14/XI0/NET34_XI14/XI0/MM5_d N_XI14/XI0/NET33_XI14/XI0/MM5_g
+ N_VDD_XI14/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI0/MM4 N_XI14/XI0/NET33_XI14/XI0/MM4_d N_XI14/XI0/NET34_XI14/XI0/MM4_g
+ N_VDD_XI14/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI0/MM10 N_XI14/XI0/NET35_XI14/XI0/MM10_d N_XI14/XI0/NET36_XI14/XI0/MM10_g
+ N_VDD_XI14/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI0/MM11 N_XI14/XI0/NET36_XI14/XI0/MM11_d N_XI14/XI0/NET35_XI14/XI0/MM11_g
+ N_VDD_XI14/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI1/MM2 N_XI14/XI1/NET34_XI14/XI1/MM2_d N_XI14/XI1/NET33_XI14/XI1/MM2_g
+ N_VSS_XI14/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI1/MM3 N_XI14/XI1/NET33_XI14/XI1/MM3_d N_WL<24>_XI14/XI1/MM3_g
+ N_BLN<14>_XI14/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI1/MM0 N_XI14/XI1/NET34_XI14/XI1/MM0_d N_WL<24>_XI14/XI1/MM0_g
+ N_BL<14>_XI14/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI1/MM1 N_XI14/XI1/NET33_XI14/XI1/MM1_d N_XI14/XI1/NET34_XI14/XI1/MM1_g
+ N_VSS_XI14/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI1/MM9 N_XI14/XI1/NET36_XI14/XI1/MM9_d N_WL<25>_XI14/XI1/MM9_g
+ N_BL<14>_XI14/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI1/MM6 N_XI14/XI1/NET35_XI14/XI1/MM6_d N_XI14/XI1/NET36_XI14/XI1/MM6_g
+ N_VSS_XI14/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI1/MM7 N_XI14/XI1/NET36_XI14/XI1/MM7_d N_XI14/XI1/NET35_XI14/XI1/MM7_g
+ N_VSS_XI14/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI1/MM8 N_XI14/XI1/NET35_XI14/XI1/MM8_d N_WL<25>_XI14/XI1/MM8_g
+ N_BLN<14>_XI14/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI1/MM5 N_XI14/XI1/NET34_XI14/XI1/MM5_d N_XI14/XI1/NET33_XI14/XI1/MM5_g
+ N_VDD_XI14/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI1/MM4 N_XI14/XI1/NET33_XI14/XI1/MM4_d N_XI14/XI1/NET34_XI14/XI1/MM4_g
+ N_VDD_XI14/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI1/MM10 N_XI14/XI1/NET35_XI14/XI1/MM10_d N_XI14/XI1/NET36_XI14/XI1/MM10_g
+ N_VDD_XI14/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI1/MM11 N_XI14/XI1/NET36_XI14/XI1/MM11_d N_XI14/XI1/NET35_XI14/XI1/MM11_g
+ N_VDD_XI14/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI2/MM2 N_XI14/XI2/NET34_XI14/XI2/MM2_d N_XI14/XI2/NET33_XI14/XI2/MM2_g
+ N_VSS_XI14/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI2/MM3 N_XI14/XI2/NET33_XI14/XI2/MM3_d N_WL<24>_XI14/XI2/MM3_g
+ N_BLN<13>_XI14/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI2/MM0 N_XI14/XI2/NET34_XI14/XI2/MM0_d N_WL<24>_XI14/XI2/MM0_g
+ N_BL<13>_XI14/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI2/MM1 N_XI14/XI2/NET33_XI14/XI2/MM1_d N_XI14/XI2/NET34_XI14/XI2/MM1_g
+ N_VSS_XI14/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI2/MM9 N_XI14/XI2/NET36_XI14/XI2/MM9_d N_WL<25>_XI14/XI2/MM9_g
+ N_BL<13>_XI14/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI2/MM6 N_XI14/XI2/NET35_XI14/XI2/MM6_d N_XI14/XI2/NET36_XI14/XI2/MM6_g
+ N_VSS_XI14/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI2/MM7 N_XI14/XI2/NET36_XI14/XI2/MM7_d N_XI14/XI2/NET35_XI14/XI2/MM7_g
+ N_VSS_XI14/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI2/MM8 N_XI14/XI2/NET35_XI14/XI2/MM8_d N_WL<25>_XI14/XI2/MM8_g
+ N_BLN<13>_XI14/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI2/MM5 N_XI14/XI2/NET34_XI14/XI2/MM5_d N_XI14/XI2/NET33_XI14/XI2/MM5_g
+ N_VDD_XI14/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI2/MM4 N_XI14/XI2/NET33_XI14/XI2/MM4_d N_XI14/XI2/NET34_XI14/XI2/MM4_g
+ N_VDD_XI14/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI2/MM10 N_XI14/XI2/NET35_XI14/XI2/MM10_d N_XI14/XI2/NET36_XI14/XI2/MM10_g
+ N_VDD_XI14/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI2/MM11 N_XI14/XI2/NET36_XI14/XI2/MM11_d N_XI14/XI2/NET35_XI14/XI2/MM11_g
+ N_VDD_XI14/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI3/MM2 N_XI14/XI3/NET34_XI14/XI3/MM2_d N_XI14/XI3/NET33_XI14/XI3/MM2_g
+ N_VSS_XI14/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI3/MM3 N_XI14/XI3/NET33_XI14/XI3/MM3_d N_WL<24>_XI14/XI3/MM3_g
+ N_BLN<12>_XI14/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI3/MM0 N_XI14/XI3/NET34_XI14/XI3/MM0_d N_WL<24>_XI14/XI3/MM0_g
+ N_BL<12>_XI14/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI3/MM1 N_XI14/XI3/NET33_XI14/XI3/MM1_d N_XI14/XI3/NET34_XI14/XI3/MM1_g
+ N_VSS_XI14/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI3/MM9 N_XI14/XI3/NET36_XI14/XI3/MM9_d N_WL<25>_XI14/XI3/MM9_g
+ N_BL<12>_XI14/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI3/MM6 N_XI14/XI3/NET35_XI14/XI3/MM6_d N_XI14/XI3/NET36_XI14/XI3/MM6_g
+ N_VSS_XI14/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI3/MM7 N_XI14/XI3/NET36_XI14/XI3/MM7_d N_XI14/XI3/NET35_XI14/XI3/MM7_g
+ N_VSS_XI14/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI3/MM8 N_XI14/XI3/NET35_XI14/XI3/MM8_d N_WL<25>_XI14/XI3/MM8_g
+ N_BLN<12>_XI14/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI3/MM5 N_XI14/XI3/NET34_XI14/XI3/MM5_d N_XI14/XI3/NET33_XI14/XI3/MM5_g
+ N_VDD_XI14/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI3/MM4 N_XI14/XI3/NET33_XI14/XI3/MM4_d N_XI14/XI3/NET34_XI14/XI3/MM4_g
+ N_VDD_XI14/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI3/MM10 N_XI14/XI3/NET35_XI14/XI3/MM10_d N_XI14/XI3/NET36_XI14/XI3/MM10_g
+ N_VDD_XI14/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI3/MM11 N_XI14/XI3/NET36_XI14/XI3/MM11_d N_XI14/XI3/NET35_XI14/XI3/MM11_g
+ N_VDD_XI14/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI4/MM2 N_XI14/XI4/NET34_XI14/XI4/MM2_d N_XI14/XI4/NET33_XI14/XI4/MM2_g
+ N_VSS_XI14/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI4/MM3 N_XI14/XI4/NET33_XI14/XI4/MM3_d N_WL<24>_XI14/XI4/MM3_g
+ N_BLN<11>_XI14/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI4/MM0 N_XI14/XI4/NET34_XI14/XI4/MM0_d N_WL<24>_XI14/XI4/MM0_g
+ N_BL<11>_XI14/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI4/MM1 N_XI14/XI4/NET33_XI14/XI4/MM1_d N_XI14/XI4/NET34_XI14/XI4/MM1_g
+ N_VSS_XI14/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI4/MM9 N_XI14/XI4/NET36_XI14/XI4/MM9_d N_WL<25>_XI14/XI4/MM9_g
+ N_BL<11>_XI14/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI4/MM6 N_XI14/XI4/NET35_XI14/XI4/MM6_d N_XI14/XI4/NET36_XI14/XI4/MM6_g
+ N_VSS_XI14/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI4/MM7 N_XI14/XI4/NET36_XI14/XI4/MM7_d N_XI14/XI4/NET35_XI14/XI4/MM7_g
+ N_VSS_XI14/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI4/MM8 N_XI14/XI4/NET35_XI14/XI4/MM8_d N_WL<25>_XI14/XI4/MM8_g
+ N_BLN<11>_XI14/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI4/MM5 N_XI14/XI4/NET34_XI14/XI4/MM5_d N_XI14/XI4/NET33_XI14/XI4/MM5_g
+ N_VDD_XI14/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI4/MM4 N_XI14/XI4/NET33_XI14/XI4/MM4_d N_XI14/XI4/NET34_XI14/XI4/MM4_g
+ N_VDD_XI14/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI4/MM10 N_XI14/XI4/NET35_XI14/XI4/MM10_d N_XI14/XI4/NET36_XI14/XI4/MM10_g
+ N_VDD_XI14/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI4/MM11 N_XI14/XI4/NET36_XI14/XI4/MM11_d N_XI14/XI4/NET35_XI14/XI4/MM11_g
+ N_VDD_XI14/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI5/MM2 N_XI14/XI5/NET34_XI14/XI5/MM2_d N_XI14/XI5/NET33_XI14/XI5/MM2_g
+ N_VSS_XI14/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI5/MM3 N_XI14/XI5/NET33_XI14/XI5/MM3_d N_WL<24>_XI14/XI5/MM3_g
+ N_BLN<10>_XI14/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI5/MM0 N_XI14/XI5/NET34_XI14/XI5/MM0_d N_WL<24>_XI14/XI5/MM0_g
+ N_BL<10>_XI14/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI5/MM1 N_XI14/XI5/NET33_XI14/XI5/MM1_d N_XI14/XI5/NET34_XI14/XI5/MM1_g
+ N_VSS_XI14/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI5/MM9 N_XI14/XI5/NET36_XI14/XI5/MM9_d N_WL<25>_XI14/XI5/MM9_g
+ N_BL<10>_XI14/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI5/MM6 N_XI14/XI5/NET35_XI14/XI5/MM6_d N_XI14/XI5/NET36_XI14/XI5/MM6_g
+ N_VSS_XI14/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI5/MM7 N_XI14/XI5/NET36_XI14/XI5/MM7_d N_XI14/XI5/NET35_XI14/XI5/MM7_g
+ N_VSS_XI14/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI5/MM8 N_XI14/XI5/NET35_XI14/XI5/MM8_d N_WL<25>_XI14/XI5/MM8_g
+ N_BLN<10>_XI14/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI5/MM5 N_XI14/XI5/NET34_XI14/XI5/MM5_d N_XI14/XI5/NET33_XI14/XI5/MM5_g
+ N_VDD_XI14/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI5/MM4 N_XI14/XI5/NET33_XI14/XI5/MM4_d N_XI14/XI5/NET34_XI14/XI5/MM4_g
+ N_VDD_XI14/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI5/MM10 N_XI14/XI5/NET35_XI14/XI5/MM10_d N_XI14/XI5/NET36_XI14/XI5/MM10_g
+ N_VDD_XI14/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI5/MM11 N_XI14/XI5/NET36_XI14/XI5/MM11_d N_XI14/XI5/NET35_XI14/XI5/MM11_g
+ N_VDD_XI14/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI6/MM2 N_XI14/XI6/NET34_XI14/XI6/MM2_d N_XI14/XI6/NET33_XI14/XI6/MM2_g
+ N_VSS_XI14/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM3 N_XI14/XI6/NET33_XI14/XI6/MM3_d N_WL<24>_XI14/XI6/MM3_g
+ N_BLN<9>_XI14/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM0 N_XI14/XI6/NET34_XI14/XI6/MM0_d N_WL<24>_XI14/XI6/MM0_g
+ N_BL<9>_XI14/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM1 N_XI14/XI6/NET33_XI14/XI6/MM1_d N_XI14/XI6/NET34_XI14/XI6/MM1_g
+ N_VSS_XI14/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM9 N_XI14/XI6/NET36_XI14/XI6/MM9_d N_WL<25>_XI14/XI6/MM9_g
+ N_BL<9>_XI14/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM6 N_XI14/XI6/NET35_XI14/XI6/MM6_d N_XI14/XI6/NET36_XI14/XI6/MM6_g
+ N_VSS_XI14/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM7 N_XI14/XI6/NET36_XI14/XI6/MM7_d N_XI14/XI6/NET35_XI14/XI6/MM7_g
+ N_VSS_XI14/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM8 N_XI14/XI6/NET35_XI14/XI6/MM8_d N_WL<25>_XI14/XI6/MM8_g
+ N_BLN<9>_XI14/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI6/MM5 N_XI14/XI6/NET34_XI14/XI6/MM5_d N_XI14/XI6/NET33_XI14/XI6/MM5_g
+ N_VDD_XI14/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI6/MM4 N_XI14/XI6/NET33_XI14/XI6/MM4_d N_XI14/XI6/NET34_XI14/XI6/MM4_g
+ N_VDD_XI14/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI6/MM10 N_XI14/XI6/NET35_XI14/XI6/MM10_d N_XI14/XI6/NET36_XI14/XI6/MM10_g
+ N_VDD_XI14/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI6/MM11 N_XI14/XI6/NET36_XI14/XI6/MM11_d N_XI14/XI6/NET35_XI14/XI6/MM11_g
+ N_VDD_XI14/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI7/MM2 N_XI14/XI7/NET34_XI14/XI7/MM2_d N_XI14/XI7/NET33_XI14/XI7/MM2_g
+ N_VSS_XI14/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM3 N_XI14/XI7/NET33_XI14/XI7/MM3_d N_WL<24>_XI14/XI7/MM3_g
+ N_BLN<8>_XI14/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM0 N_XI14/XI7/NET34_XI14/XI7/MM0_d N_WL<24>_XI14/XI7/MM0_g
+ N_BL<8>_XI14/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM1 N_XI14/XI7/NET33_XI14/XI7/MM1_d N_XI14/XI7/NET34_XI14/XI7/MM1_g
+ N_VSS_XI14/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM9 N_XI14/XI7/NET36_XI14/XI7/MM9_d N_WL<25>_XI14/XI7/MM9_g
+ N_BL<8>_XI14/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM6 N_XI14/XI7/NET35_XI14/XI7/MM6_d N_XI14/XI7/NET36_XI14/XI7/MM6_g
+ N_VSS_XI14/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM7 N_XI14/XI7/NET36_XI14/XI7/MM7_d N_XI14/XI7/NET35_XI14/XI7/MM7_g
+ N_VSS_XI14/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM8 N_XI14/XI7/NET35_XI14/XI7/MM8_d N_WL<25>_XI14/XI7/MM8_g
+ N_BLN<8>_XI14/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI7/MM5 N_XI14/XI7/NET34_XI14/XI7/MM5_d N_XI14/XI7/NET33_XI14/XI7/MM5_g
+ N_VDD_XI14/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI7/MM4 N_XI14/XI7/NET33_XI14/XI7/MM4_d N_XI14/XI7/NET34_XI14/XI7/MM4_g
+ N_VDD_XI14/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI7/MM10 N_XI14/XI7/NET35_XI14/XI7/MM10_d N_XI14/XI7/NET36_XI14/XI7/MM10_g
+ N_VDD_XI14/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI7/MM11 N_XI14/XI7/NET36_XI14/XI7/MM11_d N_XI14/XI7/NET35_XI14/XI7/MM11_g
+ N_VDD_XI14/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI8/MM2 N_XI14/XI8/NET34_XI14/XI8/MM2_d N_XI14/XI8/NET33_XI14/XI8/MM2_g
+ N_VSS_XI14/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM3 N_XI14/XI8/NET33_XI14/XI8/MM3_d N_WL<24>_XI14/XI8/MM3_g
+ N_BLN<7>_XI14/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM0 N_XI14/XI8/NET34_XI14/XI8/MM0_d N_WL<24>_XI14/XI8/MM0_g
+ N_BL<7>_XI14/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM1 N_XI14/XI8/NET33_XI14/XI8/MM1_d N_XI14/XI8/NET34_XI14/XI8/MM1_g
+ N_VSS_XI14/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM9 N_XI14/XI8/NET36_XI14/XI8/MM9_d N_WL<25>_XI14/XI8/MM9_g
+ N_BL<7>_XI14/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM6 N_XI14/XI8/NET35_XI14/XI8/MM6_d N_XI14/XI8/NET36_XI14/XI8/MM6_g
+ N_VSS_XI14/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM7 N_XI14/XI8/NET36_XI14/XI8/MM7_d N_XI14/XI8/NET35_XI14/XI8/MM7_g
+ N_VSS_XI14/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM8 N_XI14/XI8/NET35_XI14/XI8/MM8_d N_WL<25>_XI14/XI8/MM8_g
+ N_BLN<7>_XI14/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI8/MM5 N_XI14/XI8/NET34_XI14/XI8/MM5_d N_XI14/XI8/NET33_XI14/XI8/MM5_g
+ N_VDD_XI14/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI8/MM4 N_XI14/XI8/NET33_XI14/XI8/MM4_d N_XI14/XI8/NET34_XI14/XI8/MM4_g
+ N_VDD_XI14/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI8/MM10 N_XI14/XI8/NET35_XI14/XI8/MM10_d N_XI14/XI8/NET36_XI14/XI8/MM10_g
+ N_VDD_XI14/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI8/MM11 N_XI14/XI8/NET36_XI14/XI8/MM11_d N_XI14/XI8/NET35_XI14/XI8/MM11_g
+ N_VDD_XI14/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI9/MM2 N_XI14/XI9/NET34_XI14/XI9/MM2_d N_XI14/XI9/NET33_XI14/XI9/MM2_g
+ N_VSS_XI14/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM3 N_XI14/XI9/NET33_XI14/XI9/MM3_d N_WL<24>_XI14/XI9/MM3_g
+ N_BLN<6>_XI14/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM0 N_XI14/XI9/NET34_XI14/XI9/MM0_d N_WL<24>_XI14/XI9/MM0_g
+ N_BL<6>_XI14/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM1 N_XI14/XI9/NET33_XI14/XI9/MM1_d N_XI14/XI9/NET34_XI14/XI9/MM1_g
+ N_VSS_XI14/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM9 N_XI14/XI9/NET36_XI14/XI9/MM9_d N_WL<25>_XI14/XI9/MM9_g
+ N_BL<6>_XI14/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM6 N_XI14/XI9/NET35_XI14/XI9/MM6_d N_XI14/XI9/NET36_XI14/XI9/MM6_g
+ N_VSS_XI14/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM7 N_XI14/XI9/NET36_XI14/XI9/MM7_d N_XI14/XI9/NET35_XI14/XI9/MM7_g
+ N_VSS_XI14/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM8 N_XI14/XI9/NET35_XI14/XI9/MM8_d N_WL<25>_XI14/XI9/MM8_g
+ N_BLN<6>_XI14/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI9/MM5 N_XI14/XI9/NET34_XI14/XI9/MM5_d N_XI14/XI9/NET33_XI14/XI9/MM5_g
+ N_VDD_XI14/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI9/MM4 N_XI14/XI9/NET33_XI14/XI9/MM4_d N_XI14/XI9/NET34_XI14/XI9/MM4_g
+ N_VDD_XI14/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI9/MM10 N_XI14/XI9/NET35_XI14/XI9/MM10_d N_XI14/XI9/NET36_XI14/XI9/MM10_g
+ N_VDD_XI14/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI9/MM11 N_XI14/XI9/NET36_XI14/XI9/MM11_d N_XI14/XI9/NET35_XI14/XI9/MM11_g
+ N_VDD_XI14/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI10/MM2 N_XI14/XI10/NET34_XI14/XI10/MM2_d
+ N_XI14/XI10/NET33_XI14/XI10/MM2_g N_VSS_XI14/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI10/MM3 N_XI14/XI10/NET33_XI14/XI10/MM3_d N_WL<24>_XI14/XI10/MM3_g
+ N_BLN<5>_XI14/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI10/MM0 N_XI14/XI10/NET34_XI14/XI10/MM0_d N_WL<24>_XI14/XI10/MM0_g
+ N_BL<5>_XI14/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI10/MM1 N_XI14/XI10/NET33_XI14/XI10/MM1_d
+ N_XI14/XI10/NET34_XI14/XI10/MM1_g N_VSS_XI14/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI10/MM9 N_XI14/XI10/NET36_XI14/XI10/MM9_d N_WL<25>_XI14/XI10/MM9_g
+ N_BL<5>_XI14/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI10/MM6 N_XI14/XI10/NET35_XI14/XI10/MM6_d
+ N_XI14/XI10/NET36_XI14/XI10/MM6_g N_VSS_XI14/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI10/MM7 N_XI14/XI10/NET36_XI14/XI10/MM7_d
+ N_XI14/XI10/NET35_XI14/XI10/MM7_g N_VSS_XI14/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI10/MM8 N_XI14/XI10/NET35_XI14/XI10/MM8_d N_WL<25>_XI14/XI10/MM8_g
+ N_BLN<5>_XI14/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI10/MM5 N_XI14/XI10/NET34_XI14/XI10/MM5_d
+ N_XI14/XI10/NET33_XI14/XI10/MM5_g N_VDD_XI14/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI10/MM4 N_XI14/XI10/NET33_XI14/XI10/MM4_d
+ N_XI14/XI10/NET34_XI14/XI10/MM4_g N_VDD_XI14/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI10/MM10 N_XI14/XI10/NET35_XI14/XI10/MM10_d
+ N_XI14/XI10/NET36_XI14/XI10/MM10_g N_VDD_XI14/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI10/MM11 N_XI14/XI10/NET36_XI14/XI10/MM11_d
+ N_XI14/XI10/NET35_XI14/XI10/MM11_g N_VDD_XI14/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI11/MM2 N_XI14/XI11/NET34_XI14/XI11/MM2_d
+ N_XI14/XI11/NET33_XI14/XI11/MM2_g N_VSS_XI14/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI11/MM3 N_XI14/XI11/NET33_XI14/XI11/MM3_d N_WL<24>_XI14/XI11/MM3_g
+ N_BLN<4>_XI14/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI11/MM0 N_XI14/XI11/NET34_XI14/XI11/MM0_d N_WL<24>_XI14/XI11/MM0_g
+ N_BL<4>_XI14/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI11/MM1 N_XI14/XI11/NET33_XI14/XI11/MM1_d
+ N_XI14/XI11/NET34_XI14/XI11/MM1_g N_VSS_XI14/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI11/MM9 N_XI14/XI11/NET36_XI14/XI11/MM9_d N_WL<25>_XI14/XI11/MM9_g
+ N_BL<4>_XI14/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI11/MM6 N_XI14/XI11/NET35_XI14/XI11/MM6_d
+ N_XI14/XI11/NET36_XI14/XI11/MM6_g N_VSS_XI14/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI11/MM7 N_XI14/XI11/NET36_XI14/XI11/MM7_d
+ N_XI14/XI11/NET35_XI14/XI11/MM7_g N_VSS_XI14/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI11/MM8 N_XI14/XI11/NET35_XI14/XI11/MM8_d N_WL<25>_XI14/XI11/MM8_g
+ N_BLN<4>_XI14/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI11/MM5 N_XI14/XI11/NET34_XI14/XI11/MM5_d
+ N_XI14/XI11/NET33_XI14/XI11/MM5_g N_VDD_XI14/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI11/MM4 N_XI14/XI11/NET33_XI14/XI11/MM4_d
+ N_XI14/XI11/NET34_XI14/XI11/MM4_g N_VDD_XI14/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI11/MM10 N_XI14/XI11/NET35_XI14/XI11/MM10_d
+ N_XI14/XI11/NET36_XI14/XI11/MM10_g N_VDD_XI14/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI11/MM11 N_XI14/XI11/NET36_XI14/XI11/MM11_d
+ N_XI14/XI11/NET35_XI14/XI11/MM11_g N_VDD_XI14/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI12/MM2 N_XI14/XI12/NET34_XI14/XI12/MM2_d
+ N_XI14/XI12/NET33_XI14/XI12/MM2_g N_VSS_XI14/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI12/MM3 N_XI14/XI12/NET33_XI14/XI12/MM3_d N_WL<24>_XI14/XI12/MM3_g
+ N_BLN<3>_XI14/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI12/MM0 N_XI14/XI12/NET34_XI14/XI12/MM0_d N_WL<24>_XI14/XI12/MM0_g
+ N_BL<3>_XI14/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI12/MM1 N_XI14/XI12/NET33_XI14/XI12/MM1_d
+ N_XI14/XI12/NET34_XI14/XI12/MM1_g N_VSS_XI14/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI12/MM9 N_XI14/XI12/NET36_XI14/XI12/MM9_d N_WL<25>_XI14/XI12/MM9_g
+ N_BL<3>_XI14/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI12/MM6 N_XI14/XI12/NET35_XI14/XI12/MM6_d
+ N_XI14/XI12/NET36_XI14/XI12/MM6_g N_VSS_XI14/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI12/MM7 N_XI14/XI12/NET36_XI14/XI12/MM7_d
+ N_XI14/XI12/NET35_XI14/XI12/MM7_g N_VSS_XI14/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI12/MM8 N_XI14/XI12/NET35_XI14/XI12/MM8_d N_WL<25>_XI14/XI12/MM8_g
+ N_BLN<3>_XI14/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI12/MM5 N_XI14/XI12/NET34_XI14/XI12/MM5_d
+ N_XI14/XI12/NET33_XI14/XI12/MM5_g N_VDD_XI14/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI12/MM4 N_XI14/XI12/NET33_XI14/XI12/MM4_d
+ N_XI14/XI12/NET34_XI14/XI12/MM4_g N_VDD_XI14/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI12/MM10 N_XI14/XI12/NET35_XI14/XI12/MM10_d
+ N_XI14/XI12/NET36_XI14/XI12/MM10_g N_VDD_XI14/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI12/MM11 N_XI14/XI12/NET36_XI14/XI12/MM11_d
+ N_XI14/XI12/NET35_XI14/XI12/MM11_g N_VDD_XI14/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI13/MM2 N_XI14/XI13/NET34_XI14/XI13/MM2_d
+ N_XI14/XI13/NET33_XI14/XI13/MM2_g N_VSS_XI14/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI13/MM3 N_XI14/XI13/NET33_XI14/XI13/MM3_d N_WL<24>_XI14/XI13/MM3_g
+ N_BLN<2>_XI14/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI13/MM0 N_XI14/XI13/NET34_XI14/XI13/MM0_d N_WL<24>_XI14/XI13/MM0_g
+ N_BL<2>_XI14/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI13/MM1 N_XI14/XI13/NET33_XI14/XI13/MM1_d
+ N_XI14/XI13/NET34_XI14/XI13/MM1_g N_VSS_XI14/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI13/MM9 N_XI14/XI13/NET36_XI14/XI13/MM9_d N_WL<25>_XI14/XI13/MM9_g
+ N_BL<2>_XI14/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI13/MM6 N_XI14/XI13/NET35_XI14/XI13/MM6_d
+ N_XI14/XI13/NET36_XI14/XI13/MM6_g N_VSS_XI14/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI13/MM7 N_XI14/XI13/NET36_XI14/XI13/MM7_d
+ N_XI14/XI13/NET35_XI14/XI13/MM7_g N_VSS_XI14/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI13/MM8 N_XI14/XI13/NET35_XI14/XI13/MM8_d N_WL<25>_XI14/XI13/MM8_g
+ N_BLN<2>_XI14/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI13/MM5 N_XI14/XI13/NET34_XI14/XI13/MM5_d
+ N_XI14/XI13/NET33_XI14/XI13/MM5_g N_VDD_XI14/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI13/MM4 N_XI14/XI13/NET33_XI14/XI13/MM4_d
+ N_XI14/XI13/NET34_XI14/XI13/MM4_g N_VDD_XI14/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI13/MM10 N_XI14/XI13/NET35_XI14/XI13/MM10_d
+ N_XI14/XI13/NET36_XI14/XI13/MM10_g N_VDD_XI14/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI13/MM11 N_XI14/XI13/NET36_XI14/XI13/MM11_d
+ N_XI14/XI13/NET35_XI14/XI13/MM11_g N_VDD_XI14/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI14/MM2 N_XI14/XI14/NET34_XI14/XI14/MM2_d
+ N_XI14/XI14/NET33_XI14/XI14/MM2_g N_VSS_XI14/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI14/MM3 N_XI14/XI14/NET33_XI14/XI14/MM3_d N_WL<24>_XI14/XI14/MM3_g
+ N_BLN<1>_XI14/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI14/MM0 N_XI14/XI14/NET34_XI14/XI14/MM0_d N_WL<24>_XI14/XI14/MM0_g
+ N_BL<1>_XI14/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI14/MM1 N_XI14/XI14/NET33_XI14/XI14/MM1_d
+ N_XI14/XI14/NET34_XI14/XI14/MM1_g N_VSS_XI14/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI14/MM9 N_XI14/XI14/NET36_XI14/XI14/MM9_d N_WL<25>_XI14/XI14/MM9_g
+ N_BL<1>_XI14/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI14/MM6 N_XI14/XI14/NET35_XI14/XI14/MM6_d
+ N_XI14/XI14/NET36_XI14/XI14/MM6_g N_VSS_XI14/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI14/MM7 N_XI14/XI14/NET36_XI14/XI14/MM7_d
+ N_XI14/XI14/NET35_XI14/XI14/MM7_g N_VSS_XI14/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI14/MM8 N_XI14/XI14/NET35_XI14/XI14/MM8_d N_WL<25>_XI14/XI14/MM8_g
+ N_BLN<1>_XI14/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI14/MM5 N_XI14/XI14/NET34_XI14/XI14/MM5_d
+ N_XI14/XI14/NET33_XI14/XI14/MM5_g N_VDD_XI14/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI14/MM4 N_XI14/XI14/NET33_XI14/XI14/MM4_d
+ N_XI14/XI14/NET34_XI14/XI14/MM4_g N_VDD_XI14/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI14/MM10 N_XI14/XI14/NET35_XI14/XI14/MM10_d
+ N_XI14/XI14/NET36_XI14/XI14/MM10_g N_VDD_XI14/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI14/MM11 N_XI14/XI14/NET36_XI14/XI14/MM11_d
+ N_XI14/XI14/NET35_XI14/XI14/MM11_g N_VDD_XI14/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI15/MM2 N_XI14/XI15/NET34_XI14/XI15/MM2_d
+ N_XI14/XI15/NET33_XI14/XI15/MM2_g N_VSS_XI14/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI15/MM3 N_XI14/XI15/NET33_XI14/XI15/MM3_d N_WL<24>_XI14/XI15/MM3_g
+ N_BLN<0>_XI14/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI15/MM0 N_XI14/XI15/NET34_XI14/XI15/MM0_d N_WL<24>_XI14/XI15/MM0_g
+ N_BL<0>_XI14/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI15/MM1 N_XI14/XI15/NET33_XI14/XI15/MM1_d
+ N_XI14/XI15/NET34_XI14/XI15/MM1_g N_VSS_XI14/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI15/MM9 N_XI14/XI15/NET36_XI14/XI15/MM9_d N_WL<25>_XI14/XI15/MM9_g
+ N_BL<0>_XI14/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI15/MM6 N_XI14/XI15/NET35_XI14/XI15/MM6_d
+ N_XI14/XI15/NET36_XI14/XI15/MM6_g N_VSS_XI14/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI15/MM7 N_XI14/XI15/NET36_XI14/XI15/MM7_d
+ N_XI14/XI15/NET35_XI14/XI15/MM7_g N_VSS_XI14/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/XI15/MM8 N_XI14/XI15/NET35_XI14/XI15/MM8_d N_WL<25>_XI14/XI15/MM8_g
+ N_BLN<0>_XI14/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI14/XI15/MM5 N_XI14/XI15/NET34_XI14/XI15/MM5_d
+ N_XI14/XI15/NET33_XI14/XI15/MM5_g N_VDD_XI14/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI15/MM4 N_XI14/XI15/NET33_XI14/XI15/MM4_d
+ N_XI14/XI15/NET34_XI14/XI15/MM4_g N_VDD_XI14/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI15/MM10 N_XI14/XI15/NET35_XI14/XI15/MM10_d
+ N_XI14/XI15/NET36_XI14/XI15/MM10_g N_VDD_XI14/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/XI15/MM11 N_XI14/XI15/NET36_XI14/XI15/MM11_d
+ N_XI14/XI15/NET35_XI14/XI15/MM11_g N_VDD_XI14/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI0/MM2 N_XI15/XI0/NET34_XI15/XI0/MM2_d N_XI15/XI0/NET33_XI15/XI0/MM2_g
+ N_VSS_XI15/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI0/MM3 N_XI15/XI0/NET33_XI15/XI0/MM3_d N_WL<26>_XI15/XI0/MM3_g
+ N_BLN<15>_XI15/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI0/MM0 N_XI15/XI0/NET34_XI15/XI0/MM0_d N_WL<26>_XI15/XI0/MM0_g
+ N_BL<15>_XI15/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI0/MM1 N_XI15/XI0/NET33_XI15/XI0/MM1_d N_XI15/XI0/NET34_XI15/XI0/MM1_g
+ N_VSS_XI15/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI0/MM9 N_XI15/XI0/NET36_XI15/XI0/MM9_d N_WL<27>_XI15/XI0/MM9_g
+ N_BL<15>_XI15/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI0/MM6 N_XI15/XI0/NET35_XI15/XI0/MM6_d N_XI15/XI0/NET36_XI15/XI0/MM6_g
+ N_VSS_XI15/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI0/MM7 N_XI15/XI0/NET36_XI15/XI0/MM7_d N_XI15/XI0/NET35_XI15/XI0/MM7_g
+ N_VSS_XI15/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI0/MM8 N_XI15/XI0/NET35_XI15/XI0/MM8_d N_WL<27>_XI15/XI0/MM8_g
+ N_BLN<15>_XI15/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI0/MM5 N_XI15/XI0/NET34_XI15/XI0/MM5_d N_XI15/XI0/NET33_XI15/XI0/MM5_g
+ N_VDD_XI15/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI0/MM4 N_XI15/XI0/NET33_XI15/XI0/MM4_d N_XI15/XI0/NET34_XI15/XI0/MM4_g
+ N_VDD_XI15/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI0/MM10 N_XI15/XI0/NET35_XI15/XI0/MM10_d N_XI15/XI0/NET36_XI15/XI0/MM10_g
+ N_VDD_XI15/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI0/MM11 N_XI15/XI0/NET36_XI15/XI0/MM11_d N_XI15/XI0/NET35_XI15/XI0/MM11_g
+ N_VDD_XI15/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI1/MM2 N_XI15/XI1/NET34_XI15/XI1/MM2_d N_XI15/XI1/NET33_XI15/XI1/MM2_g
+ N_VSS_XI15/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI1/MM3 N_XI15/XI1/NET33_XI15/XI1/MM3_d N_WL<26>_XI15/XI1/MM3_g
+ N_BLN<14>_XI15/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI1/MM0 N_XI15/XI1/NET34_XI15/XI1/MM0_d N_WL<26>_XI15/XI1/MM0_g
+ N_BL<14>_XI15/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI1/MM1 N_XI15/XI1/NET33_XI15/XI1/MM1_d N_XI15/XI1/NET34_XI15/XI1/MM1_g
+ N_VSS_XI15/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI1/MM9 N_XI15/XI1/NET36_XI15/XI1/MM9_d N_WL<27>_XI15/XI1/MM9_g
+ N_BL<14>_XI15/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI1/MM6 N_XI15/XI1/NET35_XI15/XI1/MM6_d N_XI15/XI1/NET36_XI15/XI1/MM6_g
+ N_VSS_XI15/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI1/MM7 N_XI15/XI1/NET36_XI15/XI1/MM7_d N_XI15/XI1/NET35_XI15/XI1/MM7_g
+ N_VSS_XI15/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI1/MM8 N_XI15/XI1/NET35_XI15/XI1/MM8_d N_WL<27>_XI15/XI1/MM8_g
+ N_BLN<14>_XI15/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI1/MM5 N_XI15/XI1/NET34_XI15/XI1/MM5_d N_XI15/XI1/NET33_XI15/XI1/MM5_g
+ N_VDD_XI15/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI1/MM4 N_XI15/XI1/NET33_XI15/XI1/MM4_d N_XI15/XI1/NET34_XI15/XI1/MM4_g
+ N_VDD_XI15/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI1/MM10 N_XI15/XI1/NET35_XI15/XI1/MM10_d N_XI15/XI1/NET36_XI15/XI1/MM10_g
+ N_VDD_XI15/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI1/MM11 N_XI15/XI1/NET36_XI15/XI1/MM11_d N_XI15/XI1/NET35_XI15/XI1/MM11_g
+ N_VDD_XI15/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI2/MM2 N_XI15/XI2/NET34_XI15/XI2/MM2_d N_XI15/XI2/NET33_XI15/XI2/MM2_g
+ N_VSS_XI15/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI2/MM3 N_XI15/XI2/NET33_XI15/XI2/MM3_d N_WL<26>_XI15/XI2/MM3_g
+ N_BLN<13>_XI15/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI2/MM0 N_XI15/XI2/NET34_XI15/XI2/MM0_d N_WL<26>_XI15/XI2/MM0_g
+ N_BL<13>_XI15/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI2/MM1 N_XI15/XI2/NET33_XI15/XI2/MM1_d N_XI15/XI2/NET34_XI15/XI2/MM1_g
+ N_VSS_XI15/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI2/MM9 N_XI15/XI2/NET36_XI15/XI2/MM9_d N_WL<27>_XI15/XI2/MM9_g
+ N_BL<13>_XI15/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI2/MM6 N_XI15/XI2/NET35_XI15/XI2/MM6_d N_XI15/XI2/NET36_XI15/XI2/MM6_g
+ N_VSS_XI15/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI2/MM7 N_XI15/XI2/NET36_XI15/XI2/MM7_d N_XI15/XI2/NET35_XI15/XI2/MM7_g
+ N_VSS_XI15/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI2/MM8 N_XI15/XI2/NET35_XI15/XI2/MM8_d N_WL<27>_XI15/XI2/MM8_g
+ N_BLN<13>_XI15/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI2/MM5 N_XI15/XI2/NET34_XI15/XI2/MM5_d N_XI15/XI2/NET33_XI15/XI2/MM5_g
+ N_VDD_XI15/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI2/MM4 N_XI15/XI2/NET33_XI15/XI2/MM4_d N_XI15/XI2/NET34_XI15/XI2/MM4_g
+ N_VDD_XI15/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI2/MM10 N_XI15/XI2/NET35_XI15/XI2/MM10_d N_XI15/XI2/NET36_XI15/XI2/MM10_g
+ N_VDD_XI15/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI2/MM11 N_XI15/XI2/NET36_XI15/XI2/MM11_d N_XI15/XI2/NET35_XI15/XI2/MM11_g
+ N_VDD_XI15/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI3/MM2 N_XI15/XI3/NET34_XI15/XI3/MM2_d N_XI15/XI3/NET33_XI15/XI3/MM2_g
+ N_VSS_XI15/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI3/MM3 N_XI15/XI3/NET33_XI15/XI3/MM3_d N_WL<26>_XI15/XI3/MM3_g
+ N_BLN<12>_XI15/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI3/MM0 N_XI15/XI3/NET34_XI15/XI3/MM0_d N_WL<26>_XI15/XI3/MM0_g
+ N_BL<12>_XI15/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI3/MM1 N_XI15/XI3/NET33_XI15/XI3/MM1_d N_XI15/XI3/NET34_XI15/XI3/MM1_g
+ N_VSS_XI15/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI3/MM9 N_XI15/XI3/NET36_XI15/XI3/MM9_d N_WL<27>_XI15/XI3/MM9_g
+ N_BL<12>_XI15/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI3/MM6 N_XI15/XI3/NET35_XI15/XI3/MM6_d N_XI15/XI3/NET36_XI15/XI3/MM6_g
+ N_VSS_XI15/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI3/MM7 N_XI15/XI3/NET36_XI15/XI3/MM7_d N_XI15/XI3/NET35_XI15/XI3/MM7_g
+ N_VSS_XI15/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI3/MM8 N_XI15/XI3/NET35_XI15/XI3/MM8_d N_WL<27>_XI15/XI3/MM8_g
+ N_BLN<12>_XI15/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI3/MM5 N_XI15/XI3/NET34_XI15/XI3/MM5_d N_XI15/XI3/NET33_XI15/XI3/MM5_g
+ N_VDD_XI15/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI3/MM4 N_XI15/XI3/NET33_XI15/XI3/MM4_d N_XI15/XI3/NET34_XI15/XI3/MM4_g
+ N_VDD_XI15/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI3/MM10 N_XI15/XI3/NET35_XI15/XI3/MM10_d N_XI15/XI3/NET36_XI15/XI3/MM10_g
+ N_VDD_XI15/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI3/MM11 N_XI15/XI3/NET36_XI15/XI3/MM11_d N_XI15/XI3/NET35_XI15/XI3/MM11_g
+ N_VDD_XI15/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI4/MM2 N_XI15/XI4/NET34_XI15/XI4/MM2_d N_XI15/XI4/NET33_XI15/XI4/MM2_g
+ N_VSS_XI15/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI4/MM3 N_XI15/XI4/NET33_XI15/XI4/MM3_d N_WL<26>_XI15/XI4/MM3_g
+ N_BLN<11>_XI15/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI4/MM0 N_XI15/XI4/NET34_XI15/XI4/MM0_d N_WL<26>_XI15/XI4/MM0_g
+ N_BL<11>_XI15/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI4/MM1 N_XI15/XI4/NET33_XI15/XI4/MM1_d N_XI15/XI4/NET34_XI15/XI4/MM1_g
+ N_VSS_XI15/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI4/MM9 N_XI15/XI4/NET36_XI15/XI4/MM9_d N_WL<27>_XI15/XI4/MM9_g
+ N_BL<11>_XI15/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI4/MM6 N_XI15/XI4/NET35_XI15/XI4/MM6_d N_XI15/XI4/NET36_XI15/XI4/MM6_g
+ N_VSS_XI15/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI4/MM7 N_XI15/XI4/NET36_XI15/XI4/MM7_d N_XI15/XI4/NET35_XI15/XI4/MM7_g
+ N_VSS_XI15/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI4/MM8 N_XI15/XI4/NET35_XI15/XI4/MM8_d N_WL<27>_XI15/XI4/MM8_g
+ N_BLN<11>_XI15/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI4/MM5 N_XI15/XI4/NET34_XI15/XI4/MM5_d N_XI15/XI4/NET33_XI15/XI4/MM5_g
+ N_VDD_XI15/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI4/MM4 N_XI15/XI4/NET33_XI15/XI4/MM4_d N_XI15/XI4/NET34_XI15/XI4/MM4_g
+ N_VDD_XI15/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI4/MM10 N_XI15/XI4/NET35_XI15/XI4/MM10_d N_XI15/XI4/NET36_XI15/XI4/MM10_g
+ N_VDD_XI15/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI4/MM11 N_XI15/XI4/NET36_XI15/XI4/MM11_d N_XI15/XI4/NET35_XI15/XI4/MM11_g
+ N_VDD_XI15/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI5/MM2 N_XI15/XI5/NET34_XI15/XI5/MM2_d N_XI15/XI5/NET33_XI15/XI5/MM2_g
+ N_VSS_XI15/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI5/MM3 N_XI15/XI5/NET33_XI15/XI5/MM3_d N_WL<26>_XI15/XI5/MM3_g
+ N_BLN<10>_XI15/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI5/MM0 N_XI15/XI5/NET34_XI15/XI5/MM0_d N_WL<26>_XI15/XI5/MM0_g
+ N_BL<10>_XI15/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI5/MM1 N_XI15/XI5/NET33_XI15/XI5/MM1_d N_XI15/XI5/NET34_XI15/XI5/MM1_g
+ N_VSS_XI15/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI5/MM9 N_XI15/XI5/NET36_XI15/XI5/MM9_d N_WL<27>_XI15/XI5/MM9_g
+ N_BL<10>_XI15/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI5/MM6 N_XI15/XI5/NET35_XI15/XI5/MM6_d N_XI15/XI5/NET36_XI15/XI5/MM6_g
+ N_VSS_XI15/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI5/MM7 N_XI15/XI5/NET36_XI15/XI5/MM7_d N_XI15/XI5/NET35_XI15/XI5/MM7_g
+ N_VSS_XI15/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI5/MM8 N_XI15/XI5/NET35_XI15/XI5/MM8_d N_WL<27>_XI15/XI5/MM8_g
+ N_BLN<10>_XI15/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI5/MM5 N_XI15/XI5/NET34_XI15/XI5/MM5_d N_XI15/XI5/NET33_XI15/XI5/MM5_g
+ N_VDD_XI15/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI5/MM4 N_XI15/XI5/NET33_XI15/XI5/MM4_d N_XI15/XI5/NET34_XI15/XI5/MM4_g
+ N_VDD_XI15/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI5/MM10 N_XI15/XI5/NET35_XI15/XI5/MM10_d N_XI15/XI5/NET36_XI15/XI5/MM10_g
+ N_VDD_XI15/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI5/MM11 N_XI15/XI5/NET36_XI15/XI5/MM11_d N_XI15/XI5/NET35_XI15/XI5/MM11_g
+ N_VDD_XI15/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI6/MM2 N_XI15/XI6/NET34_XI15/XI6/MM2_d N_XI15/XI6/NET33_XI15/XI6/MM2_g
+ N_VSS_XI15/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM3 N_XI15/XI6/NET33_XI15/XI6/MM3_d N_WL<26>_XI15/XI6/MM3_g
+ N_BLN<9>_XI15/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM0 N_XI15/XI6/NET34_XI15/XI6/MM0_d N_WL<26>_XI15/XI6/MM0_g
+ N_BL<9>_XI15/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM1 N_XI15/XI6/NET33_XI15/XI6/MM1_d N_XI15/XI6/NET34_XI15/XI6/MM1_g
+ N_VSS_XI15/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM9 N_XI15/XI6/NET36_XI15/XI6/MM9_d N_WL<27>_XI15/XI6/MM9_g
+ N_BL<9>_XI15/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM6 N_XI15/XI6/NET35_XI15/XI6/MM6_d N_XI15/XI6/NET36_XI15/XI6/MM6_g
+ N_VSS_XI15/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM7 N_XI15/XI6/NET36_XI15/XI6/MM7_d N_XI15/XI6/NET35_XI15/XI6/MM7_g
+ N_VSS_XI15/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM8 N_XI15/XI6/NET35_XI15/XI6/MM8_d N_WL<27>_XI15/XI6/MM8_g
+ N_BLN<9>_XI15/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI6/MM5 N_XI15/XI6/NET34_XI15/XI6/MM5_d N_XI15/XI6/NET33_XI15/XI6/MM5_g
+ N_VDD_XI15/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI6/MM4 N_XI15/XI6/NET33_XI15/XI6/MM4_d N_XI15/XI6/NET34_XI15/XI6/MM4_g
+ N_VDD_XI15/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI6/MM10 N_XI15/XI6/NET35_XI15/XI6/MM10_d N_XI15/XI6/NET36_XI15/XI6/MM10_g
+ N_VDD_XI15/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI6/MM11 N_XI15/XI6/NET36_XI15/XI6/MM11_d N_XI15/XI6/NET35_XI15/XI6/MM11_g
+ N_VDD_XI15/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI7/MM2 N_XI15/XI7/NET34_XI15/XI7/MM2_d N_XI15/XI7/NET33_XI15/XI7/MM2_g
+ N_VSS_XI15/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM3 N_XI15/XI7/NET33_XI15/XI7/MM3_d N_WL<26>_XI15/XI7/MM3_g
+ N_BLN<8>_XI15/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM0 N_XI15/XI7/NET34_XI15/XI7/MM0_d N_WL<26>_XI15/XI7/MM0_g
+ N_BL<8>_XI15/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM1 N_XI15/XI7/NET33_XI15/XI7/MM1_d N_XI15/XI7/NET34_XI15/XI7/MM1_g
+ N_VSS_XI15/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM9 N_XI15/XI7/NET36_XI15/XI7/MM9_d N_WL<27>_XI15/XI7/MM9_g
+ N_BL<8>_XI15/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM6 N_XI15/XI7/NET35_XI15/XI7/MM6_d N_XI15/XI7/NET36_XI15/XI7/MM6_g
+ N_VSS_XI15/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM7 N_XI15/XI7/NET36_XI15/XI7/MM7_d N_XI15/XI7/NET35_XI15/XI7/MM7_g
+ N_VSS_XI15/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM8 N_XI15/XI7/NET35_XI15/XI7/MM8_d N_WL<27>_XI15/XI7/MM8_g
+ N_BLN<8>_XI15/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI7/MM5 N_XI15/XI7/NET34_XI15/XI7/MM5_d N_XI15/XI7/NET33_XI15/XI7/MM5_g
+ N_VDD_XI15/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI7/MM4 N_XI15/XI7/NET33_XI15/XI7/MM4_d N_XI15/XI7/NET34_XI15/XI7/MM4_g
+ N_VDD_XI15/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI7/MM10 N_XI15/XI7/NET35_XI15/XI7/MM10_d N_XI15/XI7/NET36_XI15/XI7/MM10_g
+ N_VDD_XI15/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI7/MM11 N_XI15/XI7/NET36_XI15/XI7/MM11_d N_XI15/XI7/NET35_XI15/XI7/MM11_g
+ N_VDD_XI15/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI8/MM2 N_XI15/XI8/NET34_XI15/XI8/MM2_d N_XI15/XI8/NET33_XI15/XI8/MM2_g
+ N_VSS_XI15/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM3 N_XI15/XI8/NET33_XI15/XI8/MM3_d N_WL<26>_XI15/XI8/MM3_g
+ N_BLN<7>_XI15/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM0 N_XI15/XI8/NET34_XI15/XI8/MM0_d N_WL<26>_XI15/XI8/MM0_g
+ N_BL<7>_XI15/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM1 N_XI15/XI8/NET33_XI15/XI8/MM1_d N_XI15/XI8/NET34_XI15/XI8/MM1_g
+ N_VSS_XI15/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM9 N_XI15/XI8/NET36_XI15/XI8/MM9_d N_WL<27>_XI15/XI8/MM9_g
+ N_BL<7>_XI15/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM6 N_XI15/XI8/NET35_XI15/XI8/MM6_d N_XI15/XI8/NET36_XI15/XI8/MM6_g
+ N_VSS_XI15/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM7 N_XI15/XI8/NET36_XI15/XI8/MM7_d N_XI15/XI8/NET35_XI15/XI8/MM7_g
+ N_VSS_XI15/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM8 N_XI15/XI8/NET35_XI15/XI8/MM8_d N_WL<27>_XI15/XI8/MM8_g
+ N_BLN<7>_XI15/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI8/MM5 N_XI15/XI8/NET34_XI15/XI8/MM5_d N_XI15/XI8/NET33_XI15/XI8/MM5_g
+ N_VDD_XI15/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI8/MM4 N_XI15/XI8/NET33_XI15/XI8/MM4_d N_XI15/XI8/NET34_XI15/XI8/MM4_g
+ N_VDD_XI15/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI8/MM10 N_XI15/XI8/NET35_XI15/XI8/MM10_d N_XI15/XI8/NET36_XI15/XI8/MM10_g
+ N_VDD_XI15/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI8/MM11 N_XI15/XI8/NET36_XI15/XI8/MM11_d N_XI15/XI8/NET35_XI15/XI8/MM11_g
+ N_VDD_XI15/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI9/MM2 N_XI15/XI9/NET34_XI15/XI9/MM2_d N_XI15/XI9/NET33_XI15/XI9/MM2_g
+ N_VSS_XI15/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM3 N_XI15/XI9/NET33_XI15/XI9/MM3_d N_WL<26>_XI15/XI9/MM3_g
+ N_BLN<6>_XI15/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM0 N_XI15/XI9/NET34_XI15/XI9/MM0_d N_WL<26>_XI15/XI9/MM0_g
+ N_BL<6>_XI15/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM1 N_XI15/XI9/NET33_XI15/XI9/MM1_d N_XI15/XI9/NET34_XI15/XI9/MM1_g
+ N_VSS_XI15/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM9 N_XI15/XI9/NET36_XI15/XI9/MM9_d N_WL<27>_XI15/XI9/MM9_g
+ N_BL<6>_XI15/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM6 N_XI15/XI9/NET35_XI15/XI9/MM6_d N_XI15/XI9/NET36_XI15/XI9/MM6_g
+ N_VSS_XI15/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM7 N_XI15/XI9/NET36_XI15/XI9/MM7_d N_XI15/XI9/NET35_XI15/XI9/MM7_g
+ N_VSS_XI15/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM8 N_XI15/XI9/NET35_XI15/XI9/MM8_d N_WL<27>_XI15/XI9/MM8_g
+ N_BLN<6>_XI15/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI9/MM5 N_XI15/XI9/NET34_XI15/XI9/MM5_d N_XI15/XI9/NET33_XI15/XI9/MM5_g
+ N_VDD_XI15/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI9/MM4 N_XI15/XI9/NET33_XI15/XI9/MM4_d N_XI15/XI9/NET34_XI15/XI9/MM4_g
+ N_VDD_XI15/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI9/MM10 N_XI15/XI9/NET35_XI15/XI9/MM10_d N_XI15/XI9/NET36_XI15/XI9/MM10_g
+ N_VDD_XI15/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI9/MM11 N_XI15/XI9/NET36_XI15/XI9/MM11_d N_XI15/XI9/NET35_XI15/XI9/MM11_g
+ N_VDD_XI15/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI10/MM2 N_XI15/XI10/NET34_XI15/XI10/MM2_d
+ N_XI15/XI10/NET33_XI15/XI10/MM2_g N_VSS_XI15/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI10/MM3 N_XI15/XI10/NET33_XI15/XI10/MM3_d N_WL<26>_XI15/XI10/MM3_g
+ N_BLN<5>_XI15/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI10/MM0 N_XI15/XI10/NET34_XI15/XI10/MM0_d N_WL<26>_XI15/XI10/MM0_g
+ N_BL<5>_XI15/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI10/MM1 N_XI15/XI10/NET33_XI15/XI10/MM1_d
+ N_XI15/XI10/NET34_XI15/XI10/MM1_g N_VSS_XI15/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI10/MM9 N_XI15/XI10/NET36_XI15/XI10/MM9_d N_WL<27>_XI15/XI10/MM9_g
+ N_BL<5>_XI15/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI10/MM6 N_XI15/XI10/NET35_XI15/XI10/MM6_d
+ N_XI15/XI10/NET36_XI15/XI10/MM6_g N_VSS_XI15/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI10/MM7 N_XI15/XI10/NET36_XI15/XI10/MM7_d
+ N_XI15/XI10/NET35_XI15/XI10/MM7_g N_VSS_XI15/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI10/MM8 N_XI15/XI10/NET35_XI15/XI10/MM8_d N_WL<27>_XI15/XI10/MM8_g
+ N_BLN<5>_XI15/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI10/MM5 N_XI15/XI10/NET34_XI15/XI10/MM5_d
+ N_XI15/XI10/NET33_XI15/XI10/MM5_g N_VDD_XI15/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI10/MM4 N_XI15/XI10/NET33_XI15/XI10/MM4_d
+ N_XI15/XI10/NET34_XI15/XI10/MM4_g N_VDD_XI15/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI10/MM10 N_XI15/XI10/NET35_XI15/XI10/MM10_d
+ N_XI15/XI10/NET36_XI15/XI10/MM10_g N_VDD_XI15/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI10/MM11 N_XI15/XI10/NET36_XI15/XI10/MM11_d
+ N_XI15/XI10/NET35_XI15/XI10/MM11_g N_VDD_XI15/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI11/MM2 N_XI15/XI11/NET34_XI15/XI11/MM2_d
+ N_XI15/XI11/NET33_XI15/XI11/MM2_g N_VSS_XI15/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI11/MM3 N_XI15/XI11/NET33_XI15/XI11/MM3_d N_WL<26>_XI15/XI11/MM3_g
+ N_BLN<4>_XI15/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI11/MM0 N_XI15/XI11/NET34_XI15/XI11/MM0_d N_WL<26>_XI15/XI11/MM0_g
+ N_BL<4>_XI15/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI11/MM1 N_XI15/XI11/NET33_XI15/XI11/MM1_d
+ N_XI15/XI11/NET34_XI15/XI11/MM1_g N_VSS_XI15/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI11/MM9 N_XI15/XI11/NET36_XI15/XI11/MM9_d N_WL<27>_XI15/XI11/MM9_g
+ N_BL<4>_XI15/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI11/MM6 N_XI15/XI11/NET35_XI15/XI11/MM6_d
+ N_XI15/XI11/NET36_XI15/XI11/MM6_g N_VSS_XI15/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI11/MM7 N_XI15/XI11/NET36_XI15/XI11/MM7_d
+ N_XI15/XI11/NET35_XI15/XI11/MM7_g N_VSS_XI15/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI11/MM8 N_XI15/XI11/NET35_XI15/XI11/MM8_d N_WL<27>_XI15/XI11/MM8_g
+ N_BLN<4>_XI15/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI11/MM5 N_XI15/XI11/NET34_XI15/XI11/MM5_d
+ N_XI15/XI11/NET33_XI15/XI11/MM5_g N_VDD_XI15/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI11/MM4 N_XI15/XI11/NET33_XI15/XI11/MM4_d
+ N_XI15/XI11/NET34_XI15/XI11/MM4_g N_VDD_XI15/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI11/MM10 N_XI15/XI11/NET35_XI15/XI11/MM10_d
+ N_XI15/XI11/NET36_XI15/XI11/MM10_g N_VDD_XI15/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI11/MM11 N_XI15/XI11/NET36_XI15/XI11/MM11_d
+ N_XI15/XI11/NET35_XI15/XI11/MM11_g N_VDD_XI15/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI12/MM2 N_XI15/XI12/NET34_XI15/XI12/MM2_d
+ N_XI15/XI12/NET33_XI15/XI12/MM2_g N_VSS_XI15/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI12/MM3 N_XI15/XI12/NET33_XI15/XI12/MM3_d N_WL<26>_XI15/XI12/MM3_g
+ N_BLN<3>_XI15/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI12/MM0 N_XI15/XI12/NET34_XI15/XI12/MM0_d N_WL<26>_XI15/XI12/MM0_g
+ N_BL<3>_XI15/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI12/MM1 N_XI15/XI12/NET33_XI15/XI12/MM1_d
+ N_XI15/XI12/NET34_XI15/XI12/MM1_g N_VSS_XI15/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI12/MM9 N_XI15/XI12/NET36_XI15/XI12/MM9_d N_WL<27>_XI15/XI12/MM9_g
+ N_BL<3>_XI15/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI12/MM6 N_XI15/XI12/NET35_XI15/XI12/MM6_d
+ N_XI15/XI12/NET36_XI15/XI12/MM6_g N_VSS_XI15/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI12/MM7 N_XI15/XI12/NET36_XI15/XI12/MM7_d
+ N_XI15/XI12/NET35_XI15/XI12/MM7_g N_VSS_XI15/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI12/MM8 N_XI15/XI12/NET35_XI15/XI12/MM8_d N_WL<27>_XI15/XI12/MM8_g
+ N_BLN<3>_XI15/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI12/MM5 N_XI15/XI12/NET34_XI15/XI12/MM5_d
+ N_XI15/XI12/NET33_XI15/XI12/MM5_g N_VDD_XI15/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI12/MM4 N_XI15/XI12/NET33_XI15/XI12/MM4_d
+ N_XI15/XI12/NET34_XI15/XI12/MM4_g N_VDD_XI15/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI12/MM10 N_XI15/XI12/NET35_XI15/XI12/MM10_d
+ N_XI15/XI12/NET36_XI15/XI12/MM10_g N_VDD_XI15/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI12/MM11 N_XI15/XI12/NET36_XI15/XI12/MM11_d
+ N_XI15/XI12/NET35_XI15/XI12/MM11_g N_VDD_XI15/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI13/MM2 N_XI15/XI13/NET34_XI15/XI13/MM2_d
+ N_XI15/XI13/NET33_XI15/XI13/MM2_g N_VSS_XI15/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI13/MM3 N_XI15/XI13/NET33_XI15/XI13/MM3_d N_WL<26>_XI15/XI13/MM3_g
+ N_BLN<2>_XI15/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI13/MM0 N_XI15/XI13/NET34_XI15/XI13/MM0_d N_WL<26>_XI15/XI13/MM0_g
+ N_BL<2>_XI15/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI13/MM1 N_XI15/XI13/NET33_XI15/XI13/MM1_d
+ N_XI15/XI13/NET34_XI15/XI13/MM1_g N_VSS_XI15/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI13/MM9 N_XI15/XI13/NET36_XI15/XI13/MM9_d N_WL<27>_XI15/XI13/MM9_g
+ N_BL<2>_XI15/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI13/MM6 N_XI15/XI13/NET35_XI15/XI13/MM6_d
+ N_XI15/XI13/NET36_XI15/XI13/MM6_g N_VSS_XI15/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI13/MM7 N_XI15/XI13/NET36_XI15/XI13/MM7_d
+ N_XI15/XI13/NET35_XI15/XI13/MM7_g N_VSS_XI15/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI13/MM8 N_XI15/XI13/NET35_XI15/XI13/MM8_d N_WL<27>_XI15/XI13/MM8_g
+ N_BLN<2>_XI15/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI13/MM5 N_XI15/XI13/NET34_XI15/XI13/MM5_d
+ N_XI15/XI13/NET33_XI15/XI13/MM5_g N_VDD_XI15/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI13/MM4 N_XI15/XI13/NET33_XI15/XI13/MM4_d
+ N_XI15/XI13/NET34_XI15/XI13/MM4_g N_VDD_XI15/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI13/MM10 N_XI15/XI13/NET35_XI15/XI13/MM10_d
+ N_XI15/XI13/NET36_XI15/XI13/MM10_g N_VDD_XI15/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI13/MM11 N_XI15/XI13/NET36_XI15/XI13/MM11_d
+ N_XI15/XI13/NET35_XI15/XI13/MM11_g N_VDD_XI15/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI14/MM2 N_XI15/XI14/NET34_XI15/XI14/MM2_d
+ N_XI15/XI14/NET33_XI15/XI14/MM2_g N_VSS_XI15/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI14/MM3 N_XI15/XI14/NET33_XI15/XI14/MM3_d N_WL<26>_XI15/XI14/MM3_g
+ N_BLN<1>_XI15/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI14/MM0 N_XI15/XI14/NET34_XI15/XI14/MM0_d N_WL<26>_XI15/XI14/MM0_g
+ N_BL<1>_XI15/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI14/MM1 N_XI15/XI14/NET33_XI15/XI14/MM1_d
+ N_XI15/XI14/NET34_XI15/XI14/MM1_g N_VSS_XI15/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI14/MM9 N_XI15/XI14/NET36_XI15/XI14/MM9_d N_WL<27>_XI15/XI14/MM9_g
+ N_BL<1>_XI15/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI14/MM6 N_XI15/XI14/NET35_XI15/XI14/MM6_d
+ N_XI15/XI14/NET36_XI15/XI14/MM6_g N_VSS_XI15/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI14/MM7 N_XI15/XI14/NET36_XI15/XI14/MM7_d
+ N_XI15/XI14/NET35_XI15/XI14/MM7_g N_VSS_XI15/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI14/MM8 N_XI15/XI14/NET35_XI15/XI14/MM8_d N_WL<27>_XI15/XI14/MM8_g
+ N_BLN<1>_XI15/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI14/MM5 N_XI15/XI14/NET34_XI15/XI14/MM5_d
+ N_XI15/XI14/NET33_XI15/XI14/MM5_g N_VDD_XI15/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI14/MM4 N_XI15/XI14/NET33_XI15/XI14/MM4_d
+ N_XI15/XI14/NET34_XI15/XI14/MM4_g N_VDD_XI15/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI14/MM10 N_XI15/XI14/NET35_XI15/XI14/MM10_d
+ N_XI15/XI14/NET36_XI15/XI14/MM10_g N_VDD_XI15/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI14/MM11 N_XI15/XI14/NET36_XI15/XI14/MM11_d
+ N_XI15/XI14/NET35_XI15/XI14/MM11_g N_VDD_XI15/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI15/MM2 N_XI15/XI15/NET34_XI15/XI15/MM2_d
+ N_XI15/XI15/NET33_XI15/XI15/MM2_g N_VSS_XI15/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI15/MM3 N_XI15/XI15/NET33_XI15/XI15/MM3_d N_WL<26>_XI15/XI15/MM3_g
+ N_BLN<0>_XI15/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI15/MM0 N_XI15/XI15/NET34_XI15/XI15/MM0_d N_WL<26>_XI15/XI15/MM0_g
+ N_BL<0>_XI15/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI15/MM1 N_XI15/XI15/NET33_XI15/XI15/MM1_d
+ N_XI15/XI15/NET34_XI15/XI15/MM1_g N_VSS_XI15/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI15/MM9 N_XI15/XI15/NET36_XI15/XI15/MM9_d N_WL<27>_XI15/XI15/MM9_g
+ N_BL<0>_XI15/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI15/MM6 N_XI15/XI15/NET35_XI15/XI15/MM6_d
+ N_XI15/XI15/NET36_XI15/XI15/MM6_g N_VSS_XI15/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI15/MM7 N_XI15/XI15/NET36_XI15/XI15/MM7_d
+ N_XI15/XI15/NET35_XI15/XI15/MM7_g N_VSS_XI15/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/XI15/MM8 N_XI15/XI15/NET35_XI15/XI15/MM8_d N_WL<27>_XI15/XI15/MM8_g
+ N_BLN<0>_XI15/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI15/XI15/MM5 N_XI15/XI15/NET34_XI15/XI15/MM5_d
+ N_XI15/XI15/NET33_XI15/XI15/MM5_g N_VDD_XI15/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI15/MM4 N_XI15/XI15/NET33_XI15/XI15/MM4_d
+ N_XI15/XI15/NET34_XI15/XI15/MM4_g N_VDD_XI15/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI15/MM10 N_XI15/XI15/NET35_XI15/XI15/MM10_d
+ N_XI15/XI15/NET36_XI15/XI15/MM10_g N_VDD_XI15/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/XI15/MM11 N_XI15/XI15/NET36_XI15/XI15/MM11_d
+ N_XI15/XI15/NET35_XI15/XI15/MM11_g N_VDD_XI15/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI0/MM2 N_XI16/XI0/NET34_XI16/XI0/MM2_d N_XI16/XI0/NET33_XI16/XI0/MM2_g
+ N_VSS_XI16/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI0/MM3 N_XI16/XI0/NET33_XI16/XI0/MM3_d N_WL<28>_XI16/XI0/MM3_g
+ N_BLN<15>_XI16/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI0/MM0 N_XI16/XI0/NET34_XI16/XI0/MM0_d N_WL<28>_XI16/XI0/MM0_g
+ N_BL<15>_XI16/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI0/MM1 N_XI16/XI0/NET33_XI16/XI0/MM1_d N_XI16/XI0/NET34_XI16/XI0/MM1_g
+ N_VSS_XI16/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI0/MM9 N_XI16/XI0/NET36_XI16/XI0/MM9_d N_WL<29>_XI16/XI0/MM9_g
+ N_BL<15>_XI16/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI0/MM6 N_XI16/XI0/NET35_XI16/XI0/MM6_d N_XI16/XI0/NET36_XI16/XI0/MM6_g
+ N_VSS_XI16/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI0/MM7 N_XI16/XI0/NET36_XI16/XI0/MM7_d N_XI16/XI0/NET35_XI16/XI0/MM7_g
+ N_VSS_XI16/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI0/MM8 N_XI16/XI0/NET35_XI16/XI0/MM8_d N_WL<29>_XI16/XI0/MM8_g
+ N_BLN<15>_XI16/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI0/MM5 N_XI16/XI0/NET34_XI16/XI0/MM5_d N_XI16/XI0/NET33_XI16/XI0/MM5_g
+ N_VDD_XI16/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI0/MM4 N_XI16/XI0/NET33_XI16/XI0/MM4_d N_XI16/XI0/NET34_XI16/XI0/MM4_g
+ N_VDD_XI16/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI0/MM10 N_XI16/XI0/NET35_XI16/XI0/MM10_d N_XI16/XI0/NET36_XI16/XI0/MM10_g
+ N_VDD_XI16/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI0/MM11 N_XI16/XI0/NET36_XI16/XI0/MM11_d N_XI16/XI0/NET35_XI16/XI0/MM11_g
+ N_VDD_XI16/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI1/MM2 N_XI16/XI1/NET34_XI16/XI1/MM2_d N_XI16/XI1/NET33_XI16/XI1/MM2_g
+ N_VSS_XI16/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI1/MM3 N_XI16/XI1/NET33_XI16/XI1/MM3_d N_WL<28>_XI16/XI1/MM3_g
+ N_BLN<14>_XI16/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI1/MM0 N_XI16/XI1/NET34_XI16/XI1/MM0_d N_WL<28>_XI16/XI1/MM0_g
+ N_BL<14>_XI16/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI1/MM1 N_XI16/XI1/NET33_XI16/XI1/MM1_d N_XI16/XI1/NET34_XI16/XI1/MM1_g
+ N_VSS_XI16/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI1/MM9 N_XI16/XI1/NET36_XI16/XI1/MM9_d N_WL<29>_XI16/XI1/MM9_g
+ N_BL<14>_XI16/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI1/MM6 N_XI16/XI1/NET35_XI16/XI1/MM6_d N_XI16/XI1/NET36_XI16/XI1/MM6_g
+ N_VSS_XI16/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI1/MM7 N_XI16/XI1/NET36_XI16/XI1/MM7_d N_XI16/XI1/NET35_XI16/XI1/MM7_g
+ N_VSS_XI16/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI1/MM8 N_XI16/XI1/NET35_XI16/XI1/MM8_d N_WL<29>_XI16/XI1/MM8_g
+ N_BLN<14>_XI16/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI1/MM5 N_XI16/XI1/NET34_XI16/XI1/MM5_d N_XI16/XI1/NET33_XI16/XI1/MM5_g
+ N_VDD_XI16/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI1/MM4 N_XI16/XI1/NET33_XI16/XI1/MM4_d N_XI16/XI1/NET34_XI16/XI1/MM4_g
+ N_VDD_XI16/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI1/MM10 N_XI16/XI1/NET35_XI16/XI1/MM10_d N_XI16/XI1/NET36_XI16/XI1/MM10_g
+ N_VDD_XI16/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI1/MM11 N_XI16/XI1/NET36_XI16/XI1/MM11_d N_XI16/XI1/NET35_XI16/XI1/MM11_g
+ N_VDD_XI16/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI2/MM2 N_XI16/XI2/NET34_XI16/XI2/MM2_d N_XI16/XI2/NET33_XI16/XI2/MM2_g
+ N_VSS_XI16/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI2/MM3 N_XI16/XI2/NET33_XI16/XI2/MM3_d N_WL<28>_XI16/XI2/MM3_g
+ N_BLN<13>_XI16/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI2/MM0 N_XI16/XI2/NET34_XI16/XI2/MM0_d N_WL<28>_XI16/XI2/MM0_g
+ N_BL<13>_XI16/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI2/MM1 N_XI16/XI2/NET33_XI16/XI2/MM1_d N_XI16/XI2/NET34_XI16/XI2/MM1_g
+ N_VSS_XI16/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI2/MM9 N_XI16/XI2/NET36_XI16/XI2/MM9_d N_WL<29>_XI16/XI2/MM9_g
+ N_BL<13>_XI16/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI2/MM6 N_XI16/XI2/NET35_XI16/XI2/MM6_d N_XI16/XI2/NET36_XI16/XI2/MM6_g
+ N_VSS_XI16/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI2/MM7 N_XI16/XI2/NET36_XI16/XI2/MM7_d N_XI16/XI2/NET35_XI16/XI2/MM7_g
+ N_VSS_XI16/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI2/MM8 N_XI16/XI2/NET35_XI16/XI2/MM8_d N_WL<29>_XI16/XI2/MM8_g
+ N_BLN<13>_XI16/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI2/MM5 N_XI16/XI2/NET34_XI16/XI2/MM5_d N_XI16/XI2/NET33_XI16/XI2/MM5_g
+ N_VDD_XI16/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI2/MM4 N_XI16/XI2/NET33_XI16/XI2/MM4_d N_XI16/XI2/NET34_XI16/XI2/MM4_g
+ N_VDD_XI16/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI2/MM10 N_XI16/XI2/NET35_XI16/XI2/MM10_d N_XI16/XI2/NET36_XI16/XI2/MM10_g
+ N_VDD_XI16/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI2/MM11 N_XI16/XI2/NET36_XI16/XI2/MM11_d N_XI16/XI2/NET35_XI16/XI2/MM11_g
+ N_VDD_XI16/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI3/MM2 N_XI16/XI3/NET34_XI16/XI3/MM2_d N_XI16/XI3/NET33_XI16/XI3/MM2_g
+ N_VSS_XI16/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI3/MM3 N_XI16/XI3/NET33_XI16/XI3/MM3_d N_WL<28>_XI16/XI3/MM3_g
+ N_BLN<12>_XI16/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI3/MM0 N_XI16/XI3/NET34_XI16/XI3/MM0_d N_WL<28>_XI16/XI3/MM0_g
+ N_BL<12>_XI16/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI3/MM1 N_XI16/XI3/NET33_XI16/XI3/MM1_d N_XI16/XI3/NET34_XI16/XI3/MM1_g
+ N_VSS_XI16/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI3/MM9 N_XI16/XI3/NET36_XI16/XI3/MM9_d N_WL<29>_XI16/XI3/MM9_g
+ N_BL<12>_XI16/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI3/MM6 N_XI16/XI3/NET35_XI16/XI3/MM6_d N_XI16/XI3/NET36_XI16/XI3/MM6_g
+ N_VSS_XI16/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI3/MM7 N_XI16/XI3/NET36_XI16/XI3/MM7_d N_XI16/XI3/NET35_XI16/XI3/MM7_g
+ N_VSS_XI16/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI3/MM8 N_XI16/XI3/NET35_XI16/XI3/MM8_d N_WL<29>_XI16/XI3/MM8_g
+ N_BLN<12>_XI16/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI3/MM5 N_XI16/XI3/NET34_XI16/XI3/MM5_d N_XI16/XI3/NET33_XI16/XI3/MM5_g
+ N_VDD_XI16/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI3/MM4 N_XI16/XI3/NET33_XI16/XI3/MM4_d N_XI16/XI3/NET34_XI16/XI3/MM4_g
+ N_VDD_XI16/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI3/MM10 N_XI16/XI3/NET35_XI16/XI3/MM10_d N_XI16/XI3/NET36_XI16/XI3/MM10_g
+ N_VDD_XI16/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI3/MM11 N_XI16/XI3/NET36_XI16/XI3/MM11_d N_XI16/XI3/NET35_XI16/XI3/MM11_g
+ N_VDD_XI16/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI4/MM2 N_XI16/XI4/NET34_XI16/XI4/MM2_d N_XI16/XI4/NET33_XI16/XI4/MM2_g
+ N_VSS_XI16/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI4/MM3 N_XI16/XI4/NET33_XI16/XI4/MM3_d N_WL<28>_XI16/XI4/MM3_g
+ N_BLN<11>_XI16/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI4/MM0 N_XI16/XI4/NET34_XI16/XI4/MM0_d N_WL<28>_XI16/XI4/MM0_g
+ N_BL<11>_XI16/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI4/MM1 N_XI16/XI4/NET33_XI16/XI4/MM1_d N_XI16/XI4/NET34_XI16/XI4/MM1_g
+ N_VSS_XI16/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI4/MM9 N_XI16/XI4/NET36_XI16/XI4/MM9_d N_WL<29>_XI16/XI4/MM9_g
+ N_BL<11>_XI16/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI4/MM6 N_XI16/XI4/NET35_XI16/XI4/MM6_d N_XI16/XI4/NET36_XI16/XI4/MM6_g
+ N_VSS_XI16/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI4/MM7 N_XI16/XI4/NET36_XI16/XI4/MM7_d N_XI16/XI4/NET35_XI16/XI4/MM7_g
+ N_VSS_XI16/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI4/MM8 N_XI16/XI4/NET35_XI16/XI4/MM8_d N_WL<29>_XI16/XI4/MM8_g
+ N_BLN<11>_XI16/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI4/MM5 N_XI16/XI4/NET34_XI16/XI4/MM5_d N_XI16/XI4/NET33_XI16/XI4/MM5_g
+ N_VDD_XI16/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI4/MM4 N_XI16/XI4/NET33_XI16/XI4/MM4_d N_XI16/XI4/NET34_XI16/XI4/MM4_g
+ N_VDD_XI16/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI4/MM10 N_XI16/XI4/NET35_XI16/XI4/MM10_d N_XI16/XI4/NET36_XI16/XI4/MM10_g
+ N_VDD_XI16/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI4/MM11 N_XI16/XI4/NET36_XI16/XI4/MM11_d N_XI16/XI4/NET35_XI16/XI4/MM11_g
+ N_VDD_XI16/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI5/MM2 N_XI16/XI5/NET34_XI16/XI5/MM2_d N_XI16/XI5/NET33_XI16/XI5/MM2_g
+ N_VSS_XI16/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI5/MM3 N_XI16/XI5/NET33_XI16/XI5/MM3_d N_WL<28>_XI16/XI5/MM3_g
+ N_BLN<10>_XI16/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI5/MM0 N_XI16/XI5/NET34_XI16/XI5/MM0_d N_WL<28>_XI16/XI5/MM0_g
+ N_BL<10>_XI16/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI5/MM1 N_XI16/XI5/NET33_XI16/XI5/MM1_d N_XI16/XI5/NET34_XI16/XI5/MM1_g
+ N_VSS_XI16/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI5/MM9 N_XI16/XI5/NET36_XI16/XI5/MM9_d N_WL<29>_XI16/XI5/MM9_g
+ N_BL<10>_XI16/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI5/MM6 N_XI16/XI5/NET35_XI16/XI5/MM6_d N_XI16/XI5/NET36_XI16/XI5/MM6_g
+ N_VSS_XI16/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI5/MM7 N_XI16/XI5/NET36_XI16/XI5/MM7_d N_XI16/XI5/NET35_XI16/XI5/MM7_g
+ N_VSS_XI16/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI5/MM8 N_XI16/XI5/NET35_XI16/XI5/MM8_d N_WL<29>_XI16/XI5/MM8_g
+ N_BLN<10>_XI16/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI5/MM5 N_XI16/XI5/NET34_XI16/XI5/MM5_d N_XI16/XI5/NET33_XI16/XI5/MM5_g
+ N_VDD_XI16/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI5/MM4 N_XI16/XI5/NET33_XI16/XI5/MM4_d N_XI16/XI5/NET34_XI16/XI5/MM4_g
+ N_VDD_XI16/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI5/MM10 N_XI16/XI5/NET35_XI16/XI5/MM10_d N_XI16/XI5/NET36_XI16/XI5/MM10_g
+ N_VDD_XI16/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI5/MM11 N_XI16/XI5/NET36_XI16/XI5/MM11_d N_XI16/XI5/NET35_XI16/XI5/MM11_g
+ N_VDD_XI16/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI6/MM2 N_XI16/XI6/NET34_XI16/XI6/MM2_d N_XI16/XI6/NET33_XI16/XI6/MM2_g
+ N_VSS_XI16/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM3 N_XI16/XI6/NET33_XI16/XI6/MM3_d N_WL<28>_XI16/XI6/MM3_g
+ N_BLN<9>_XI16/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM0 N_XI16/XI6/NET34_XI16/XI6/MM0_d N_WL<28>_XI16/XI6/MM0_g
+ N_BL<9>_XI16/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM1 N_XI16/XI6/NET33_XI16/XI6/MM1_d N_XI16/XI6/NET34_XI16/XI6/MM1_g
+ N_VSS_XI16/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM9 N_XI16/XI6/NET36_XI16/XI6/MM9_d N_WL<29>_XI16/XI6/MM9_g
+ N_BL<9>_XI16/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM6 N_XI16/XI6/NET35_XI16/XI6/MM6_d N_XI16/XI6/NET36_XI16/XI6/MM6_g
+ N_VSS_XI16/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM7 N_XI16/XI6/NET36_XI16/XI6/MM7_d N_XI16/XI6/NET35_XI16/XI6/MM7_g
+ N_VSS_XI16/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM8 N_XI16/XI6/NET35_XI16/XI6/MM8_d N_WL<29>_XI16/XI6/MM8_g
+ N_BLN<9>_XI16/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI6/MM5 N_XI16/XI6/NET34_XI16/XI6/MM5_d N_XI16/XI6/NET33_XI16/XI6/MM5_g
+ N_VDD_XI16/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI6/MM4 N_XI16/XI6/NET33_XI16/XI6/MM4_d N_XI16/XI6/NET34_XI16/XI6/MM4_g
+ N_VDD_XI16/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI6/MM10 N_XI16/XI6/NET35_XI16/XI6/MM10_d N_XI16/XI6/NET36_XI16/XI6/MM10_g
+ N_VDD_XI16/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI6/MM11 N_XI16/XI6/NET36_XI16/XI6/MM11_d N_XI16/XI6/NET35_XI16/XI6/MM11_g
+ N_VDD_XI16/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI7/MM2 N_XI16/XI7/NET34_XI16/XI7/MM2_d N_XI16/XI7/NET33_XI16/XI7/MM2_g
+ N_VSS_XI16/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM3 N_XI16/XI7/NET33_XI16/XI7/MM3_d N_WL<28>_XI16/XI7/MM3_g
+ N_BLN<8>_XI16/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM0 N_XI16/XI7/NET34_XI16/XI7/MM0_d N_WL<28>_XI16/XI7/MM0_g
+ N_BL<8>_XI16/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM1 N_XI16/XI7/NET33_XI16/XI7/MM1_d N_XI16/XI7/NET34_XI16/XI7/MM1_g
+ N_VSS_XI16/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM9 N_XI16/XI7/NET36_XI16/XI7/MM9_d N_WL<29>_XI16/XI7/MM9_g
+ N_BL<8>_XI16/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM6 N_XI16/XI7/NET35_XI16/XI7/MM6_d N_XI16/XI7/NET36_XI16/XI7/MM6_g
+ N_VSS_XI16/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM7 N_XI16/XI7/NET36_XI16/XI7/MM7_d N_XI16/XI7/NET35_XI16/XI7/MM7_g
+ N_VSS_XI16/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM8 N_XI16/XI7/NET35_XI16/XI7/MM8_d N_WL<29>_XI16/XI7/MM8_g
+ N_BLN<8>_XI16/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI7/MM5 N_XI16/XI7/NET34_XI16/XI7/MM5_d N_XI16/XI7/NET33_XI16/XI7/MM5_g
+ N_VDD_XI16/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI7/MM4 N_XI16/XI7/NET33_XI16/XI7/MM4_d N_XI16/XI7/NET34_XI16/XI7/MM4_g
+ N_VDD_XI16/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI7/MM10 N_XI16/XI7/NET35_XI16/XI7/MM10_d N_XI16/XI7/NET36_XI16/XI7/MM10_g
+ N_VDD_XI16/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI7/MM11 N_XI16/XI7/NET36_XI16/XI7/MM11_d N_XI16/XI7/NET35_XI16/XI7/MM11_g
+ N_VDD_XI16/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI8/MM2 N_XI16/XI8/NET34_XI16/XI8/MM2_d N_XI16/XI8/NET33_XI16/XI8/MM2_g
+ N_VSS_XI16/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM3 N_XI16/XI8/NET33_XI16/XI8/MM3_d N_WL<28>_XI16/XI8/MM3_g
+ N_BLN<7>_XI16/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM0 N_XI16/XI8/NET34_XI16/XI8/MM0_d N_WL<28>_XI16/XI8/MM0_g
+ N_BL<7>_XI16/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM1 N_XI16/XI8/NET33_XI16/XI8/MM1_d N_XI16/XI8/NET34_XI16/XI8/MM1_g
+ N_VSS_XI16/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM9 N_XI16/XI8/NET36_XI16/XI8/MM9_d N_WL<29>_XI16/XI8/MM9_g
+ N_BL<7>_XI16/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM6 N_XI16/XI8/NET35_XI16/XI8/MM6_d N_XI16/XI8/NET36_XI16/XI8/MM6_g
+ N_VSS_XI16/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM7 N_XI16/XI8/NET36_XI16/XI8/MM7_d N_XI16/XI8/NET35_XI16/XI8/MM7_g
+ N_VSS_XI16/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM8 N_XI16/XI8/NET35_XI16/XI8/MM8_d N_WL<29>_XI16/XI8/MM8_g
+ N_BLN<7>_XI16/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI8/MM5 N_XI16/XI8/NET34_XI16/XI8/MM5_d N_XI16/XI8/NET33_XI16/XI8/MM5_g
+ N_VDD_XI16/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI8/MM4 N_XI16/XI8/NET33_XI16/XI8/MM4_d N_XI16/XI8/NET34_XI16/XI8/MM4_g
+ N_VDD_XI16/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI8/MM10 N_XI16/XI8/NET35_XI16/XI8/MM10_d N_XI16/XI8/NET36_XI16/XI8/MM10_g
+ N_VDD_XI16/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI8/MM11 N_XI16/XI8/NET36_XI16/XI8/MM11_d N_XI16/XI8/NET35_XI16/XI8/MM11_g
+ N_VDD_XI16/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI9/MM2 N_XI16/XI9/NET34_XI16/XI9/MM2_d N_XI16/XI9/NET33_XI16/XI9/MM2_g
+ N_VSS_XI16/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM3 N_XI16/XI9/NET33_XI16/XI9/MM3_d N_WL<28>_XI16/XI9/MM3_g
+ N_BLN<6>_XI16/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM0 N_XI16/XI9/NET34_XI16/XI9/MM0_d N_WL<28>_XI16/XI9/MM0_g
+ N_BL<6>_XI16/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM1 N_XI16/XI9/NET33_XI16/XI9/MM1_d N_XI16/XI9/NET34_XI16/XI9/MM1_g
+ N_VSS_XI16/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM9 N_XI16/XI9/NET36_XI16/XI9/MM9_d N_WL<29>_XI16/XI9/MM9_g
+ N_BL<6>_XI16/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM6 N_XI16/XI9/NET35_XI16/XI9/MM6_d N_XI16/XI9/NET36_XI16/XI9/MM6_g
+ N_VSS_XI16/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM7 N_XI16/XI9/NET36_XI16/XI9/MM7_d N_XI16/XI9/NET35_XI16/XI9/MM7_g
+ N_VSS_XI16/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM8 N_XI16/XI9/NET35_XI16/XI9/MM8_d N_WL<29>_XI16/XI9/MM8_g
+ N_BLN<6>_XI16/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI9/MM5 N_XI16/XI9/NET34_XI16/XI9/MM5_d N_XI16/XI9/NET33_XI16/XI9/MM5_g
+ N_VDD_XI16/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI9/MM4 N_XI16/XI9/NET33_XI16/XI9/MM4_d N_XI16/XI9/NET34_XI16/XI9/MM4_g
+ N_VDD_XI16/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI9/MM10 N_XI16/XI9/NET35_XI16/XI9/MM10_d N_XI16/XI9/NET36_XI16/XI9/MM10_g
+ N_VDD_XI16/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI9/MM11 N_XI16/XI9/NET36_XI16/XI9/MM11_d N_XI16/XI9/NET35_XI16/XI9/MM11_g
+ N_VDD_XI16/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI10/MM2 N_XI16/XI10/NET34_XI16/XI10/MM2_d
+ N_XI16/XI10/NET33_XI16/XI10/MM2_g N_VSS_XI16/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI10/MM3 N_XI16/XI10/NET33_XI16/XI10/MM3_d N_WL<28>_XI16/XI10/MM3_g
+ N_BLN<5>_XI16/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI10/MM0 N_XI16/XI10/NET34_XI16/XI10/MM0_d N_WL<28>_XI16/XI10/MM0_g
+ N_BL<5>_XI16/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI10/MM1 N_XI16/XI10/NET33_XI16/XI10/MM1_d
+ N_XI16/XI10/NET34_XI16/XI10/MM1_g N_VSS_XI16/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI10/MM9 N_XI16/XI10/NET36_XI16/XI10/MM9_d N_WL<29>_XI16/XI10/MM9_g
+ N_BL<5>_XI16/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI10/MM6 N_XI16/XI10/NET35_XI16/XI10/MM6_d
+ N_XI16/XI10/NET36_XI16/XI10/MM6_g N_VSS_XI16/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI10/MM7 N_XI16/XI10/NET36_XI16/XI10/MM7_d
+ N_XI16/XI10/NET35_XI16/XI10/MM7_g N_VSS_XI16/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI10/MM8 N_XI16/XI10/NET35_XI16/XI10/MM8_d N_WL<29>_XI16/XI10/MM8_g
+ N_BLN<5>_XI16/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI10/MM5 N_XI16/XI10/NET34_XI16/XI10/MM5_d
+ N_XI16/XI10/NET33_XI16/XI10/MM5_g N_VDD_XI16/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI10/MM4 N_XI16/XI10/NET33_XI16/XI10/MM4_d
+ N_XI16/XI10/NET34_XI16/XI10/MM4_g N_VDD_XI16/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI10/MM10 N_XI16/XI10/NET35_XI16/XI10/MM10_d
+ N_XI16/XI10/NET36_XI16/XI10/MM10_g N_VDD_XI16/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI10/MM11 N_XI16/XI10/NET36_XI16/XI10/MM11_d
+ N_XI16/XI10/NET35_XI16/XI10/MM11_g N_VDD_XI16/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI11/MM2 N_XI16/XI11/NET34_XI16/XI11/MM2_d
+ N_XI16/XI11/NET33_XI16/XI11/MM2_g N_VSS_XI16/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI11/MM3 N_XI16/XI11/NET33_XI16/XI11/MM3_d N_WL<28>_XI16/XI11/MM3_g
+ N_BLN<4>_XI16/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI11/MM0 N_XI16/XI11/NET34_XI16/XI11/MM0_d N_WL<28>_XI16/XI11/MM0_g
+ N_BL<4>_XI16/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI11/MM1 N_XI16/XI11/NET33_XI16/XI11/MM1_d
+ N_XI16/XI11/NET34_XI16/XI11/MM1_g N_VSS_XI16/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI11/MM9 N_XI16/XI11/NET36_XI16/XI11/MM9_d N_WL<29>_XI16/XI11/MM9_g
+ N_BL<4>_XI16/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI11/MM6 N_XI16/XI11/NET35_XI16/XI11/MM6_d
+ N_XI16/XI11/NET36_XI16/XI11/MM6_g N_VSS_XI16/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI11/MM7 N_XI16/XI11/NET36_XI16/XI11/MM7_d
+ N_XI16/XI11/NET35_XI16/XI11/MM7_g N_VSS_XI16/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI11/MM8 N_XI16/XI11/NET35_XI16/XI11/MM8_d N_WL<29>_XI16/XI11/MM8_g
+ N_BLN<4>_XI16/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI11/MM5 N_XI16/XI11/NET34_XI16/XI11/MM5_d
+ N_XI16/XI11/NET33_XI16/XI11/MM5_g N_VDD_XI16/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI11/MM4 N_XI16/XI11/NET33_XI16/XI11/MM4_d
+ N_XI16/XI11/NET34_XI16/XI11/MM4_g N_VDD_XI16/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI11/MM10 N_XI16/XI11/NET35_XI16/XI11/MM10_d
+ N_XI16/XI11/NET36_XI16/XI11/MM10_g N_VDD_XI16/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI11/MM11 N_XI16/XI11/NET36_XI16/XI11/MM11_d
+ N_XI16/XI11/NET35_XI16/XI11/MM11_g N_VDD_XI16/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI12/MM2 N_XI16/XI12/NET34_XI16/XI12/MM2_d
+ N_XI16/XI12/NET33_XI16/XI12/MM2_g N_VSS_XI16/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI12/MM3 N_XI16/XI12/NET33_XI16/XI12/MM3_d N_WL<28>_XI16/XI12/MM3_g
+ N_BLN<3>_XI16/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI12/MM0 N_XI16/XI12/NET34_XI16/XI12/MM0_d N_WL<28>_XI16/XI12/MM0_g
+ N_BL<3>_XI16/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI12/MM1 N_XI16/XI12/NET33_XI16/XI12/MM1_d
+ N_XI16/XI12/NET34_XI16/XI12/MM1_g N_VSS_XI16/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI12/MM9 N_XI16/XI12/NET36_XI16/XI12/MM9_d N_WL<29>_XI16/XI12/MM9_g
+ N_BL<3>_XI16/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI12/MM6 N_XI16/XI12/NET35_XI16/XI12/MM6_d
+ N_XI16/XI12/NET36_XI16/XI12/MM6_g N_VSS_XI16/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI12/MM7 N_XI16/XI12/NET36_XI16/XI12/MM7_d
+ N_XI16/XI12/NET35_XI16/XI12/MM7_g N_VSS_XI16/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI12/MM8 N_XI16/XI12/NET35_XI16/XI12/MM8_d N_WL<29>_XI16/XI12/MM8_g
+ N_BLN<3>_XI16/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI12/MM5 N_XI16/XI12/NET34_XI16/XI12/MM5_d
+ N_XI16/XI12/NET33_XI16/XI12/MM5_g N_VDD_XI16/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI12/MM4 N_XI16/XI12/NET33_XI16/XI12/MM4_d
+ N_XI16/XI12/NET34_XI16/XI12/MM4_g N_VDD_XI16/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI12/MM10 N_XI16/XI12/NET35_XI16/XI12/MM10_d
+ N_XI16/XI12/NET36_XI16/XI12/MM10_g N_VDD_XI16/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI12/MM11 N_XI16/XI12/NET36_XI16/XI12/MM11_d
+ N_XI16/XI12/NET35_XI16/XI12/MM11_g N_VDD_XI16/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI13/MM2 N_XI16/XI13/NET34_XI16/XI13/MM2_d
+ N_XI16/XI13/NET33_XI16/XI13/MM2_g N_VSS_XI16/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI13/MM3 N_XI16/XI13/NET33_XI16/XI13/MM3_d N_WL<28>_XI16/XI13/MM3_g
+ N_BLN<2>_XI16/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI13/MM0 N_XI16/XI13/NET34_XI16/XI13/MM0_d N_WL<28>_XI16/XI13/MM0_g
+ N_BL<2>_XI16/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI13/MM1 N_XI16/XI13/NET33_XI16/XI13/MM1_d
+ N_XI16/XI13/NET34_XI16/XI13/MM1_g N_VSS_XI16/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI13/MM9 N_XI16/XI13/NET36_XI16/XI13/MM9_d N_WL<29>_XI16/XI13/MM9_g
+ N_BL<2>_XI16/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI13/MM6 N_XI16/XI13/NET35_XI16/XI13/MM6_d
+ N_XI16/XI13/NET36_XI16/XI13/MM6_g N_VSS_XI16/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI13/MM7 N_XI16/XI13/NET36_XI16/XI13/MM7_d
+ N_XI16/XI13/NET35_XI16/XI13/MM7_g N_VSS_XI16/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI13/MM8 N_XI16/XI13/NET35_XI16/XI13/MM8_d N_WL<29>_XI16/XI13/MM8_g
+ N_BLN<2>_XI16/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI13/MM5 N_XI16/XI13/NET34_XI16/XI13/MM5_d
+ N_XI16/XI13/NET33_XI16/XI13/MM5_g N_VDD_XI16/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI13/MM4 N_XI16/XI13/NET33_XI16/XI13/MM4_d
+ N_XI16/XI13/NET34_XI16/XI13/MM4_g N_VDD_XI16/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI13/MM10 N_XI16/XI13/NET35_XI16/XI13/MM10_d
+ N_XI16/XI13/NET36_XI16/XI13/MM10_g N_VDD_XI16/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI13/MM11 N_XI16/XI13/NET36_XI16/XI13/MM11_d
+ N_XI16/XI13/NET35_XI16/XI13/MM11_g N_VDD_XI16/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI14/MM2 N_XI16/XI14/NET34_XI16/XI14/MM2_d
+ N_XI16/XI14/NET33_XI16/XI14/MM2_g N_VSS_XI16/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI14/MM3 N_XI16/XI14/NET33_XI16/XI14/MM3_d N_WL<28>_XI16/XI14/MM3_g
+ N_BLN<1>_XI16/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI14/MM0 N_XI16/XI14/NET34_XI16/XI14/MM0_d N_WL<28>_XI16/XI14/MM0_g
+ N_BL<1>_XI16/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI14/MM1 N_XI16/XI14/NET33_XI16/XI14/MM1_d
+ N_XI16/XI14/NET34_XI16/XI14/MM1_g N_VSS_XI16/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI14/MM9 N_XI16/XI14/NET36_XI16/XI14/MM9_d N_WL<29>_XI16/XI14/MM9_g
+ N_BL<1>_XI16/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI14/MM6 N_XI16/XI14/NET35_XI16/XI14/MM6_d
+ N_XI16/XI14/NET36_XI16/XI14/MM6_g N_VSS_XI16/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI14/MM7 N_XI16/XI14/NET36_XI16/XI14/MM7_d
+ N_XI16/XI14/NET35_XI16/XI14/MM7_g N_VSS_XI16/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI14/MM8 N_XI16/XI14/NET35_XI16/XI14/MM8_d N_WL<29>_XI16/XI14/MM8_g
+ N_BLN<1>_XI16/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI14/MM5 N_XI16/XI14/NET34_XI16/XI14/MM5_d
+ N_XI16/XI14/NET33_XI16/XI14/MM5_g N_VDD_XI16/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI14/MM4 N_XI16/XI14/NET33_XI16/XI14/MM4_d
+ N_XI16/XI14/NET34_XI16/XI14/MM4_g N_VDD_XI16/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI14/MM10 N_XI16/XI14/NET35_XI16/XI14/MM10_d
+ N_XI16/XI14/NET36_XI16/XI14/MM10_g N_VDD_XI16/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI14/MM11 N_XI16/XI14/NET36_XI16/XI14/MM11_d
+ N_XI16/XI14/NET35_XI16/XI14/MM11_g N_VDD_XI16/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI15/MM2 N_XI16/XI15/NET34_XI16/XI15/MM2_d
+ N_XI16/XI15/NET33_XI16/XI15/MM2_g N_VSS_XI16/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI15/MM3 N_XI16/XI15/NET33_XI16/XI15/MM3_d N_WL<28>_XI16/XI15/MM3_g
+ N_BLN<0>_XI16/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI15/MM0 N_XI16/XI15/NET34_XI16/XI15/MM0_d N_WL<28>_XI16/XI15/MM0_g
+ N_BL<0>_XI16/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI15/MM1 N_XI16/XI15/NET33_XI16/XI15/MM1_d
+ N_XI16/XI15/NET34_XI16/XI15/MM1_g N_VSS_XI16/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI15/MM9 N_XI16/XI15/NET36_XI16/XI15/MM9_d N_WL<29>_XI16/XI15/MM9_g
+ N_BL<0>_XI16/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI15/MM6 N_XI16/XI15/NET35_XI16/XI15/MM6_d
+ N_XI16/XI15/NET36_XI16/XI15/MM6_g N_VSS_XI16/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI15/MM7 N_XI16/XI15/NET36_XI16/XI15/MM7_d
+ N_XI16/XI15/NET35_XI16/XI15/MM7_g N_VSS_XI16/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI16/XI15/MM8 N_XI16/XI15/NET35_XI16/XI15/MM8_d N_WL<29>_XI16/XI15/MM8_g
+ N_BLN<0>_XI16/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI16/XI15/MM5 N_XI16/XI15/NET34_XI16/XI15/MM5_d
+ N_XI16/XI15/NET33_XI16/XI15/MM5_g N_VDD_XI16/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI15/MM4 N_XI16/XI15/NET33_XI16/XI15/MM4_d
+ N_XI16/XI15/NET34_XI16/XI15/MM4_g N_VDD_XI16/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI15/MM10 N_XI16/XI15/NET35_XI16/XI15/MM10_d
+ N_XI16/XI15/NET36_XI16/XI15/MM10_g N_VDD_XI16/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI16/XI15/MM11 N_XI16/XI15/NET36_XI16/XI15/MM11_d
+ N_XI16/XI15/NET35_XI16/XI15/MM11_g N_VDD_XI16/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI0/MM2 N_XI17/XI0/NET34_XI17/XI0/MM2_d N_XI17/XI0/NET33_XI17/XI0/MM2_g
+ N_VSS_XI17/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI0/MM3 N_XI17/XI0/NET33_XI17/XI0/MM3_d N_WL<30>_XI17/XI0/MM3_g
+ N_BLN<15>_XI17/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI0/MM0 N_XI17/XI0/NET34_XI17/XI0/MM0_d N_WL<30>_XI17/XI0/MM0_g
+ N_BL<15>_XI17/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI0/MM1 N_XI17/XI0/NET33_XI17/XI0/MM1_d N_XI17/XI0/NET34_XI17/XI0/MM1_g
+ N_VSS_XI17/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI0/MM9 N_XI17/XI0/NET36_XI17/XI0/MM9_d N_WL<31>_XI17/XI0/MM9_g
+ N_BL<15>_XI17/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI0/MM6 N_XI17/XI0/NET35_XI17/XI0/MM6_d N_XI17/XI0/NET36_XI17/XI0/MM6_g
+ N_VSS_XI17/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI0/MM7 N_XI17/XI0/NET36_XI17/XI0/MM7_d N_XI17/XI0/NET35_XI17/XI0/MM7_g
+ N_VSS_XI17/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI0/MM8 N_XI17/XI0/NET35_XI17/XI0/MM8_d N_WL<31>_XI17/XI0/MM8_g
+ N_BLN<15>_XI17/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI0/MM5 N_XI17/XI0/NET34_XI17/XI0/MM5_d N_XI17/XI0/NET33_XI17/XI0/MM5_g
+ N_VDD_XI17/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI0/MM4 N_XI17/XI0/NET33_XI17/XI0/MM4_d N_XI17/XI0/NET34_XI17/XI0/MM4_g
+ N_VDD_XI17/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI0/MM10 N_XI17/XI0/NET35_XI17/XI0/MM10_d N_XI17/XI0/NET36_XI17/XI0/MM10_g
+ N_VDD_XI17/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI0/MM11 N_XI17/XI0/NET36_XI17/XI0/MM11_d N_XI17/XI0/NET35_XI17/XI0/MM11_g
+ N_VDD_XI17/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI1/MM2 N_XI17/XI1/NET34_XI17/XI1/MM2_d N_XI17/XI1/NET33_XI17/XI1/MM2_g
+ N_VSS_XI17/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI1/MM3 N_XI17/XI1/NET33_XI17/XI1/MM3_d N_WL<30>_XI17/XI1/MM3_g
+ N_BLN<14>_XI17/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI1/MM0 N_XI17/XI1/NET34_XI17/XI1/MM0_d N_WL<30>_XI17/XI1/MM0_g
+ N_BL<14>_XI17/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI1/MM1 N_XI17/XI1/NET33_XI17/XI1/MM1_d N_XI17/XI1/NET34_XI17/XI1/MM1_g
+ N_VSS_XI17/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI1/MM9 N_XI17/XI1/NET36_XI17/XI1/MM9_d N_WL<31>_XI17/XI1/MM9_g
+ N_BL<14>_XI17/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI1/MM6 N_XI17/XI1/NET35_XI17/XI1/MM6_d N_XI17/XI1/NET36_XI17/XI1/MM6_g
+ N_VSS_XI17/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI1/MM7 N_XI17/XI1/NET36_XI17/XI1/MM7_d N_XI17/XI1/NET35_XI17/XI1/MM7_g
+ N_VSS_XI17/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI1/MM8 N_XI17/XI1/NET35_XI17/XI1/MM8_d N_WL<31>_XI17/XI1/MM8_g
+ N_BLN<14>_XI17/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI1/MM5 N_XI17/XI1/NET34_XI17/XI1/MM5_d N_XI17/XI1/NET33_XI17/XI1/MM5_g
+ N_VDD_XI17/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI1/MM4 N_XI17/XI1/NET33_XI17/XI1/MM4_d N_XI17/XI1/NET34_XI17/XI1/MM4_g
+ N_VDD_XI17/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI1/MM10 N_XI17/XI1/NET35_XI17/XI1/MM10_d N_XI17/XI1/NET36_XI17/XI1/MM10_g
+ N_VDD_XI17/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI1/MM11 N_XI17/XI1/NET36_XI17/XI1/MM11_d N_XI17/XI1/NET35_XI17/XI1/MM11_g
+ N_VDD_XI17/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI2/MM2 N_XI17/XI2/NET34_XI17/XI2/MM2_d N_XI17/XI2/NET33_XI17/XI2/MM2_g
+ N_VSS_XI17/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI2/MM3 N_XI17/XI2/NET33_XI17/XI2/MM3_d N_WL<30>_XI17/XI2/MM3_g
+ N_BLN<13>_XI17/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI2/MM0 N_XI17/XI2/NET34_XI17/XI2/MM0_d N_WL<30>_XI17/XI2/MM0_g
+ N_BL<13>_XI17/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI2/MM1 N_XI17/XI2/NET33_XI17/XI2/MM1_d N_XI17/XI2/NET34_XI17/XI2/MM1_g
+ N_VSS_XI17/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI2/MM9 N_XI17/XI2/NET36_XI17/XI2/MM9_d N_WL<31>_XI17/XI2/MM9_g
+ N_BL<13>_XI17/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI2/MM6 N_XI17/XI2/NET35_XI17/XI2/MM6_d N_XI17/XI2/NET36_XI17/XI2/MM6_g
+ N_VSS_XI17/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI2/MM7 N_XI17/XI2/NET36_XI17/XI2/MM7_d N_XI17/XI2/NET35_XI17/XI2/MM7_g
+ N_VSS_XI17/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI2/MM8 N_XI17/XI2/NET35_XI17/XI2/MM8_d N_WL<31>_XI17/XI2/MM8_g
+ N_BLN<13>_XI17/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI2/MM5 N_XI17/XI2/NET34_XI17/XI2/MM5_d N_XI17/XI2/NET33_XI17/XI2/MM5_g
+ N_VDD_XI17/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI2/MM4 N_XI17/XI2/NET33_XI17/XI2/MM4_d N_XI17/XI2/NET34_XI17/XI2/MM4_g
+ N_VDD_XI17/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI2/MM10 N_XI17/XI2/NET35_XI17/XI2/MM10_d N_XI17/XI2/NET36_XI17/XI2/MM10_g
+ N_VDD_XI17/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI2/MM11 N_XI17/XI2/NET36_XI17/XI2/MM11_d N_XI17/XI2/NET35_XI17/XI2/MM11_g
+ N_VDD_XI17/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI3/MM2 N_XI17/XI3/NET34_XI17/XI3/MM2_d N_XI17/XI3/NET33_XI17/XI3/MM2_g
+ N_VSS_XI17/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI3/MM3 N_XI17/XI3/NET33_XI17/XI3/MM3_d N_WL<30>_XI17/XI3/MM3_g
+ N_BLN<12>_XI17/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI3/MM0 N_XI17/XI3/NET34_XI17/XI3/MM0_d N_WL<30>_XI17/XI3/MM0_g
+ N_BL<12>_XI17/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI3/MM1 N_XI17/XI3/NET33_XI17/XI3/MM1_d N_XI17/XI3/NET34_XI17/XI3/MM1_g
+ N_VSS_XI17/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI3/MM9 N_XI17/XI3/NET36_XI17/XI3/MM9_d N_WL<31>_XI17/XI3/MM9_g
+ N_BL<12>_XI17/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI3/MM6 N_XI17/XI3/NET35_XI17/XI3/MM6_d N_XI17/XI3/NET36_XI17/XI3/MM6_g
+ N_VSS_XI17/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI3/MM7 N_XI17/XI3/NET36_XI17/XI3/MM7_d N_XI17/XI3/NET35_XI17/XI3/MM7_g
+ N_VSS_XI17/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI3/MM8 N_XI17/XI3/NET35_XI17/XI3/MM8_d N_WL<31>_XI17/XI3/MM8_g
+ N_BLN<12>_XI17/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI3/MM5 N_XI17/XI3/NET34_XI17/XI3/MM5_d N_XI17/XI3/NET33_XI17/XI3/MM5_g
+ N_VDD_XI17/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI3/MM4 N_XI17/XI3/NET33_XI17/XI3/MM4_d N_XI17/XI3/NET34_XI17/XI3/MM4_g
+ N_VDD_XI17/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI3/MM10 N_XI17/XI3/NET35_XI17/XI3/MM10_d N_XI17/XI3/NET36_XI17/XI3/MM10_g
+ N_VDD_XI17/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI3/MM11 N_XI17/XI3/NET36_XI17/XI3/MM11_d N_XI17/XI3/NET35_XI17/XI3/MM11_g
+ N_VDD_XI17/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI4/MM2 N_XI17/XI4/NET34_XI17/XI4/MM2_d N_XI17/XI4/NET33_XI17/XI4/MM2_g
+ N_VSS_XI17/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI4/MM3 N_XI17/XI4/NET33_XI17/XI4/MM3_d N_WL<30>_XI17/XI4/MM3_g
+ N_BLN<11>_XI17/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI4/MM0 N_XI17/XI4/NET34_XI17/XI4/MM0_d N_WL<30>_XI17/XI4/MM0_g
+ N_BL<11>_XI17/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI4/MM1 N_XI17/XI4/NET33_XI17/XI4/MM1_d N_XI17/XI4/NET34_XI17/XI4/MM1_g
+ N_VSS_XI17/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI4/MM9 N_XI17/XI4/NET36_XI17/XI4/MM9_d N_WL<31>_XI17/XI4/MM9_g
+ N_BL<11>_XI17/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI4/MM6 N_XI17/XI4/NET35_XI17/XI4/MM6_d N_XI17/XI4/NET36_XI17/XI4/MM6_g
+ N_VSS_XI17/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI4/MM7 N_XI17/XI4/NET36_XI17/XI4/MM7_d N_XI17/XI4/NET35_XI17/XI4/MM7_g
+ N_VSS_XI17/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI4/MM8 N_XI17/XI4/NET35_XI17/XI4/MM8_d N_WL<31>_XI17/XI4/MM8_g
+ N_BLN<11>_XI17/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI4/MM5 N_XI17/XI4/NET34_XI17/XI4/MM5_d N_XI17/XI4/NET33_XI17/XI4/MM5_g
+ N_VDD_XI17/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI4/MM4 N_XI17/XI4/NET33_XI17/XI4/MM4_d N_XI17/XI4/NET34_XI17/XI4/MM4_g
+ N_VDD_XI17/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI4/MM10 N_XI17/XI4/NET35_XI17/XI4/MM10_d N_XI17/XI4/NET36_XI17/XI4/MM10_g
+ N_VDD_XI17/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI4/MM11 N_XI17/XI4/NET36_XI17/XI4/MM11_d N_XI17/XI4/NET35_XI17/XI4/MM11_g
+ N_VDD_XI17/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI5/MM2 N_XI17/XI5/NET34_XI17/XI5/MM2_d N_XI17/XI5/NET33_XI17/XI5/MM2_g
+ N_VSS_XI17/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI5/MM3 N_XI17/XI5/NET33_XI17/XI5/MM3_d N_WL<30>_XI17/XI5/MM3_g
+ N_BLN<10>_XI17/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI5/MM0 N_XI17/XI5/NET34_XI17/XI5/MM0_d N_WL<30>_XI17/XI5/MM0_g
+ N_BL<10>_XI17/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI5/MM1 N_XI17/XI5/NET33_XI17/XI5/MM1_d N_XI17/XI5/NET34_XI17/XI5/MM1_g
+ N_VSS_XI17/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI5/MM9 N_XI17/XI5/NET36_XI17/XI5/MM9_d N_WL<31>_XI17/XI5/MM9_g
+ N_BL<10>_XI17/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI5/MM6 N_XI17/XI5/NET35_XI17/XI5/MM6_d N_XI17/XI5/NET36_XI17/XI5/MM6_g
+ N_VSS_XI17/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI5/MM7 N_XI17/XI5/NET36_XI17/XI5/MM7_d N_XI17/XI5/NET35_XI17/XI5/MM7_g
+ N_VSS_XI17/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI5/MM8 N_XI17/XI5/NET35_XI17/XI5/MM8_d N_WL<31>_XI17/XI5/MM8_g
+ N_BLN<10>_XI17/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI5/MM5 N_XI17/XI5/NET34_XI17/XI5/MM5_d N_XI17/XI5/NET33_XI17/XI5/MM5_g
+ N_VDD_XI17/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI5/MM4 N_XI17/XI5/NET33_XI17/XI5/MM4_d N_XI17/XI5/NET34_XI17/XI5/MM4_g
+ N_VDD_XI17/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI5/MM10 N_XI17/XI5/NET35_XI17/XI5/MM10_d N_XI17/XI5/NET36_XI17/XI5/MM10_g
+ N_VDD_XI17/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI5/MM11 N_XI17/XI5/NET36_XI17/XI5/MM11_d N_XI17/XI5/NET35_XI17/XI5/MM11_g
+ N_VDD_XI17/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI6/MM2 N_XI17/XI6/NET34_XI17/XI6/MM2_d N_XI17/XI6/NET33_XI17/XI6/MM2_g
+ N_VSS_XI17/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM3 N_XI17/XI6/NET33_XI17/XI6/MM3_d N_WL<30>_XI17/XI6/MM3_g
+ N_BLN<9>_XI17/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM0 N_XI17/XI6/NET34_XI17/XI6/MM0_d N_WL<30>_XI17/XI6/MM0_g
+ N_BL<9>_XI17/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM1 N_XI17/XI6/NET33_XI17/XI6/MM1_d N_XI17/XI6/NET34_XI17/XI6/MM1_g
+ N_VSS_XI17/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM9 N_XI17/XI6/NET36_XI17/XI6/MM9_d N_WL<31>_XI17/XI6/MM9_g
+ N_BL<9>_XI17/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM6 N_XI17/XI6/NET35_XI17/XI6/MM6_d N_XI17/XI6/NET36_XI17/XI6/MM6_g
+ N_VSS_XI17/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM7 N_XI17/XI6/NET36_XI17/XI6/MM7_d N_XI17/XI6/NET35_XI17/XI6/MM7_g
+ N_VSS_XI17/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM8 N_XI17/XI6/NET35_XI17/XI6/MM8_d N_WL<31>_XI17/XI6/MM8_g
+ N_BLN<9>_XI17/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI6/MM5 N_XI17/XI6/NET34_XI17/XI6/MM5_d N_XI17/XI6/NET33_XI17/XI6/MM5_g
+ N_VDD_XI17/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI6/MM4 N_XI17/XI6/NET33_XI17/XI6/MM4_d N_XI17/XI6/NET34_XI17/XI6/MM4_g
+ N_VDD_XI17/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI6/MM10 N_XI17/XI6/NET35_XI17/XI6/MM10_d N_XI17/XI6/NET36_XI17/XI6/MM10_g
+ N_VDD_XI17/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI6/MM11 N_XI17/XI6/NET36_XI17/XI6/MM11_d N_XI17/XI6/NET35_XI17/XI6/MM11_g
+ N_VDD_XI17/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI7/MM2 N_XI17/XI7/NET34_XI17/XI7/MM2_d N_XI17/XI7/NET33_XI17/XI7/MM2_g
+ N_VSS_XI17/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM3 N_XI17/XI7/NET33_XI17/XI7/MM3_d N_WL<30>_XI17/XI7/MM3_g
+ N_BLN<8>_XI17/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM0 N_XI17/XI7/NET34_XI17/XI7/MM0_d N_WL<30>_XI17/XI7/MM0_g
+ N_BL<8>_XI17/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM1 N_XI17/XI7/NET33_XI17/XI7/MM1_d N_XI17/XI7/NET34_XI17/XI7/MM1_g
+ N_VSS_XI17/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM9 N_XI17/XI7/NET36_XI17/XI7/MM9_d N_WL<31>_XI17/XI7/MM9_g
+ N_BL<8>_XI17/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM6 N_XI17/XI7/NET35_XI17/XI7/MM6_d N_XI17/XI7/NET36_XI17/XI7/MM6_g
+ N_VSS_XI17/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM7 N_XI17/XI7/NET36_XI17/XI7/MM7_d N_XI17/XI7/NET35_XI17/XI7/MM7_g
+ N_VSS_XI17/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM8 N_XI17/XI7/NET35_XI17/XI7/MM8_d N_WL<31>_XI17/XI7/MM8_g
+ N_BLN<8>_XI17/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI7/MM5 N_XI17/XI7/NET34_XI17/XI7/MM5_d N_XI17/XI7/NET33_XI17/XI7/MM5_g
+ N_VDD_XI17/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI7/MM4 N_XI17/XI7/NET33_XI17/XI7/MM4_d N_XI17/XI7/NET34_XI17/XI7/MM4_g
+ N_VDD_XI17/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI7/MM10 N_XI17/XI7/NET35_XI17/XI7/MM10_d N_XI17/XI7/NET36_XI17/XI7/MM10_g
+ N_VDD_XI17/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI7/MM11 N_XI17/XI7/NET36_XI17/XI7/MM11_d N_XI17/XI7/NET35_XI17/XI7/MM11_g
+ N_VDD_XI17/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI8/MM2 N_XI17/XI8/NET34_XI17/XI8/MM2_d N_XI17/XI8/NET33_XI17/XI8/MM2_g
+ N_VSS_XI17/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM3 N_XI17/XI8/NET33_XI17/XI8/MM3_d N_WL<30>_XI17/XI8/MM3_g
+ N_BLN<7>_XI17/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM0 N_XI17/XI8/NET34_XI17/XI8/MM0_d N_WL<30>_XI17/XI8/MM0_g
+ N_BL<7>_XI17/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM1 N_XI17/XI8/NET33_XI17/XI8/MM1_d N_XI17/XI8/NET34_XI17/XI8/MM1_g
+ N_VSS_XI17/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM9 N_XI17/XI8/NET36_XI17/XI8/MM9_d N_WL<31>_XI17/XI8/MM9_g
+ N_BL<7>_XI17/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM6 N_XI17/XI8/NET35_XI17/XI8/MM6_d N_XI17/XI8/NET36_XI17/XI8/MM6_g
+ N_VSS_XI17/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM7 N_XI17/XI8/NET36_XI17/XI8/MM7_d N_XI17/XI8/NET35_XI17/XI8/MM7_g
+ N_VSS_XI17/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM8 N_XI17/XI8/NET35_XI17/XI8/MM8_d N_WL<31>_XI17/XI8/MM8_g
+ N_BLN<7>_XI17/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI8/MM5 N_XI17/XI8/NET34_XI17/XI8/MM5_d N_XI17/XI8/NET33_XI17/XI8/MM5_g
+ N_VDD_XI17/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI8/MM4 N_XI17/XI8/NET33_XI17/XI8/MM4_d N_XI17/XI8/NET34_XI17/XI8/MM4_g
+ N_VDD_XI17/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI8/MM10 N_XI17/XI8/NET35_XI17/XI8/MM10_d N_XI17/XI8/NET36_XI17/XI8/MM10_g
+ N_VDD_XI17/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI8/MM11 N_XI17/XI8/NET36_XI17/XI8/MM11_d N_XI17/XI8/NET35_XI17/XI8/MM11_g
+ N_VDD_XI17/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI9/MM2 N_XI17/XI9/NET34_XI17/XI9/MM2_d N_XI17/XI9/NET33_XI17/XI9/MM2_g
+ N_VSS_XI17/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM3 N_XI17/XI9/NET33_XI17/XI9/MM3_d N_WL<30>_XI17/XI9/MM3_g
+ N_BLN<6>_XI17/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM0 N_XI17/XI9/NET34_XI17/XI9/MM0_d N_WL<30>_XI17/XI9/MM0_g
+ N_BL<6>_XI17/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM1 N_XI17/XI9/NET33_XI17/XI9/MM1_d N_XI17/XI9/NET34_XI17/XI9/MM1_g
+ N_VSS_XI17/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM9 N_XI17/XI9/NET36_XI17/XI9/MM9_d N_WL<31>_XI17/XI9/MM9_g
+ N_BL<6>_XI17/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM6 N_XI17/XI9/NET35_XI17/XI9/MM6_d N_XI17/XI9/NET36_XI17/XI9/MM6_g
+ N_VSS_XI17/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM7 N_XI17/XI9/NET36_XI17/XI9/MM7_d N_XI17/XI9/NET35_XI17/XI9/MM7_g
+ N_VSS_XI17/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM8 N_XI17/XI9/NET35_XI17/XI9/MM8_d N_WL<31>_XI17/XI9/MM8_g
+ N_BLN<6>_XI17/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI9/MM5 N_XI17/XI9/NET34_XI17/XI9/MM5_d N_XI17/XI9/NET33_XI17/XI9/MM5_g
+ N_VDD_XI17/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI9/MM4 N_XI17/XI9/NET33_XI17/XI9/MM4_d N_XI17/XI9/NET34_XI17/XI9/MM4_g
+ N_VDD_XI17/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI9/MM10 N_XI17/XI9/NET35_XI17/XI9/MM10_d N_XI17/XI9/NET36_XI17/XI9/MM10_g
+ N_VDD_XI17/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI9/MM11 N_XI17/XI9/NET36_XI17/XI9/MM11_d N_XI17/XI9/NET35_XI17/XI9/MM11_g
+ N_VDD_XI17/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI10/MM2 N_XI17/XI10/NET34_XI17/XI10/MM2_d
+ N_XI17/XI10/NET33_XI17/XI10/MM2_g N_VSS_XI17/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI10/MM3 N_XI17/XI10/NET33_XI17/XI10/MM3_d N_WL<30>_XI17/XI10/MM3_g
+ N_BLN<5>_XI17/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI10/MM0 N_XI17/XI10/NET34_XI17/XI10/MM0_d N_WL<30>_XI17/XI10/MM0_g
+ N_BL<5>_XI17/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI10/MM1 N_XI17/XI10/NET33_XI17/XI10/MM1_d
+ N_XI17/XI10/NET34_XI17/XI10/MM1_g N_VSS_XI17/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI10/MM9 N_XI17/XI10/NET36_XI17/XI10/MM9_d N_WL<31>_XI17/XI10/MM9_g
+ N_BL<5>_XI17/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI10/MM6 N_XI17/XI10/NET35_XI17/XI10/MM6_d
+ N_XI17/XI10/NET36_XI17/XI10/MM6_g N_VSS_XI17/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI10/MM7 N_XI17/XI10/NET36_XI17/XI10/MM7_d
+ N_XI17/XI10/NET35_XI17/XI10/MM7_g N_VSS_XI17/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI10/MM8 N_XI17/XI10/NET35_XI17/XI10/MM8_d N_WL<31>_XI17/XI10/MM8_g
+ N_BLN<5>_XI17/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI10/MM5 N_XI17/XI10/NET34_XI17/XI10/MM5_d
+ N_XI17/XI10/NET33_XI17/XI10/MM5_g N_VDD_XI17/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI10/MM4 N_XI17/XI10/NET33_XI17/XI10/MM4_d
+ N_XI17/XI10/NET34_XI17/XI10/MM4_g N_VDD_XI17/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI10/MM10 N_XI17/XI10/NET35_XI17/XI10/MM10_d
+ N_XI17/XI10/NET36_XI17/XI10/MM10_g N_VDD_XI17/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI10/MM11 N_XI17/XI10/NET36_XI17/XI10/MM11_d
+ N_XI17/XI10/NET35_XI17/XI10/MM11_g N_VDD_XI17/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI11/MM2 N_XI17/XI11/NET34_XI17/XI11/MM2_d
+ N_XI17/XI11/NET33_XI17/XI11/MM2_g N_VSS_XI17/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI11/MM3 N_XI17/XI11/NET33_XI17/XI11/MM3_d N_WL<30>_XI17/XI11/MM3_g
+ N_BLN<4>_XI17/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI11/MM0 N_XI17/XI11/NET34_XI17/XI11/MM0_d N_WL<30>_XI17/XI11/MM0_g
+ N_BL<4>_XI17/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI11/MM1 N_XI17/XI11/NET33_XI17/XI11/MM1_d
+ N_XI17/XI11/NET34_XI17/XI11/MM1_g N_VSS_XI17/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI11/MM9 N_XI17/XI11/NET36_XI17/XI11/MM9_d N_WL<31>_XI17/XI11/MM9_g
+ N_BL<4>_XI17/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI11/MM6 N_XI17/XI11/NET35_XI17/XI11/MM6_d
+ N_XI17/XI11/NET36_XI17/XI11/MM6_g N_VSS_XI17/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI11/MM7 N_XI17/XI11/NET36_XI17/XI11/MM7_d
+ N_XI17/XI11/NET35_XI17/XI11/MM7_g N_VSS_XI17/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI11/MM8 N_XI17/XI11/NET35_XI17/XI11/MM8_d N_WL<31>_XI17/XI11/MM8_g
+ N_BLN<4>_XI17/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI11/MM5 N_XI17/XI11/NET34_XI17/XI11/MM5_d
+ N_XI17/XI11/NET33_XI17/XI11/MM5_g N_VDD_XI17/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI11/MM4 N_XI17/XI11/NET33_XI17/XI11/MM4_d
+ N_XI17/XI11/NET34_XI17/XI11/MM4_g N_VDD_XI17/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI11/MM10 N_XI17/XI11/NET35_XI17/XI11/MM10_d
+ N_XI17/XI11/NET36_XI17/XI11/MM10_g N_VDD_XI17/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI11/MM11 N_XI17/XI11/NET36_XI17/XI11/MM11_d
+ N_XI17/XI11/NET35_XI17/XI11/MM11_g N_VDD_XI17/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI12/MM2 N_XI17/XI12/NET34_XI17/XI12/MM2_d
+ N_XI17/XI12/NET33_XI17/XI12/MM2_g N_VSS_XI17/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI12/MM3 N_XI17/XI12/NET33_XI17/XI12/MM3_d N_WL<30>_XI17/XI12/MM3_g
+ N_BLN<3>_XI17/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI12/MM0 N_XI17/XI12/NET34_XI17/XI12/MM0_d N_WL<30>_XI17/XI12/MM0_g
+ N_BL<3>_XI17/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI12/MM1 N_XI17/XI12/NET33_XI17/XI12/MM1_d
+ N_XI17/XI12/NET34_XI17/XI12/MM1_g N_VSS_XI17/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI12/MM9 N_XI17/XI12/NET36_XI17/XI12/MM9_d N_WL<31>_XI17/XI12/MM9_g
+ N_BL<3>_XI17/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI12/MM6 N_XI17/XI12/NET35_XI17/XI12/MM6_d
+ N_XI17/XI12/NET36_XI17/XI12/MM6_g N_VSS_XI17/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI12/MM7 N_XI17/XI12/NET36_XI17/XI12/MM7_d
+ N_XI17/XI12/NET35_XI17/XI12/MM7_g N_VSS_XI17/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI12/MM8 N_XI17/XI12/NET35_XI17/XI12/MM8_d N_WL<31>_XI17/XI12/MM8_g
+ N_BLN<3>_XI17/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI12/MM5 N_XI17/XI12/NET34_XI17/XI12/MM5_d
+ N_XI17/XI12/NET33_XI17/XI12/MM5_g N_VDD_XI17/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI12/MM4 N_XI17/XI12/NET33_XI17/XI12/MM4_d
+ N_XI17/XI12/NET34_XI17/XI12/MM4_g N_VDD_XI17/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI12/MM10 N_XI17/XI12/NET35_XI17/XI12/MM10_d
+ N_XI17/XI12/NET36_XI17/XI12/MM10_g N_VDD_XI17/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI12/MM11 N_XI17/XI12/NET36_XI17/XI12/MM11_d
+ N_XI17/XI12/NET35_XI17/XI12/MM11_g N_VDD_XI17/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI13/MM2 N_XI17/XI13/NET34_XI17/XI13/MM2_d
+ N_XI17/XI13/NET33_XI17/XI13/MM2_g N_VSS_XI17/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI13/MM3 N_XI17/XI13/NET33_XI17/XI13/MM3_d N_WL<30>_XI17/XI13/MM3_g
+ N_BLN<2>_XI17/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI13/MM0 N_XI17/XI13/NET34_XI17/XI13/MM0_d N_WL<30>_XI17/XI13/MM0_g
+ N_BL<2>_XI17/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI13/MM1 N_XI17/XI13/NET33_XI17/XI13/MM1_d
+ N_XI17/XI13/NET34_XI17/XI13/MM1_g N_VSS_XI17/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI13/MM9 N_XI17/XI13/NET36_XI17/XI13/MM9_d N_WL<31>_XI17/XI13/MM9_g
+ N_BL<2>_XI17/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI13/MM6 N_XI17/XI13/NET35_XI17/XI13/MM6_d
+ N_XI17/XI13/NET36_XI17/XI13/MM6_g N_VSS_XI17/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI13/MM7 N_XI17/XI13/NET36_XI17/XI13/MM7_d
+ N_XI17/XI13/NET35_XI17/XI13/MM7_g N_VSS_XI17/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI13/MM8 N_XI17/XI13/NET35_XI17/XI13/MM8_d N_WL<31>_XI17/XI13/MM8_g
+ N_BLN<2>_XI17/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI13/MM5 N_XI17/XI13/NET34_XI17/XI13/MM5_d
+ N_XI17/XI13/NET33_XI17/XI13/MM5_g N_VDD_XI17/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI13/MM4 N_XI17/XI13/NET33_XI17/XI13/MM4_d
+ N_XI17/XI13/NET34_XI17/XI13/MM4_g N_VDD_XI17/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI13/MM10 N_XI17/XI13/NET35_XI17/XI13/MM10_d
+ N_XI17/XI13/NET36_XI17/XI13/MM10_g N_VDD_XI17/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI13/MM11 N_XI17/XI13/NET36_XI17/XI13/MM11_d
+ N_XI17/XI13/NET35_XI17/XI13/MM11_g N_VDD_XI17/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI14/MM2 N_XI17/XI14/NET34_XI17/XI14/MM2_d
+ N_XI17/XI14/NET33_XI17/XI14/MM2_g N_VSS_XI17/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI14/MM3 N_XI17/XI14/NET33_XI17/XI14/MM3_d N_WL<30>_XI17/XI14/MM3_g
+ N_BLN<1>_XI17/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI14/MM0 N_XI17/XI14/NET34_XI17/XI14/MM0_d N_WL<30>_XI17/XI14/MM0_g
+ N_BL<1>_XI17/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI14/MM1 N_XI17/XI14/NET33_XI17/XI14/MM1_d
+ N_XI17/XI14/NET34_XI17/XI14/MM1_g N_VSS_XI17/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI14/MM9 N_XI17/XI14/NET36_XI17/XI14/MM9_d N_WL<31>_XI17/XI14/MM9_g
+ N_BL<1>_XI17/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI14/MM6 N_XI17/XI14/NET35_XI17/XI14/MM6_d
+ N_XI17/XI14/NET36_XI17/XI14/MM6_g N_VSS_XI17/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI14/MM7 N_XI17/XI14/NET36_XI17/XI14/MM7_d
+ N_XI17/XI14/NET35_XI17/XI14/MM7_g N_VSS_XI17/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI14/MM8 N_XI17/XI14/NET35_XI17/XI14/MM8_d N_WL<31>_XI17/XI14/MM8_g
+ N_BLN<1>_XI17/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI14/MM5 N_XI17/XI14/NET34_XI17/XI14/MM5_d
+ N_XI17/XI14/NET33_XI17/XI14/MM5_g N_VDD_XI17/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI14/MM4 N_XI17/XI14/NET33_XI17/XI14/MM4_d
+ N_XI17/XI14/NET34_XI17/XI14/MM4_g N_VDD_XI17/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI14/MM10 N_XI17/XI14/NET35_XI17/XI14/MM10_d
+ N_XI17/XI14/NET36_XI17/XI14/MM10_g N_VDD_XI17/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI14/MM11 N_XI17/XI14/NET36_XI17/XI14/MM11_d
+ N_XI17/XI14/NET35_XI17/XI14/MM11_g N_VDD_XI17/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI15/MM2 N_XI17/XI15/NET34_XI17/XI15/MM2_d
+ N_XI17/XI15/NET33_XI17/XI15/MM2_g N_VSS_XI17/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI15/MM3 N_XI17/XI15/NET33_XI17/XI15/MM3_d N_WL<30>_XI17/XI15/MM3_g
+ N_BLN<0>_XI17/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI15/MM0 N_XI17/XI15/NET34_XI17/XI15/MM0_d N_WL<30>_XI17/XI15/MM0_g
+ N_BL<0>_XI17/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI15/MM1 N_XI17/XI15/NET33_XI17/XI15/MM1_d
+ N_XI17/XI15/NET34_XI17/XI15/MM1_g N_VSS_XI17/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI15/MM9 N_XI17/XI15/NET36_XI17/XI15/MM9_d N_WL<31>_XI17/XI15/MM9_g
+ N_BL<0>_XI17/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI15/MM6 N_XI17/XI15/NET35_XI17/XI15/MM6_d
+ N_XI17/XI15/NET36_XI17/XI15/MM6_g N_VSS_XI17/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI15/MM7 N_XI17/XI15/NET36_XI17/XI15/MM7_d
+ N_XI17/XI15/NET35_XI17/XI15/MM7_g N_VSS_XI17/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI17/XI15/MM8 N_XI17/XI15/NET35_XI17/XI15/MM8_d N_WL<31>_XI17/XI15/MM8_g
+ N_BLN<0>_XI17/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI17/XI15/MM5 N_XI17/XI15/NET34_XI17/XI15/MM5_d
+ N_XI17/XI15/NET33_XI17/XI15/MM5_g N_VDD_XI17/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI15/MM4 N_XI17/XI15/NET33_XI17/XI15/MM4_d
+ N_XI17/XI15/NET34_XI17/XI15/MM4_g N_VDD_XI17/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI15/MM10 N_XI17/XI15/NET35_XI17/XI15/MM10_d
+ N_XI17/XI15/NET36_XI17/XI15/MM10_g N_VDD_XI17/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI17/XI15/MM11 N_XI17/XI15/NET36_XI17/XI15/MM11_d
+ N_XI17/XI15/NET35_XI17/XI15/MM11_g N_VDD_XI17/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI0/MM2 N_XI18/XI0/NET34_XI18/XI0/MM2_d N_XI18/XI0/NET33_XI18/XI0/MM2_g
+ N_VSS_XI18/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI0/MM3 N_XI18/XI0/NET33_XI18/XI0/MM3_d N_WL<32>_XI18/XI0/MM3_g
+ N_BLN<15>_XI18/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI0/MM0 N_XI18/XI0/NET34_XI18/XI0/MM0_d N_WL<32>_XI18/XI0/MM0_g
+ N_BL<15>_XI18/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI0/MM1 N_XI18/XI0/NET33_XI18/XI0/MM1_d N_XI18/XI0/NET34_XI18/XI0/MM1_g
+ N_VSS_XI18/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI0/MM9 N_XI18/XI0/NET36_XI18/XI0/MM9_d N_WL<33>_XI18/XI0/MM9_g
+ N_BL<15>_XI18/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI0/MM6 N_XI18/XI0/NET35_XI18/XI0/MM6_d N_XI18/XI0/NET36_XI18/XI0/MM6_g
+ N_VSS_XI18/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI0/MM7 N_XI18/XI0/NET36_XI18/XI0/MM7_d N_XI18/XI0/NET35_XI18/XI0/MM7_g
+ N_VSS_XI18/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI0/MM8 N_XI18/XI0/NET35_XI18/XI0/MM8_d N_WL<33>_XI18/XI0/MM8_g
+ N_BLN<15>_XI18/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI0/MM5 N_XI18/XI0/NET34_XI18/XI0/MM5_d N_XI18/XI0/NET33_XI18/XI0/MM5_g
+ N_VDD_XI18/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI0/MM4 N_XI18/XI0/NET33_XI18/XI0/MM4_d N_XI18/XI0/NET34_XI18/XI0/MM4_g
+ N_VDD_XI18/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI0/MM10 N_XI18/XI0/NET35_XI18/XI0/MM10_d N_XI18/XI0/NET36_XI18/XI0/MM10_g
+ N_VDD_XI18/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI0/MM11 N_XI18/XI0/NET36_XI18/XI0/MM11_d N_XI18/XI0/NET35_XI18/XI0/MM11_g
+ N_VDD_XI18/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI1/MM2 N_XI18/XI1/NET34_XI18/XI1/MM2_d N_XI18/XI1/NET33_XI18/XI1/MM2_g
+ N_VSS_XI18/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI1/MM3 N_XI18/XI1/NET33_XI18/XI1/MM3_d N_WL<32>_XI18/XI1/MM3_g
+ N_BLN<14>_XI18/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI1/MM0 N_XI18/XI1/NET34_XI18/XI1/MM0_d N_WL<32>_XI18/XI1/MM0_g
+ N_BL<14>_XI18/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI1/MM1 N_XI18/XI1/NET33_XI18/XI1/MM1_d N_XI18/XI1/NET34_XI18/XI1/MM1_g
+ N_VSS_XI18/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI1/MM9 N_XI18/XI1/NET36_XI18/XI1/MM9_d N_WL<33>_XI18/XI1/MM9_g
+ N_BL<14>_XI18/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI1/MM6 N_XI18/XI1/NET35_XI18/XI1/MM6_d N_XI18/XI1/NET36_XI18/XI1/MM6_g
+ N_VSS_XI18/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI1/MM7 N_XI18/XI1/NET36_XI18/XI1/MM7_d N_XI18/XI1/NET35_XI18/XI1/MM7_g
+ N_VSS_XI18/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI1/MM8 N_XI18/XI1/NET35_XI18/XI1/MM8_d N_WL<33>_XI18/XI1/MM8_g
+ N_BLN<14>_XI18/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI1/MM5 N_XI18/XI1/NET34_XI18/XI1/MM5_d N_XI18/XI1/NET33_XI18/XI1/MM5_g
+ N_VDD_XI18/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI1/MM4 N_XI18/XI1/NET33_XI18/XI1/MM4_d N_XI18/XI1/NET34_XI18/XI1/MM4_g
+ N_VDD_XI18/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI1/MM10 N_XI18/XI1/NET35_XI18/XI1/MM10_d N_XI18/XI1/NET36_XI18/XI1/MM10_g
+ N_VDD_XI18/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI1/MM11 N_XI18/XI1/NET36_XI18/XI1/MM11_d N_XI18/XI1/NET35_XI18/XI1/MM11_g
+ N_VDD_XI18/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI2/MM2 N_XI18/XI2/NET34_XI18/XI2/MM2_d N_XI18/XI2/NET33_XI18/XI2/MM2_g
+ N_VSS_XI18/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI2/MM3 N_XI18/XI2/NET33_XI18/XI2/MM3_d N_WL<32>_XI18/XI2/MM3_g
+ N_BLN<13>_XI18/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI2/MM0 N_XI18/XI2/NET34_XI18/XI2/MM0_d N_WL<32>_XI18/XI2/MM0_g
+ N_BL<13>_XI18/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI2/MM1 N_XI18/XI2/NET33_XI18/XI2/MM1_d N_XI18/XI2/NET34_XI18/XI2/MM1_g
+ N_VSS_XI18/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI2/MM9 N_XI18/XI2/NET36_XI18/XI2/MM9_d N_WL<33>_XI18/XI2/MM9_g
+ N_BL<13>_XI18/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI2/MM6 N_XI18/XI2/NET35_XI18/XI2/MM6_d N_XI18/XI2/NET36_XI18/XI2/MM6_g
+ N_VSS_XI18/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI2/MM7 N_XI18/XI2/NET36_XI18/XI2/MM7_d N_XI18/XI2/NET35_XI18/XI2/MM7_g
+ N_VSS_XI18/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI2/MM8 N_XI18/XI2/NET35_XI18/XI2/MM8_d N_WL<33>_XI18/XI2/MM8_g
+ N_BLN<13>_XI18/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI2/MM5 N_XI18/XI2/NET34_XI18/XI2/MM5_d N_XI18/XI2/NET33_XI18/XI2/MM5_g
+ N_VDD_XI18/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI2/MM4 N_XI18/XI2/NET33_XI18/XI2/MM4_d N_XI18/XI2/NET34_XI18/XI2/MM4_g
+ N_VDD_XI18/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI2/MM10 N_XI18/XI2/NET35_XI18/XI2/MM10_d N_XI18/XI2/NET36_XI18/XI2/MM10_g
+ N_VDD_XI18/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI2/MM11 N_XI18/XI2/NET36_XI18/XI2/MM11_d N_XI18/XI2/NET35_XI18/XI2/MM11_g
+ N_VDD_XI18/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI3/MM2 N_XI18/XI3/NET34_XI18/XI3/MM2_d N_XI18/XI3/NET33_XI18/XI3/MM2_g
+ N_VSS_XI18/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI3/MM3 N_XI18/XI3/NET33_XI18/XI3/MM3_d N_WL<32>_XI18/XI3/MM3_g
+ N_BLN<12>_XI18/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI3/MM0 N_XI18/XI3/NET34_XI18/XI3/MM0_d N_WL<32>_XI18/XI3/MM0_g
+ N_BL<12>_XI18/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI3/MM1 N_XI18/XI3/NET33_XI18/XI3/MM1_d N_XI18/XI3/NET34_XI18/XI3/MM1_g
+ N_VSS_XI18/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI3/MM9 N_XI18/XI3/NET36_XI18/XI3/MM9_d N_WL<33>_XI18/XI3/MM9_g
+ N_BL<12>_XI18/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI3/MM6 N_XI18/XI3/NET35_XI18/XI3/MM6_d N_XI18/XI3/NET36_XI18/XI3/MM6_g
+ N_VSS_XI18/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI3/MM7 N_XI18/XI3/NET36_XI18/XI3/MM7_d N_XI18/XI3/NET35_XI18/XI3/MM7_g
+ N_VSS_XI18/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI3/MM8 N_XI18/XI3/NET35_XI18/XI3/MM8_d N_WL<33>_XI18/XI3/MM8_g
+ N_BLN<12>_XI18/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI3/MM5 N_XI18/XI3/NET34_XI18/XI3/MM5_d N_XI18/XI3/NET33_XI18/XI3/MM5_g
+ N_VDD_XI18/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI3/MM4 N_XI18/XI3/NET33_XI18/XI3/MM4_d N_XI18/XI3/NET34_XI18/XI3/MM4_g
+ N_VDD_XI18/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI3/MM10 N_XI18/XI3/NET35_XI18/XI3/MM10_d N_XI18/XI3/NET36_XI18/XI3/MM10_g
+ N_VDD_XI18/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI3/MM11 N_XI18/XI3/NET36_XI18/XI3/MM11_d N_XI18/XI3/NET35_XI18/XI3/MM11_g
+ N_VDD_XI18/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI4/MM2 N_XI18/XI4/NET34_XI18/XI4/MM2_d N_XI18/XI4/NET33_XI18/XI4/MM2_g
+ N_VSS_XI18/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI4/MM3 N_XI18/XI4/NET33_XI18/XI4/MM3_d N_WL<32>_XI18/XI4/MM3_g
+ N_BLN<11>_XI18/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI4/MM0 N_XI18/XI4/NET34_XI18/XI4/MM0_d N_WL<32>_XI18/XI4/MM0_g
+ N_BL<11>_XI18/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI4/MM1 N_XI18/XI4/NET33_XI18/XI4/MM1_d N_XI18/XI4/NET34_XI18/XI4/MM1_g
+ N_VSS_XI18/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI4/MM9 N_XI18/XI4/NET36_XI18/XI4/MM9_d N_WL<33>_XI18/XI4/MM9_g
+ N_BL<11>_XI18/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI4/MM6 N_XI18/XI4/NET35_XI18/XI4/MM6_d N_XI18/XI4/NET36_XI18/XI4/MM6_g
+ N_VSS_XI18/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI4/MM7 N_XI18/XI4/NET36_XI18/XI4/MM7_d N_XI18/XI4/NET35_XI18/XI4/MM7_g
+ N_VSS_XI18/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI4/MM8 N_XI18/XI4/NET35_XI18/XI4/MM8_d N_WL<33>_XI18/XI4/MM8_g
+ N_BLN<11>_XI18/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI4/MM5 N_XI18/XI4/NET34_XI18/XI4/MM5_d N_XI18/XI4/NET33_XI18/XI4/MM5_g
+ N_VDD_XI18/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI4/MM4 N_XI18/XI4/NET33_XI18/XI4/MM4_d N_XI18/XI4/NET34_XI18/XI4/MM4_g
+ N_VDD_XI18/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI4/MM10 N_XI18/XI4/NET35_XI18/XI4/MM10_d N_XI18/XI4/NET36_XI18/XI4/MM10_g
+ N_VDD_XI18/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI4/MM11 N_XI18/XI4/NET36_XI18/XI4/MM11_d N_XI18/XI4/NET35_XI18/XI4/MM11_g
+ N_VDD_XI18/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI5/MM2 N_XI18/XI5/NET34_XI18/XI5/MM2_d N_XI18/XI5/NET33_XI18/XI5/MM2_g
+ N_VSS_XI18/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI5/MM3 N_XI18/XI5/NET33_XI18/XI5/MM3_d N_WL<32>_XI18/XI5/MM3_g
+ N_BLN<10>_XI18/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI5/MM0 N_XI18/XI5/NET34_XI18/XI5/MM0_d N_WL<32>_XI18/XI5/MM0_g
+ N_BL<10>_XI18/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI5/MM1 N_XI18/XI5/NET33_XI18/XI5/MM1_d N_XI18/XI5/NET34_XI18/XI5/MM1_g
+ N_VSS_XI18/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI5/MM9 N_XI18/XI5/NET36_XI18/XI5/MM9_d N_WL<33>_XI18/XI5/MM9_g
+ N_BL<10>_XI18/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI5/MM6 N_XI18/XI5/NET35_XI18/XI5/MM6_d N_XI18/XI5/NET36_XI18/XI5/MM6_g
+ N_VSS_XI18/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI5/MM7 N_XI18/XI5/NET36_XI18/XI5/MM7_d N_XI18/XI5/NET35_XI18/XI5/MM7_g
+ N_VSS_XI18/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI5/MM8 N_XI18/XI5/NET35_XI18/XI5/MM8_d N_WL<33>_XI18/XI5/MM8_g
+ N_BLN<10>_XI18/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI5/MM5 N_XI18/XI5/NET34_XI18/XI5/MM5_d N_XI18/XI5/NET33_XI18/XI5/MM5_g
+ N_VDD_XI18/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI5/MM4 N_XI18/XI5/NET33_XI18/XI5/MM4_d N_XI18/XI5/NET34_XI18/XI5/MM4_g
+ N_VDD_XI18/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI5/MM10 N_XI18/XI5/NET35_XI18/XI5/MM10_d N_XI18/XI5/NET36_XI18/XI5/MM10_g
+ N_VDD_XI18/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI5/MM11 N_XI18/XI5/NET36_XI18/XI5/MM11_d N_XI18/XI5/NET35_XI18/XI5/MM11_g
+ N_VDD_XI18/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI6/MM2 N_XI18/XI6/NET34_XI18/XI6/MM2_d N_XI18/XI6/NET33_XI18/XI6/MM2_g
+ N_VSS_XI18/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM3 N_XI18/XI6/NET33_XI18/XI6/MM3_d N_WL<32>_XI18/XI6/MM3_g
+ N_BLN<9>_XI18/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM0 N_XI18/XI6/NET34_XI18/XI6/MM0_d N_WL<32>_XI18/XI6/MM0_g
+ N_BL<9>_XI18/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM1 N_XI18/XI6/NET33_XI18/XI6/MM1_d N_XI18/XI6/NET34_XI18/XI6/MM1_g
+ N_VSS_XI18/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM9 N_XI18/XI6/NET36_XI18/XI6/MM9_d N_WL<33>_XI18/XI6/MM9_g
+ N_BL<9>_XI18/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM6 N_XI18/XI6/NET35_XI18/XI6/MM6_d N_XI18/XI6/NET36_XI18/XI6/MM6_g
+ N_VSS_XI18/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM7 N_XI18/XI6/NET36_XI18/XI6/MM7_d N_XI18/XI6/NET35_XI18/XI6/MM7_g
+ N_VSS_XI18/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM8 N_XI18/XI6/NET35_XI18/XI6/MM8_d N_WL<33>_XI18/XI6/MM8_g
+ N_BLN<9>_XI18/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI6/MM5 N_XI18/XI6/NET34_XI18/XI6/MM5_d N_XI18/XI6/NET33_XI18/XI6/MM5_g
+ N_VDD_XI18/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI6/MM4 N_XI18/XI6/NET33_XI18/XI6/MM4_d N_XI18/XI6/NET34_XI18/XI6/MM4_g
+ N_VDD_XI18/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI6/MM10 N_XI18/XI6/NET35_XI18/XI6/MM10_d N_XI18/XI6/NET36_XI18/XI6/MM10_g
+ N_VDD_XI18/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI6/MM11 N_XI18/XI6/NET36_XI18/XI6/MM11_d N_XI18/XI6/NET35_XI18/XI6/MM11_g
+ N_VDD_XI18/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI7/MM2 N_XI18/XI7/NET34_XI18/XI7/MM2_d N_XI18/XI7/NET33_XI18/XI7/MM2_g
+ N_VSS_XI18/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM3 N_XI18/XI7/NET33_XI18/XI7/MM3_d N_WL<32>_XI18/XI7/MM3_g
+ N_BLN<8>_XI18/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM0 N_XI18/XI7/NET34_XI18/XI7/MM0_d N_WL<32>_XI18/XI7/MM0_g
+ N_BL<8>_XI18/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM1 N_XI18/XI7/NET33_XI18/XI7/MM1_d N_XI18/XI7/NET34_XI18/XI7/MM1_g
+ N_VSS_XI18/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM9 N_XI18/XI7/NET36_XI18/XI7/MM9_d N_WL<33>_XI18/XI7/MM9_g
+ N_BL<8>_XI18/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM6 N_XI18/XI7/NET35_XI18/XI7/MM6_d N_XI18/XI7/NET36_XI18/XI7/MM6_g
+ N_VSS_XI18/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM7 N_XI18/XI7/NET36_XI18/XI7/MM7_d N_XI18/XI7/NET35_XI18/XI7/MM7_g
+ N_VSS_XI18/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM8 N_XI18/XI7/NET35_XI18/XI7/MM8_d N_WL<33>_XI18/XI7/MM8_g
+ N_BLN<8>_XI18/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI7/MM5 N_XI18/XI7/NET34_XI18/XI7/MM5_d N_XI18/XI7/NET33_XI18/XI7/MM5_g
+ N_VDD_XI18/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI7/MM4 N_XI18/XI7/NET33_XI18/XI7/MM4_d N_XI18/XI7/NET34_XI18/XI7/MM4_g
+ N_VDD_XI18/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI7/MM10 N_XI18/XI7/NET35_XI18/XI7/MM10_d N_XI18/XI7/NET36_XI18/XI7/MM10_g
+ N_VDD_XI18/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI7/MM11 N_XI18/XI7/NET36_XI18/XI7/MM11_d N_XI18/XI7/NET35_XI18/XI7/MM11_g
+ N_VDD_XI18/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI8/MM2 N_XI18/XI8/NET34_XI18/XI8/MM2_d N_XI18/XI8/NET33_XI18/XI8/MM2_g
+ N_VSS_XI18/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM3 N_XI18/XI8/NET33_XI18/XI8/MM3_d N_WL<32>_XI18/XI8/MM3_g
+ N_BLN<7>_XI18/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM0 N_XI18/XI8/NET34_XI18/XI8/MM0_d N_WL<32>_XI18/XI8/MM0_g
+ N_BL<7>_XI18/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM1 N_XI18/XI8/NET33_XI18/XI8/MM1_d N_XI18/XI8/NET34_XI18/XI8/MM1_g
+ N_VSS_XI18/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM9 N_XI18/XI8/NET36_XI18/XI8/MM9_d N_WL<33>_XI18/XI8/MM9_g
+ N_BL<7>_XI18/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM6 N_XI18/XI8/NET35_XI18/XI8/MM6_d N_XI18/XI8/NET36_XI18/XI8/MM6_g
+ N_VSS_XI18/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM7 N_XI18/XI8/NET36_XI18/XI8/MM7_d N_XI18/XI8/NET35_XI18/XI8/MM7_g
+ N_VSS_XI18/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM8 N_XI18/XI8/NET35_XI18/XI8/MM8_d N_WL<33>_XI18/XI8/MM8_g
+ N_BLN<7>_XI18/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI8/MM5 N_XI18/XI8/NET34_XI18/XI8/MM5_d N_XI18/XI8/NET33_XI18/XI8/MM5_g
+ N_VDD_XI18/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI8/MM4 N_XI18/XI8/NET33_XI18/XI8/MM4_d N_XI18/XI8/NET34_XI18/XI8/MM4_g
+ N_VDD_XI18/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI8/MM10 N_XI18/XI8/NET35_XI18/XI8/MM10_d N_XI18/XI8/NET36_XI18/XI8/MM10_g
+ N_VDD_XI18/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI8/MM11 N_XI18/XI8/NET36_XI18/XI8/MM11_d N_XI18/XI8/NET35_XI18/XI8/MM11_g
+ N_VDD_XI18/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI9/MM2 N_XI18/XI9/NET34_XI18/XI9/MM2_d N_XI18/XI9/NET33_XI18/XI9/MM2_g
+ N_VSS_XI18/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM3 N_XI18/XI9/NET33_XI18/XI9/MM3_d N_WL<32>_XI18/XI9/MM3_g
+ N_BLN<6>_XI18/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM0 N_XI18/XI9/NET34_XI18/XI9/MM0_d N_WL<32>_XI18/XI9/MM0_g
+ N_BL<6>_XI18/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM1 N_XI18/XI9/NET33_XI18/XI9/MM1_d N_XI18/XI9/NET34_XI18/XI9/MM1_g
+ N_VSS_XI18/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM9 N_XI18/XI9/NET36_XI18/XI9/MM9_d N_WL<33>_XI18/XI9/MM9_g
+ N_BL<6>_XI18/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM6 N_XI18/XI9/NET35_XI18/XI9/MM6_d N_XI18/XI9/NET36_XI18/XI9/MM6_g
+ N_VSS_XI18/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM7 N_XI18/XI9/NET36_XI18/XI9/MM7_d N_XI18/XI9/NET35_XI18/XI9/MM7_g
+ N_VSS_XI18/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM8 N_XI18/XI9/NET35_XI18/XI9/MM8_d N_WL<33>_XI18/XI9/MM8_g
+ N_BLN<6>_XI18/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI9/MM5 N_XI18/XI9/NET34_XI18/XI9/MM5_d N_XI18/XI9/NET33_XI18/XI9/MM5_g
+ N_VDD_XI18/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI9/MM4 N_XI18/XI9/NET33_XI18/XI9/MM4_d N_XI18/XI9/NET34_XI18/XI9/MM4_g
+ N_VDD_XI18/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI9/MM10 N_XI18/XI9/NET35_XI18/XI9/MM10_d N_XI18/XI9/NET36_XI18/XI9/MM10_g
+ N_VDD_XI18/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI9/MM11 N_XI18/XI9/NET36_XI18/XI9/MM11_d N_XI18/XI9/NET35_XI18/XI9/MM11_g
+ N_VDD_XI18/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI10/MM2 N_XI18/XI10/NET34_XI18/XI10/MM2_d
+ N_XI18/XI10/NET33_XI18/XI10/MM2_g N_VSS_XI18/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI10/MM3 N_XI18/XI10/NET33_XI18/XI10/MM3_d N_WL<32>_XI18/XI10/MM3_g
+ N_BLN<5>_XI18/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI10/MM0 N_XI18/XI10/NET34_XI18/XI10/MM0_d N_WL<32>_XI18/XI10/MM0_g
+ N_BL<5>_XI18/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI10/MM1 N_XI18/XI10/NET33_XI18/XI10/MM1_d
+ N_XI18/XI10/NET34_XI18/XI10/MM1_g N_VSS_XI18/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI10/MM9 N_XI18/XI10/NET36_XI18/XI10/MM9_d N_WL<33>_XI18/XI10/MM9_g
+ N_BL<5>_XI18/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI10/MM6 N_XI18/XI10/NET35_XI18/XI10/MM6_d
+ N_XI18/XI10/NET36_XI18/XI10/MM6_g N_VSS_XI18/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI10/MM7 N_XI18/XI10/NET36_XI18/XI10/MM7_d
+ N_XI18/XI10/NET35_XI18/XI10/MM7_g N_VSS_XI18/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI10/MM8 N_XI18/XI10/NET35_XI18/XI10/MM8_d N_WL<33>_XI18/XI10/MM8_g
+ N_BLN<5>_XI18/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI10/MM5 N_XI18/XI10/NET34_XI18/XI10/MM5_d
+ N_XI18/XI10/NET33_XI18/XI10/MM5_g N_VDD_XI18/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI10/MM4 N_XI18/XI10/NET33_XI18/XI10/MM4_d
+ N_XI18/XI10/NET34_XI18/XI10/MM4_g N_VDD_XI18/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI10/MM10 N_XI18/XI10/NET35_XI18/XI10/MM10_d
+ N_XI18/XI10/NET36_XI18/XI10/MM10_g N_VDD_XI18/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI10/MM11 N_XI18/XI10/NET36_XI18/XI10/MM11_d
+ N_XI18/XI10/NET35_XI18/XI10/MM11_g N_VDD_XI18/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI11/MM2 N_XI18/XI11/NET34_XI18/XI11/MM2_d
+ N_XI18/XI11/NET33_XI18/XI11/MM2_g N_VSS_XI18/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI11/MM3 N_XI18/XI11/NET33_XI18/XI11/MM3_d N_WL<32>_XI18/XI11/MM3_g
+ N_BLN<4>_XI18/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI11/MM0 N_XI18/XI11/NET34_XI18/XI11/MM0_d N_WL<32>_XI18/XI11/MM0_g
+ N_BL<4>_XI18/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI11/MM1 N_XI18/XI11/NET33_XI18/XI11/MM1_d
+ N_XI18/XI11/NET34_XI18/XI11/MM1_g N_VSS_XI18/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI11/MM9 N_XI18/XI11/NET36_XI18/XI11/MM9_d N_WL<33>_XI18/XI11/MM9_g
+ N_BL<4>_XI18/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI11/MM6 N_XI18/XI11/NET35_XI18/XI11/MM6_d
+ N_XI18/XI11/NET36_XI18/XI11/MM6_g N_VSS_XI18/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI11/MM7 N_XI18/XI11/NET36_XI18/XI11/MM7_d
+ N_XI18/XI11/NET35_XI18/XI11/MM7_g N_VSS_XI18/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI11/MM8 N_XI18/XI11/NET35_XI18/XI11/MM8_d N_WL<33>_XI18/XI11/MM8_g
+ N_BLN<4>_XI18/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI11/MM5 N_XI18/XI11/NET34_XI18/XI11/MM5_d
+ N_XI18/XI11/NET33_XI18/XI11/MM5_g N_VDD_XI18/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI11/MM4 N_XI18/XI11/NET33_XI18/XI11/MM4_d
+ N_XI18/XI11/NET34_XI18/XI11/MM4_g N_VDD_XI18/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI11/MM10 N_XI18/XI11/NET35_XI18/XI11/MM10_d
+ N_XI18/XI11/NET36_XI18/XI11/MM10_g N_VDD_XI18/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI11/MM11 N_XI18/XI11/NET36_XI18/XI11/MM11_d
+ N_XI18/XI11/NET35_XI18/XI11/MM11_g N_VDD_XI18/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI12/MM2 N_XI18/XI12/NET34_XI18/XI12/MM2_d
+ N_XI18/XI12/NET33_XI18/XI12/MM2_g N_VSS_XI18/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI12/MM3 N_XI18/XI12/NET33_XI18/XI12/MM3_d N_WL<32>_XI18/XI12/MM3_g
+ N_BLN<3>_XI18/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI12/MM0 N_XI18/XI12/NET34_XI18/XI12/MM0_d N_WL<32>_XI18/XI12/MM0_g
+ N_BL<3>_XI18/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI12/MM1 N_XI18/XI12/NET33_XI18/XI12/MM1_d
+ N_XI18/XI12/NET34_XI18/XI12/MM1_g N_VSS_XI18/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI12/MM9 N_XI18/XI12/NET36_XI18/XI12/MM9_d N_WL<33>_XI18/XI12/MM9_g
+ N_BL<3>_XI18/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI12/MM6 N_XI18/XI12/NET35_XI18/XI12/MM6_d
+ N_XI18/XI12/NET36_XI18/XI12/MM6_g N_VSS_XI18/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI12/MM7 N_XI18/XI12/NET36_XI18/XI12/MM7_d
+ N_XI18/XI12/NET35_XI18/XI12/MM7_g N_VSS_XI18/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI12/MM8 N_XI18/XI12/NET35_XI18/XI12/MM8_d N_WL<33>_XI18/XI12/MM8_g
+ N_BLN<3>_XI18/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI12/MM5 N_XI18/XI12/NET34_XI18/XI12/MM5_d
+ N_XI18/XI12/NET33_XI18/XI12/MM5_g N_VDD_XI18/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI12/MM4 N_XI18/XI12/NET33_XI18/XI12/MM4_d
+ N_XI18/XI12/NET34_XI18/XI12/MM4_g N_VDD_XI18/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI12/MM10 N_XI18/XI12/NET35_XI18/XI12/MM10_d
+ N_XI18/XI12/NET36_XI18/XI12/MM10_g N_VDD_XI18/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI12/MM11 N_XI18/XI12/NET36_XI18/XI12/MM11_d
+ N_XI18/XI12/NET35_XI18/XI12/MM11_g N_VDD_XI18/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI13/MM2 N_XI18/XI13/NET34_XI18/XI13/MM2_d
+ N_XI18/XI13/NET33_XI18/XI13/MM2_g N_VSS_XI18/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI13/MM3 N_XI18/XI13/NET33_XI18/XI13/MM3_d N_WL<32>_XI18/XI13/MM3_g
+ N_BLN<2>_XI18/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI13/MM0 N_XI18/XI13/NET34_XI18/XI13/MM0_d N_WL<32>_XI18/XI13/MM0_g
+ N_BL<2>_XI18/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI13/MM1 N_XI18/XI13/NET33_XI18/XI13/MM1_d
+ N_XI18/XI13/NET34_XI18/XI13/MM1_g N_VSS_XI18/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI13/MM9 N_XI18/XI13/NET36_XI18/XI13/MM9_d N_WL<33>_XI18/XI13/MM9_g
+ N_BL<2>_XI18/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI13/MM6 N_XI18/XI13/NET35_XI18/XI13/MM6_d
+ N_XI18/XI13/NET36_XI18/XI13/MM6_g N_VSS_XI18/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI13/MM7 N_XI18/XI13/NET36_XI18/XI13/MM7_d
+ N_XI18/XI13/NET35_XI18/XI13/MM7_g N_VSS_XI18/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI13/MM8 N_XI18/XI13/NET35_XI18/XI13/MM8_d N_WL<33>_XI18/XI13/MM8_g
+ N_BLN<2>_XI18/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI13/MM5 N_XI18/XI13/NET34_XI18/XI13/MM5_d
+ N_XI18/XI13/NET33_XI18/XI13/MM5_g N_VDD_XI18/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI13/MM4 N_XI18/XI13/NET33_XI18/XI13/MM4_d
+ N_XI18/XI13/NET34_XI18/XI13/MM4_g N_VDD_XI18/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI13/MM10 N_XI18/XI13/NET35_XI18/XI13/MM10_d
+ N_XI18/XI13/NET36_XI18/XI13/MM10_g N_VDD_XI18/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI13/MM11 N_XI18/XI13/NET36_XI18/XI13/MM11_d
+ N_XI18/XI13/NET35_XI18/XI13/MM11_g N_VDD_XI18/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI14/MM2 N_XI18/XI14/NET34_XI18/XI14/MM2_d
+ N_XI18/XI14/NET33_XI18/XI14/MM2_g N_VSS_XI18/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI14/MM3 N_XI18/XI14/NET33_XI18/XI14/MM3_d N_WL<32>_XI18/XI14/MM3_g
+ N_BLN<1>_XI18/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI14/MM0 N_XI18/XI14/NET34_XI18/XI14/MM0_d N_WL<32>_XI18/XI14/MM0_g
+ N_BL<1>_XI18/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI14/MM1 N_XI18/XI14/NET33_XI18/XI14/MM1_d
+ N_XI18/XI14/NET34_XI18/XI14/MM1_g N_VSS_XI18/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI14/MM9 N_XI18/XI14/NET36_XI18/XI14/MM9_d N_WL<33>_XI18/XI14/MM9_g
+ N_BL<1>_XI18/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI14/MM6 N_XI18/XI14/NET35_XI18/XI14/MM6_d
+ N_XI18/XI14/NET36_XI18/XI14/MM6_g N_VSS_XI18/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI14/MM7 N_XI18/XI14/NET36_XI18/XI14/MM7_d
+ N_XI18/XI14/NET35_XI18/XI14/MM7_g N_VSS_XI18/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI14/MM8 N_XI18/XI14/NET35_XI18/XI14/MM8_d N_WL<33>_XI18/XI14/MM8_g
+ N_BLN<1>_XI18/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI14/MM5 N_XI18/XI14/NET34_XI18/XI14/MM5_d
+ N_XI18/XI14/NET33_XI18/XI14/MM5_g N_VDD_XI18/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI14/MM4 N_XI18/XI14/NET33_XI18/XI14/MM4_d
+ N_XI18/XI14/NET34_XI18/XI14/MM4_g N_VDD_XI18/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI14/MM10 N_XI18/XI14/NET35_XI18/XI14/MM10_d
+ N_XI18/XI14/NET36_XI18/XI14/MM10_g N_VDD_XI18/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI14/MM11 N_XI18/XI14/NET36_XI18/XI14/MM11_d
+ N_XI18/XI14/NET35_XI18/XI14/MM11_g N_VDD_XI18/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI15/MM2 N_XI18/XI15/NET34_XI18/XI15/MM2_d
+ N_XI18/XI15/NET33_XI18/XI15/MM2_g N_VSS_XI18/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI15/MM3 N_XI18/XI15/NET33_XI18/XI15/MM3_d N_WL<32>_XI18/XI15/MM3_g
+ N_BLN<0>_XI18/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI15/MM0 N_XI18/XI15/NET34_XI18/XI15/MM0_d N_WL<32>_XI18/XI15/MM0_g
+ N_BL<0>_XI18/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI15/MM1 N_XI18/XI15/NET33_XI18/XI15/MM1_d
+ N_XI18/XI15/NET34_XI18/XI15/MM1_g N_VSS_XI18/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI15/MM9 N_XI18/XI15/NET36_XI18/XI15/MM9_d N_WL<33>_XI18/XI15/MM9_g
+ N_BL<0>_XI18/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI15/MM6 N_XI18/XI15/NET35_XI18/XI15/MM6_d
+ N_XI18/XI15/NET36_XI18/XI15/MM6_g N_VSS_XI18/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI15/MM7 N_XI18/XI15/NET36_XI18/XI15/MM7_d
+ N_XI18/XI15/NET35_XI18/XI15/MM7_g N_VSS_XI18/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI18/XI15/MM8 N_XI18/XI15/NET35_XI18/XI15/MM8_d N_WL<33>_XI18/XI15/MM8_g
+ N_BLN<0>_XI18/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI18/XI15/MM5 N_XI18/XI15/NET34_XI18/XI15/MM5_d
+ N_XI18/XI15/NET33_XI18/XI15/MM5_g N_VDD_XI18/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI15/MM4 N_XI18/XI15/NET33_XI18/XI15/MM4_d
+ N_XI18/XI15/NET34_XI18/XI15/MM4_g N_VDD_XI18/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI15/MM10 N_XI18/XI15/NET35_XI18/XI15/MM10_d
+ N_XI18/XI15/NET36_XI18/XI15/MM10_g N_VDD_XI18/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI18/XI15/MM11 N_XI18/XI15/NET36_XI18/XI15/MM11_d
+ N_XI18/XI15/NET35_XI18/XI15/MM11_g N_VDD_XI18/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI0/MM2 N_XI19/XI0/NET34_XI19/XI0/MM2_d N_XI19/XI0/NET33_XI19/XI0/MM2_g
+ N_VSS_XI19/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI0/MM3 N_XI19/XI0/NET33_XI19/XI0/MM3_d N_WL<34>_XI19/XI0/MM3_g
+ N_BLN<15>_XI19/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI0/MM0 N_XI19/XI0/NET34_XI19/XI0/MM0_d N_WL<34>_XI19/XI0/MM0_g
+ N_BL<15>_XI19/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI0/MM1 N_XI19/XI0/NET33_XI19/XI0/MM1_d N_XI19/XI0/NET34_XI19/XI0/MM1_g
+ N_VSS_XI19/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI0/MM9 N_XI19/XI0/NET36_XI19/XI0/MM9_d N_WL<35>_XI19/XI0/MM9_g
+ N_BL<15>_XI19/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI0/MM6 N_XI19/XI0/NET35_XI19/XI0/MM6_d N_XI19/XI0/NET36_XI19/XI0/MM6_g
+ N_VSS_XI19/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI0/MM7 N_XI19/XI0/NET36_XI19/XI0/MM7_d N_XI19/XI0/NET35_XI19/XI0/MM7_g
+ N_VSS_XI19/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI0/MM8 N_XI19/XI0/NET35_XI19/XI0/MM8_d N_WL<35>_XI19/XI0/MM8_g
+ N_BLN<15>_XI19/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI0/MM5 N_XI19/XI0/NET34_XI19/XI0/MM5_d N_XI19/XI0/NET33_XI19/XI0/MM5_g
+ N_VDD_XI19/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI0/MM4 N_XI19/XI0/NET33_XI19/XI0/MM4_d N_XI19/XI0/NET34_XI19/XI0/MM4_g
+ N_VDD_XI19/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI0/MM10 N_XI19/XI0/NET35_XI19/XI0/MM10_d N_XI19/XI0/NET36_XI19/XI0/MM10_g
+ N_VDD_XI19/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI0/MM11 N_XI19/XI0/NET36_XI19/XI0/MM11_d N_XI19/XI0/NET35_XI19/XI0/MM11_g
+ N_VDD_XI19/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI1/MM2 N_XI19/XI1/NET34_XI19/XI1/MM2_d N_XI19/XI1/NET33_XI19/XI1/MM2_g
+ N_VSS_XI19/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI1/MM3 N_XI19/XI1/NET33_XI19/XI1/MM3_d N_WL<34>_XI19/XI1/MM3_g
+ N_BLN<14>_XI19/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI1/MM0 N_XI19/XI1/NET34_XI19/XI1/MM0_d N_WL<34>_XI19/XI1/MM0_g
+ N_BL<14>_XI19/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI1/MM1 N_XI19/XI1/NET33_XI19/XI1/MM1_d N_XI19/XI1/NET34_XI19/XI1/MM1_g
+ N_VSS_XI19/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI1/MM9 N_XI19/XI1/NET36_XI19/XI1/MM9_d N_WL<35>_XI19/XI1/MM9_g
+ N_BL<14>_XI19/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI1/MM6 N_XI19/XI1/NET35_XI19/XI1/MM6_d N_XI19/XI1/NET36_XI19/XI1/MM6_g
+ N_VSS_XI19/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI1/MM7 N_XI19/XI1/NET36_XI19/XI1/MM7_d N_XI19/XI1/NET35_XI19/XI1/MM7_g
+ N_VSS_XI19/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI1/MM8 N_XI19/XI1/NET35_XI19/XI1/MM8_d N_WL<35>_XI19/XI1/MM8_g
+ N_BLN<14>_XI19/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI1/MM5 N_XI19/XI1/NET34_XI19/XI1/MM5_d N_XI19/XI1/NET33_XI19/XI1/MM5_g
+ N_VDD_XI19/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI1/MM4 N_XI19/XI1/NET33_XI19/XI1/MM4_d N_XI19/XI1/NET34_XI19/XI1/MM4_g
+ N_VDD_XI19/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI1/MM10 N_XI19/XI1/NET35_XI19/XI1/MM10_d N_XI19/XI1/NET36_XI19/XI1/MM10_g
+ N_VDD_XI19/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI1/MM11 N_XI19/XI1/NET36_XI19/XI1/MM11_d N_XI19/XI1/NET35_XI19/XI1/MM11_g
+ N_VDD_XI19/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI2/MM2 N_XI19/XI2/NET34_XI19/XI2/MM2_d N_XI19/XI2/NET33_XI19/XI2/MM2_g
+ N_VSS_XI19/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI2/MM3 N_XI19/XI2/NET33_XI19/XI2/MM3_d N_WL<34>_XI19/XI2/MM3_g
+ N_BLN<13>_XI19/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI2/MM0 N_XI19/XI2/NET34_XI19/XI2/MM0_d N_WL<34>_XI19/XI2/MM0_g
+ N_BL<13>_XI19/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI2/MM1 N_XI19/XI2/NET33_XI19/XI2/MM1_d N_XI19/XI2/NET34_XI19/XI2/MM1_g
+ N_VSS_XI19/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI2/MM9 N_XI19/XI2/NET36_XI19/XI2/MM9_d N_WL<35>_XI19/XI2/MM9_g
+ N_BL<13>_XI19/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI2/MM6 N_XI19/XI2/NET35_XI19/XI2/MM6_d N_XI19/XI2/NET36_XI19/XI2/MM6_g
+ N_VSS_XI19/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI2/MM7 N_XI19/XI2/NET36_XI19/XI2/MM7_d N_XI19/XI2/NET35_XI19/XI2/MM7_g
+ N_VSS_XI19/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI2/MM8 N_XI19/XI2/NET35_XI19/XI2/MM8_d N_WL<35>_XI19/XI2/MM8_g
+ N_BLN<13>_XI19/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI2/MM5 N_XI19/XI2/NET34_XI19/XI2/MM5_d N_XI19/XI2/NET33_XI19/XI2/MM5_g
+ N_VDD_XI19/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI2/MM4 N_XI19/XI2/NET33_XI19/XI2/MM4_d N_XI19/XI2/NET34_XI19/XI2/MM4_g
+ N_VDD_XI19/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI2/MM10 N_XI19/XI2/NET35_XI19/XI2/MM10_d N_XI19/XI2/NET36_XI19/XI2/MM10_g
+ N_VDD_XI19/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI2/MM11 N_XI19/XI2/NET36_XI19/XI2/MM11_d N_XI19/XI2/NET35_XI19/XI2/MM11_g
+ N_VDD_XI19/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI3/MM2 N_XI19/XI3/NET34_XI19/XI3/MM2_d N_XI19/XI3/NET33_XI19/XI3/MM2_g
+ N_VSS_XI19/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI3/MM3 N_XI19/XI3/NET33_XI19/XI3/MM3_d N_WL<34>_XI19/XI3/MM3_g
+ N_BLN<12>_XI19/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI3/MM0 N_XI19/XI3/NET34_XI19/XI3/MM0_d N_WL<34>_XI19/XI3/MM0_g
+ N_BL<12>_XI19/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI3/MM1 N_XI19/XI3/NET33_XI19/XI3/MM1_d N_XI19/XI3/NET34_XI19/XI3/MM1_g
+ N_VSS_XI19/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI3/MM9 N_XI19/XI3/NET36_XI19/XI3/MM9_d N_WL<35>_XI19/XI3/MM9_g
+ N_BL<12>_XI19/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI3/MM6 N_XI19/XI3/NET35_XI19/XI3/MM6_d N_XI19/XI3/NET36_XI19/XI3/MM6_g
+ N_VSS_XI19/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI3/MM7 N_XI19/XI3/NET36_XI19/XI3/MM7_d N_XI19/XI3/NET35_XI19/XI3/MM7_g
+ N_VSS_XI19/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI3/MM8 N_XI19/XI3/NET35_XI19/XI3/MM8_d N_WL<35>_XI19/XI3/MM8_g
+ N_BLN<12>_XI19/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI3/MM5 N_XI19/XI3/NET34_XI19/XI3/MM5_d N_XI19/XI3/NET33_XI19/XI3/MM5_g
+ N_VDD_XI19/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI3/MM4 N_XI19/XI3/NET33_XI19/XI3/MM4_d N_XI19/XI3/NET34_XI19/XI3/MM4_g
+ N_VDD_XI19/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI3/MM10 N_XI19/XI3/NET35_XI19/XI3/MM10_d N_XI19/XI3/NET36_XI19/XI3/MM10_g
+ N_VDD_XI19/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI3/MM11 N_XI19/XI3/NET36_XI19/XI3/MM11_d N_XI19/XI3/NET35_XI19/XI3/MM11_g
+ N_VDD_XI19/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI4/MM2 N_XI19/XI4/NET34_XI19/XI4/MM2_d N_XI19/XI4/NET33_XI19/XI4/MM2_g
+ N_VSS_XI19/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI4/MM3 N_XI19/XI4/NET33_XI19/XI4/MM3_d N_WL<34>_XI19/XI4/MM3_g
+ N_BLN<11>_XI19/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI4/MM0 N_XI19/XI4/NET34_XI19/XI4/MM0_d N_WL<34>_XI19/XI4/MM0_g
+ N_BL<11>_XI19/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI4/MM1 N_XI19/XI4/NET33_XI19/XI4/MM1_d N_XI19/XI4/NET34_XI19/XI4/MM1_g
+ N_VSS_XI19/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI4/MM9 N_XI19/XI4/NET36_XI19/XI4/MM9_d N_WL<35>_XI19/XI4/MM9_g
+ N_BL<11>_XI19/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI4/MM6 N_XI19/XI4/NET35_XI19/XI4/MM6_d N_XI19/XI4/NET36_XI19/XI4/MM6_g
+ N_VSS_XI19/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI4/MM7 N_XI19/XI4/NET36_XI19/XI4/MM7_d N_XI19/XI4/NET35_XI19/XI4/MM7_g
+ N_VSS_XI19/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI4/MM8 N_XI19/XI4/NET35_XI19/XI4/MM8_d N_WL<35>_XI19/XI4/MM8_g
+ N_BLN<11>_XI19/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI4/MM5 N_XI19/XI4/NET34_XI19/XI4/MM5_d N_XI19/XI4/NET33_XI19/XI4/MM5_g
+ N_VDD_XI19/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI4/MM4 N_XI19/XI4/NET33_XI19/XI4/MM4_d N_XI19/XI4/NET34_XI19/XI4/MM4_g
+ N_VDD_XI19/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI4/MM10 N_XI19/XI4/NET35_XI19/XI4/MM10_d N_XI19/XI4/NET36_XI19/XI4/MM10_g
+ N_VDD_XI19/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI4/MM11 N_XI19/XI4/NET36_XI19/XI4/MM11_d N_XI19/XI4/NET35_XI19/XI4/MM11_g
+ N_VDD_XI19/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI5/MM2 N_XI19/XI5/NET34_XI19/XI5/MM2_d N_XI19/XI5/NET33_XI19/XI5/MM2_g
+ N_VSS_XI19/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI5/MM3 N_XI19/XI5/NET33_XI19/XI5/MM3_d N_WL<34>_XI19/XI5/MM3_g
+ N_BLN<10>_XI19/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI5/MM0 N_XI19/XI5/NET34_XI19/XI5/MM0_d N_WL<34>_XI19/XI5/MM0_g
+ N_BL<10>_XI19/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI5/MM1 N_XI19/XI5/NET33_XI19/XI5/MM1_d N_XI19/XI5/NET34_XI19/XI5/MM1_g
+ N_VSS_XI19/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI5/MM9 N_XI19/XI5/NET36_XI19/XI5/MM9_d N_WL<35>_XI19/XI5/MM9_g
+ N_BL<10>_XI19/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI5/MM6 N_XI19/XI5/NET35_XI19/XI5/MM6_d N_XI19/XI5/NET36_XI19/XI5/MM6_g
+ N_VSS_XI19/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI5/MM7 N_XI19/XI5/NET36_XI19/XI5/MM7_d N_XI19/XI5/NET35_XI19/XI5/MM7_g
+ N_VSS_XI19/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI5/MM8 N_XI19/XI5/NET35_XI19/XI5/MM8_d N_WL<35>_XI19/XI5/MM8_g
+ N_BLN<10>_XI19/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI5/MM5 N_XI19/XI5/NET34_XI19/XI5/MM5_d N_XI19/XI5/NET33_XI19/XI5/MM5_g
+ N_VDD_XI19/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI5/MM4 N_XI19/XI5/NET33_XI19/XI5/MM4_d N_XI19/XI5/NET34_XI19/XI5/MM4_g
+ N_VDD_XI19/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI5/MM10 N_XI19/XI5/NET35_XI19/XI5/MM10_d N_XI19/XI5/NET36_XI19/XI5/MM10_g
+ N_VDD_XI19/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI5/MM11 N_XI19/XI5/NET36_XI19/XI5/MM11_d N_XI19/XI5/NET35_XI19/XI5/MM11_g
+ N_VDD_XI19/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI6/MM2 N_XI19/XI6/NET34_XI19/XI6/MM2_d N_XI19/XI6/NET33_XI19/XI6/MM2_g
+ N_VSS_XI19/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM3 N_XI19/XI6/NET33_XI19/XI6/MM3_d N_WL<34>_XI19/XI6/MM3_g
+ N_BLN<9>_XI19/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM0 N_XI19/XI6/NET34_XI19/XI6/MM0_d N_WL<34>_XI19/XI6/MM0_g
+ N_BL<9>_XI19/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM1 N_XI19/XI6/NET33_XI19/XI6/MM1_d N_XI19/XI6/NET34_XI19/XI6/MM1_g
+ N_VSS_XI19/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM9 N_XI19/XI6/NET36_XI19/XI6/MM9_d N_WL<35>_XI19/XI6/MM9_g
+ N_BL<9>_XI19/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM6 N_XI19/XI6/NET35_XI19/XI6/MM6_d N_XI19/XI6/NET36_XI19/XI6/MM6_g
+ N_VSS_XI19/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM7 N_XI19/XI6/NET36_XI19/XI6/MM7_d N_XI19/XI6/NET35_XI19/XI6/MM7_g
+ N_VSS_XI19/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM8 N_XI19/XI6/NET35_XI19/XI6/MM8_d N_WL<35>_XI19/XI6/MM8_g
+ N_BLN<9>_XI19/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI6/MM5 N_XI19/XI6/NET34_XI19/XI6/MM5_d N_XI19/XI6/NET33_XI19/XI6/MM5_g
+ N_VDD_XI19/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI6/MM4 N_XI19/XI6/NET33_XI19/XI6/MM4_d N_XI19/XI6/NET34_XI19/XI6/MM4_g
+ N_VDD_XI19/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI6/MM10 N_XI19/XI6/NET35_XI19/XI6/MM10_d N_XI19/XI6/NET36_XI19/XI6/MM10_g
+ N_VDD_XI19/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI6/MM11 N_XI19/XI6/NET36_XI19/XI6/MM11_d N_XI19/XI6/NET35_XI19/XI6/MM11_g
+ N_VDD_XI19/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI7/MM2 N_XI19/XI7/NET34_XI19/XI7/MM2_d N_XI19/XI7/NET33_XI19/XI7/MM2_g
+ N_VSS_XI19/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM3 N_XI19/XI7/NET33_XI19/XI7/MM3_d N_WL<34>_XI19/XI7/MM3_g
+ N_BLN<8>_XI19/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM0 N_XI19/XI7/NET34_XI19/XI7/MM0_d N_WL<34>_XI19/XI7/MM0_g
+ N_BL<8>_XI19/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM1 N_XI19/XI7/NET33_XI19/XI7/MM1_d N_XI19/XI7/NET34_XI19/XI7/MM1_g
+ N_VSS_XI19/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM9 N_XI19/XI7/NET36_XI19/XI7/MM9_d N_WL<35>_XI19/XI7/MM9_g
+ N_BL<8>_XI19/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM6 N_XI19/XI7/NET35_XI19/XI7/MM6_d N_XI19/XI7/NET36_XI19/XI7/MM6_g
+ N_VSS_XI19/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM7 N_XI19/XI7/NET36_XI19/XI7/MM7_d N_XI19/XI7/NET35_XI19/XI7/MM7_g
+ N_VSS_XI19/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM8 N_XI19/XI7/NET35_XI19/XI7/MM8_d N_WL<35>_XI19/XI7/MM8_g
+ N_BLN<8>_XI19/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI7/MM5 N_XI19/XI7/NET34_XI19/XI7/MM5_d N_XI19/XI7/NET33_XI19/XI7/MM5_g
+ N_VDD_XI19/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI7/MM4 N_XI19/XI7/NET33_XI19/XI7/MM4_d N_XI19/XI7/NET34_XI19/XI7/MM4_g
+ N_VDD_XI19/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI7/MM10 N_XI19/XI7/NET35_XI19/XI7/MM10_d N_XI19/XI7/NET36_XI19/XI7/MM10_g
+ N_VDD_XI19/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI7/MM11 N_XI19/XI7/NET36_XI19/XI7/MM11_d N_XI19/XI7/NET35_XI19/XI7/MM11_g
+ N_VDD_XI19/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI8/MM2 N_XI19/XI8/NET34_XI19/XI8/MM2_d N_XI19/XI8/NET33_XI19/XI8/MM2_g
+ N_VSS_XI19/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM3 N_XI19/XI8/NET33_XI19/XI8/MM3_d N_WL<34>_XI19/XI8/MM3_g
+ N_BLN<7>_XI19/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM0 N_XI19/XI8/NET34_XI19/XI8/MM0_d N_WL<34>_XI19/XI8/MM0_g
+ N_BL<7>_XI19/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM1 N_XI19/XI8/NET33_XI19/XI8/MM1_d N_XI19/XI8/NET34_XI19/XI8/MM1_g
+ N_VSS_XI19/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM9 N_XI19/XI8/NET36_XI19/XI8/MM9_d N_WL<35>_XI19/XI8/MM9_g
+ N_BL<7>_XI19/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM6 N_XI19/XI8/NET35_XI19/XI8/MM6_d N_XI19/XI8/NET36_XI19/XI8/MM6_g
+ N_VSS_XI19/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM7 N_XI19/XI8/NET36_XI19/XI8/MM7_d N_XI19/XI8/NET35_XI19/XI8/MM7_g
+ N_VSS_XI19/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM8 N_XI19/XI8/NET35_XI19/XI8/MM8_d N_WL<35>_XI19/XI8/MM8_g
+ N_BLN<7>_XI19/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI8/MM5 N_XI19/XI8/NET34_XI19/XI8/MM5_d N_XI19/XI8/NET33_XI19/XI8/MM5_g
+ N_VDD_XI19/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI8/MM4 N_XI19/XI8/NET33_XI19/XI8/MM4_d N_XI19/XI8/NET34_XI19/XI8/MM4_g
+ N_VDD_XI19/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI8/MM10 N_XI19/XI8/NET35_XI19/XI8/MM10_d N_XI19/XI8/NET36_XI19/XI8/MM10_g
+ N_VDD_XI19/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI8/MM11 N_XI19/XI8/NET36_XI19/XI8/MM11_d N_XI19/XI8/NET35_XI19/XI8/MM11_g
+ N_VDD_XI19/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI9/MM2 N_XI19/XI9/NET34_XI19/XI9/MM2_d N_XI19/XI9/NET33_XI19/XI9/MM2_g
+ N_VSS_XI19/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM3 N_XI19/XI9/NET33_XI19/XI9/MM3_d N_WL<34>_XI19/XI9/MM3_g
+ N_BLN<6>_XI19/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM0 N_XI19/XI9/NET34_XI19/XI9/MM0_d N_WL<34>_XI19/XI9/MM0_g
+ N_BL<6>_XI19/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM1 N_XI19/XI9/NET33_XI19/XI9/MM1_d N_XI19/XI9/NET34_XI19/XI9/MM1_g
+ N_VSS_XI19/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM9 N_XI19/XI9/NET36_XI19/XI9/MM9_d N_WL<35>_XI19/XI9/MM9_g
+ N_BL<6>_XI19/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM6 N_XI19/XI9/NET35_XI19/XI9/MM6_d N_XI19/XI9/NET36_XI19/XI9/MM6_g
+ N_VSS_XI19/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM7 N_XI19/XI9/NET36_XI19/XI9/MM7_d N_XI19/XI9/NET35_XI19/XI9/MM7_g
+ N_VSS_XI19/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM8 N_XI19/XI9/NET35_XI19/XI9/MM8_d N_WL<35>_XI19/XI9/MM8_g
+ N_BLN<6>_XI19/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI9/MM5 N_XI19/XI9/NET34_XI19/XI9/MM5_d N_XI19/XI9/NET33_XI19/XI9/MM5_g
+ N_VDD_XI19/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI9/MM4 N_XI19/XI9/NET33_XI19/XI9/MM4_d N_XI19/XI9/NET34_XI19/XI9/MM4_g
+ N_VDD_XI19/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI9/MM10 N_XI19/XI9/NET35_XI19/XI9/MM10_d N_XI19/XI9/NET36_XI19/XI9/MM10_g
+ N_VDD_XI19/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI9/MM11 N_XI19/XI9/NET36_XI19/XI9/MM11_d N_XI19/XI9/NET35_XI19/XI9/MM11_g
+ N_VDD_XI19/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI10/MM2 N_XI19/XI10/NET34_XI19/XI10/MM2_d
+ N_XI19/XI10/NET33_XI19/XI10/MM2_g N_VSS_XI19/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI10/MM3 N_XI19/XI10/NET33_XI19/XI10/MM3_d N_WL<34>_XI19/XI10/MM3_g
+ N_BLN<5>_XI19/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI10/MM0 N_XI19/XI10/NET34_XI19/XI10/MM0_d N_WL<34>_XI19/XI10/MM0_g
+ N_BL<5>_XI19/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI10/MM1 N_XI19/XI10/NET33_XI19/XI10/MM1_d
+ N_XI19/XI10/NET34_XI19/XI10/MM1_g N_VSS_XI19/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI10/MM9 N_XI19/XI10/NET36_XI19/XI10/MM9_d N_WL<35>_XI19/XI10/MM9_g
+ N_BL<5>_XI19/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI10/MM6 N_XI19/XI10/NET35_XI19/XI10/MM6_d
+ N_XI19/XI10/NET36_XI19/XI10/MM6_g N_VSS_XI19/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI10/MM7 N_XI19/XI10/NET36_XI19/XI10/MM7_d
+ N_XI19/XI10/NET35_XI19/XI10/MM7_g N_VSS_XI19/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI10/MM8 N_XI19/XI10/NET35_XI19/XI10/MM8_d N_WL<35>_XI19/XI10/MM8_g
+ N_BLN<5>_XI19/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI10/MM5 N_XI19/XI10/NET34_XI19/XI10/MM5_d
+ N_XI19/XI10/NET33_XI19/XI10/MM5_g N_VDD_XI19/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI10/MM4 N_XI19/XI10/NET33_XI19/XI10/MM4_d
+ N_XI19/XI10/NET34_XI19/XI10/MM4_g N_VDD_XI19/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI10/MM10 N_XI19/XI10/NET35_XI19/XI10/MM10_d
+ N_XI19/XI10/NET36_XI19/XI10/MM10_g N_VDD_XI19/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI10/MM11 N_XI19/XI10/NET36_XI19/XI10/MM11_d
+ N_XI19/XI10/NET35_XI19/XI10/MM11_g N_VDD_XI19/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI11/MM2 N_XI19/XI11/NET34_XI19/XI11/MM2_d
+ N_XI19/XI11/NET33_XI19/XI11/MM2_g N_VSS_XI19/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI11/MM3 N_XI19/XI11/NET33_XI19/XI11/MM3_d N_WL<34>_XI19/XI11/MM3_g
+ N_BLN<4>_XI19/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI11/MM0 N_XI19/XI11/NET34_XI19/XI11/MM0_d N_WL<34>_XI19/XI11/MM0_g
+ N_BL<4>_XI19/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI11/MM1 N_XI19/XI11/NET33_XI19/XI11/MM1_d
+ N_XI19/XI11/NET34_XI19/XI11/MM1_g N_VSS_XI19/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI11/MM9 N_XI19/XI11/NET36_XI19/XI11/MM9_d N_WL<35>_XI19/XI11/MM9_g
+ N_BL<4>_XI19/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI11/MM6 N_XI19/XI11/NET35_XI19/XI11/MM6_d
+ N_XI19/XI11/NET36_XI19/XI11/MM6_g N_VSS_XI19/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI11/MM7 N_XI19/XI11/NET36_XI19/XI11/MM7_d
+ N_XI19/XI11/NET35_XI19/XI11/MM7_g N_VSS_XI19/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI11/MM8 N_XI19/XI11/NET35_XI19/XI11/MM8_d N_WL<35>_XI19/XI11/MM8_g
+ N_BLN<4>_XI19/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI11/MM5 N_XI19/XI11/NET34_XI19/XI11/MM5_d
+ N_XI19/XI11/NET33_XI19/XI11/MM5_g N_VDD_XI19/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI11/MM4 N_XI19/XI11/NET33_XI19/XI11/MM4_d
+ N_XI19/XI11/NET34_XI19/XI11/MM4_g N_VDD_XI19/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI11/MM10 N_XI19/XI11/NET35_XI19/XI11/MM10_d
+ N_XI19/XI11/NET36_XI19/XI11/MM10_g N_VDD_XI19/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI11/MM11 N_XI19/XI11/NET36_XI19/XI11/MM11_d
+ N_XI19/XI11/NET35_XI19/XI11/MM11_g N_VDD_XI19/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI12/MM2 N_XI19/XI12/NET34_XI19/XI12/MM2_d
+ N_XI19/XI12/NET33_XI19/XI12/MM2_g N_VSS_XI19/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI12/MM3 N_XI19/XI12/NET33_XI19/XI12/MM3_d N_WL<34>_XI19/XI12/MM3_g
+ N_BLN<3>_XI19/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI12/MM0 N_XI19/XI12/NET34_XI19/XI12/MM0_d N_WL<34>_XI19/XI12/MM0_g
+ N_BL<3>_XI19/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI12/MM1 N_XI19/XI12/NET33_XI19/XI12/MM1_d
+ N_XI19/XI12/NET34_XI19/XI12/MM1_g N_VSS_XI19/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI12/MM9 N_XI19/XI12/NET36_XI19/XI12/MM9_d N_WL<35>_XI19/XI12/MM9_g
+ N_BL<3>_XI19/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI12/MM6 N_XI19/XI12/NET35_XI19/XI12/MM6_d
+ N_XI19/XI12/NET36_XI19/XI12/MM6_g N_VSS_XI19/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI12/MM7 N_XI19/XI12/NET36_XI19/XI12/MM7_d
+ N_XI19/XI12/NET35_XI19/XI12/MM7_g N_VSS_XI19/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI12/MM8 N_XI19/XI12/NET35_XI19/XI12/MM8_d N_WL<35>_XI19/XI12/MM8_g
+ N_BLN<3>_XI19/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI12/MM5 N_XI19/XI12/NET34_XI19/XI12/MM5_d
+ N_XI19/XI12/NET33_XI19/XI12/MM5_g N_VDD_XI19/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI12/MM4 N_XI19/XI12/NET33_XI19/XI12/MM4_d
+ N_XI19/XI12/NET34_XI19/XI12/MM4_g N_VDD_XI19/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI12/MM10 N_XI19/XI12/NET35_XI19/XI12/MM10_d
+ N_XI19/XI12/NET36_XI19/XI12/MM10_g N_VDD_XI19/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI12/MM11 N_XI19/XI12/NET36_XI19/XI12/MM11_d
+ N_XI19/XI12/NET35_XI19/XI12/MM11_g N_VDD_XI19/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI13/MM2 N_XI19/XI13/NET34_XI19/XI13/MM2_d
+ N_XI19/XI13/NET33_XI19/XI13/MM2_g N_VSS_XI19/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI13/MM3 N_XI19/XI13/NET33_XI19/XI13/MM3_d N_WL<34>_XI19/XI13/MM3_g
+ N_BLN<2>_XI19/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI13/MM0 N_XI19/XI13/NET34_XI19/XI13/MM0_d N_WL<34>_XI19/XI13/MM0_g
+ N_BL<2>_XI19/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI13/MM1 N_XI19/XI13/NET33_XI19/XI13/MM1_d
+ N_XI19/XI13/NET34_XI19/XI13/MM1_g N_VSS_XI19/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI13/MM9 N_XI19/XI13/NET36_XI19/XI13/MM9_d N_WL<35>_XI19/XI13/MM9_g
+ N_BL<2>_XI19/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI13/MM6 N_XI19/XI13/NET35_XI19/XI13/MM6_d
+ N_XI19/XI13/NET36_XI19/XI13/MM6_g N_VSS_XI19/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI13/MM7 N_XI19/XI13/NET36_XI19/XI13/MM7_d
+ N_XI19/XI13/NET35_XI19/XI13/MM7_g N_VSS_XI19/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI13/MM8 N_XI19/XI13/NET35_XI19/XI13/MM8_d N_WL<35>_XI19/XI13/MM8_g
+ N_BLN<2>_XI19/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI13/MM5 N_XI19/XI13/NET34_XI19/XI13/MM5_d
+ N_XI19/XI13/NET33_XI19/XI13/MM5_g N_VDD_XI19/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI13/MM4 N_XI19/XI13/NET33_XI19/XI13/MM4_d
+ N_XI19/XI13/NET34_XI19/XI13/MM4_g N_VDD_XI19/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI13/MM10 N_XI19/XI13/NET35_XI19/XI13/MM10_d
+ N_XI19/XI13/NET36_XI19/XI13/MM10_g N_VDD_XI19/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI13/MM11 N_XI19/XI13/NET36_XI19/XI13/MM11_d
+ N_XI19/XI13/NET35_XI19/XI13/MM11_g N_VDD_XI19/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI14/MM2 N_XI19/XI14/NET34_XI19/XI14/MM2_d
+ N_XI19/XI14/NET33_XI19/XI14/MM2_g N_VSS_XI19/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI14/MM3 N_XI19/XI14/NET33_XI19/XI14/MM3_d N_WL<34>_XI19/XI14/MM3_g
+ N_BLN<1>_XI19/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI14/MM0 N_XI19/XI14/NET34_XI19/XI14/MM0_d N_WL<34>_XI19/XI14/MM0_g
+ N_BL<1>_XI19/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI14/MM1 N_XI19/XI14/NET33_XI19/XI14/MM1_d
+ N_XI19/XI14/NET34_XI19/XI14/MM1_g N_VSS_XI19/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI14/MM9 N_XI19/XI14/NET36_XI19/XI14/MM9_d N_WL<35>_XI19/XI14/MM9_g
+ N_BL<1>_XI19/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI14/MM6 N_XI19/XI14/NET35_XI19/XI14/MM6_d
+ N_XI19/XI14/NET36_XI19/XI14/MM6_g N_VSS_XI19/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI14/MM7 N_XI19/XI14/NET36_XI19/XI14/MM7_d
+ N_XI19/XI14/NET35_XI19/XI14/MM7_g N_VSS_XI19/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI14/MM8 N_XI19/XI14/NET35_XI19/XI14/MM8_d N_WL<35>_XI19/XI14/MM8_g
+ N_BLN<1>_XI19/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI14/MM5 N_XI19/XI14/NET34_XI19/XI14/MM5_d
+ N_XI19/XI14/NET33_XI19/XI14/MM5_g N_VDD_XI19/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI14/MM4 N_XI19/XI14/NET33_XI19/XI14/MM4_d
+ N_XI19/XI14/NET34_XI19/XI14/MM4_g N_VDD_XI19/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI14/MM10 N_XI19/XI14/NET35_XI19/XI14/MM10_d
+ N_XI19/XI14/NET36_XI19/XI14/MM10_g N_VDD_XI19/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI14/MM11 N_XI19/XI14/NET36_XI19/XI14/MM11_d
+ N_XI19/XI14/NET35_XI19/XI14/MM11_g N_VDD_XI19/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI15/MM2 N_XI19/XI15/NET34_XI19/XI15/MM2_d
+ N_XI19/XI15/NET33_XI19/XI15/MM2_g N_VSS_XI19/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI15/MM3 N_XI19/XI15/NET33_XI19/XI15/MM3_d N_WL<34>_XI19/XI15/MM3_g
+ N_BLN<0>_XI19/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI15/MM0 N_XI19/XI15/NET34_XI19/XI15/MM0_d N_WL<34>_XI19/XI15/MM0_g
+ N_BL<0>_XI19/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI15/MM1 N_XI19/XI15/NET33_XI19/XI15/MM1_d
+ N_XI19/XI15/NET34_XI19/XI15/MM1_g N_VSS_XI19/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI15/MM9 N_XI19/XI15/NET36_XI19/XI15/MM9_d N_WL<35>_XI19/XI15/MM9_g
+ N_BL<0>_XI19/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI15/MM6 N_XI19/XI15/NET35_XI19/XI15/MM6_d
+ N_XI19/XI15/NET36_XI19/XI15/MM6_g N_VSS_XI19/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI15/MM7 N_XI19/XI15/NET36_XI19/XI15/MM7_d
+ N_XI19/XI15/NET35_XI19/XI15/MM7_g N_VSS_XI19/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI19/XI15/MM8 N_XI19/XI15/NET35_XI19/XI15/MM8_d N_WL<35>_XI19/XI15/MM8_g
+ N_BLN<0>_XI19/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI19/XI15/MM5 N_XI19/XI15/NET34_XI19/XI15/MM5_d
+ N_XI19/XI15/NET33_XI19/XI15/MM5_g N_VDD_XI19/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI15/MM4 N_XI19/XI15/NET33_XI19/XI15/MM4_d
+ N_XI19/XI15/NET34_XI19/XI15/MM4_g N_VDD_XI19/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI15/MM10 N_XI19/XI15/NET35_XI19/XI15/MM10_d
+ N_XI19/XI15/NET36_XI19/XI15/MM10_g N_VDD_XI19/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI19/XI15/MM11 N_XI19/XI15/NET36_XI19/XI15/MM11_d
+ N_XI19/XI15/NET35_XI19/XI15/MM11_g N_VDD_XI19/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI0/MM2 N_XI20/XI0/NET34_XI20/XI0/MM2_d N_XI20/XI0/NET33_XI20/XI0/MM2_g
+ N_VSS_XI20/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI0/MM3 N_XI20/XI0/NET33_XI20/XI0/MM3_d N_WL<36>_XI20/XI0/MM3_g
+ N_BLN<15>_XI20/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI0/MM0 N_XI20/XI0/NET34_XI20/XI0/MM0_d N_WL<36>_XI20/XI0/MM0_g
+ N_BL<15>_XI20/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI0/MM1 N_XI20/XI0/NET33_XI20/XI0/MM1_d N_XI20/XI0/NET34_XI20/XI0/MM1_g
+ N_VSS_XI20/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI0/MM9 N_XI20/XI0/NET36_XI20/XI0/MM9_d N_WL<37>_XI20/XI0/MM9_g
+ N_BL<15>_XI20/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI0/MM6 N_XI20/XI0/NET35_XI20/XI0/MM6_d N_XI20/XI0/NET36_XI20/XI0/MM6_g
+ N_VSS_XI20/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI0/MM7 N_XI20/XI0/NET36_XI20/XI0/MM7_d N_XI20/XI0/NET35_XI20/XI0/MM7_g
+ N_VSS_XI20/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI0/MM8 N_XI20/XI0/NET35_XI20/XI0/MM8_d N_WL<37>_XI20/XI0/MM8_g
+ N_BLN<15>_XI20/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI0/MM5 N_XI20/XI0/NET34_XI20/XI0/MM5_d N_XI20/XI0/NET33_XI20/XI0/MM5_g
+ N_VDD_XI20/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI0/MM4 N_XI20/XI0/NET33_XI20/XI0/MM4_d N_XI20/XI0/NET34_XI20/XI0/MM4_g
+ N_VDD_XI20/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI0/MM10 N_XI20/XI0/NET35_XI20/XI0/MM10_d N_XI20/XI0/NET36_XI20/XI0/MM10_g
+ N_VDD_XI20/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI0/MM11 N_XI20/XI0/NET36_XI20/XI0/MM11_d N_XI20/XI0/NET35_XI20/XI0/MM11_g
+ N_VDD_XI20/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI1/MM2 N_XI20/XI1/NET34_XI20/XI1/MM2_d N_XI20/XI1/NET33_XI20/XI1/MM2_g
+ N_VSS_XI20/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI1/MM3 N_XI20/XI1/NET33_XI20/XI1/MM3_d N_WL<36>_XI20/XI1/MM3_g
+ N_BLN<14>_XI20/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI1/MM0 N_XI20/XI1/NET34_XI20/XI1/MM0_d N_WL<36>_XI20/XI1/MM0_g
+ N_BL<14>_XI20/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI1/MM1 N_XI20/XI1/NET33_XI20/XI1/MM1_d N_XI20/XI1/NET34_XI20/XI1/MM1_g
+ N_VSS_XI20/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI1/MM9 N_XI20/XI1/NET36_XI20/XI1/MM9_d N_WL<37>_XI20/XI1/MM9_g
+ N_BL<14>_XI20/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI1/MM6 N_XI20/XI1/NET35_XI20/XI1/MM6_d N_XI20/XI1/NET36_XI20/XI1/MM6_g
+ N_VSS_XI20/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI1/MM7 N_XI20/XI1/NET36_XI20/XI1/MM7_d N_XI20/XI1/NET35_XI20/XI1/MM7_g
+ N_VSS_XI20/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI1/MM8 N_XI20/XI1/NET35_XI20/XI1/MM8_d N_WL<37>_XI20/XI1/MM8_g
+ N_BLN<14>_XI20/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI1/MM5 N_XI20/XI1/NET34_XI20/XI1/MM5_d N_XI20/XI1/NET33_XI20/XI1/MM5_g
+ N_VDD_XI20/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI1/MM4 N_XI20/XI1/NET33_XI20/XI1/MM4_d N_XI20/XI1/NET34_XI20/XI1/MM4_g
+ N_VDD_XI20/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI1/MM10 N_XI20/XI1/NET35_XI20/XI1/MM10_d N_XI20/XI1/NET36_XI20/XI1/MM10_g
+ N_VDD_XI20/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI1/MM11 N_XI20/XI1/NET36_XI20/XI1/MM11_d N_XI20/XI1/NET35_XI20/XI1/MM11_g
+ N_VDD_XI20/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI2/MM2 N_XI20/XI2/NET34_XI20/XI2/MM2_d N_XI20/XI2/NET33_XI20/XI2/MM2_g
+ N_VSS_XI20/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI2/MM3 N_XI20/XI2/NET33_XI20/XI2/MM3_d N_WL<36>_XI20/XI2/MM3_g
+ N_BLN<13>_XI20/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI2/MM0 N_XI20/XI2/NET34_XI20/XI2/MM0_d N_WL<36>_XI20/XI2/MM0_g
+ N_BL<13>_XI20/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI2/MM1 N_XI20/XI2/NET33_XI20/XI2/MM1_d N_XI20/XI2/NET34_XI20/XI2/MM1_g
+ N_VSS_XI20/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI2/MM9 N_XI20/XI2/NET36_XI20/XI2/MM9_d N_WL<37>_XI20/XI2/MM9_g
+ N_BL<13>_XI20/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI2/MM6 N_XI20/XI2/NET35_XI20/XI2/MM6_d N_XI20/XI2/NET36_XI20/XI2/MM6_g
+ N_VSS_XI20/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI2/MM7 N_XI20/XI2/NET36_XI20/XI2/MM7_d N_XI20/XI2/NET35_XI20/XI2/MM7_g
+ N_VSS_XI20/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI2/MM8 N_XI20/XI2/NET35_XI20/XI2/MM8_d N_WL<37>_XI20/XI2/MM8_g
+ N_BLN<13>_XI20/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI2/MM5 N_XI20/XI2/NET34_XI20/XI2/MM5_d N_XI20/XI2/NET33_XI20/XI2/MM5_g
+ N_VDD_XI20/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI2/MM4 N_XI20/XI2/NET33_XI20/XI2/MM4_d N_XI20/XI2/NET34_XI20/XI2/MM4_g
+ N_VDD_XI20/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI2/MM10 N_XI20/XI2/NET35_XI20/XI2/MM10_d N_XI20/XI2/NET36_XI20/XI2/MM10_g
+ N_VDD_XI20/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI2/MM11 N_XI20/XI2/NET36_XI20/XI2/MM11_d N_XI20/XI2/NET35_XI20/XI2/MM11_g
+ N_VDD_XI20/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI3/MM2 N_XI20/XI3/NET34_XI20/XI3/MM2_d N_XI20/XI3/NET33_XI20/XI3/MM2_g
+ N_VSS_XI20/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI3/MM3 N_XI20/XI3/NET33_XI20/XI3/MM3_d N_WL<36>_XI20/XI3/MM3_g
+ N_BLN<12>_XI20/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI3/MM0 N_XI20/XI3/NET34_XI20/XI3/MM0_d N_WL<36>_XI20/XI3/MM0_g
+ N_BL<12>_XI20/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI3/MM1 N_XI20/XI3/NET33_XI20/XI3/MM1_d N_XI20/XI3/NET34_XI20/XI3/MM1_g
+ N_VSS_XI20/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI3/MM9 N_XI20/XI3/NET36_XI20/XI3/MM9_d N_WL<37>_XI20/XI3/MM9_g
+ N_BL<12>_XI20/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI3/MM6 N_XI20/XI3/NET35_XI20/XI3/MM6_d N_XI20/XI3/NET36_XI20/XI3/MM6_g
+ N_VSS_XI20/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI3/MM7 N_XI20/XI3/NET36_XI20/XI3/MM7_d N_XI20/XI3/NET35_XI20/XI3/MM7_g
+ N_VSS_XI20/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI3/MM8 N_XI20/XI3/NET35_XI20/XI3/MM8_d N_WL<37>_XI20/XI3/MM8_g
+ N_BLN<12>_XI20/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI3/MM5 N_XI20/XI3/NET34_XI20/XI3/MM5_d N_XI20/XI3/NET33_XI20/XI3/MM5_g
+ N_VDD_XI20/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI3/MM4 N_XI20/XI3/NET33_XI20/XI3/MM4_d N_XI20/XI3/NET34_XI20/XI3/MM4_g
+ N_VDD_XI20/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI3/MM10 N_XI20/XI3/NET35_XI20/XI3/MM10_d N_XI20/XI3/NET36_XI20/XI3/MM10_g
+ N_VDD_XI20/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI3/MM11 N_XI20/XI3/NET36_XI20/XI3/MM11_d N_XI20/XI3/NET35_XI20/XI3/MM11_g
+ N_VDD_XI20/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI4/MM2 N_XI20/XI4/NET34_XI20/XI4/MM2_d N_XI20/XI4/NET33_XI20/XI4/MM2_g
+ N_VSS_XI20/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI4/MM3 N_XI20/XI4/NET33_XI20/XI4/MM3_d N_WL<36>_XI20/XI4/MM3_g
+ N_BLN<11>_XI20/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI4/MM0 N_XI20/XI4/NET34_XI20/XI4/MM0_d N_WL<36>_XI20/XI4/MM0_g
+ N_BL<11>_XI20/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI4/MM1 N_XI20/XI4/NET33_XI20/XI4/MM1_d N_XI20/XI4/NET34_XI20/XI4/MM1_g
+ N_VSS_XI20/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI4/MM9 N_XI20/XI4/NET36_XI20/XI4/MM9_d N_WL<37>_XI20/XI4/MM9_g
+ N_BL<11>_XI20/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI4/MM6 N_XI20/XI4/NET35_XI20/XI4/MM6_d N_XI20/XI4/NET36_XI20/XI4/MM6_g
+ N_VSS_XI20/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI4/MM7 N_XI20/XI4/NET36_XI20/XI4/MM7_d N_XI20/XI4/NET35_XI20/XI4/MM7_g
+ N_VSS_XI20/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI4/MM8 N_XI20/XI4/NET35_XI20/XI4/MM8_d N_WL<37>_XI20/XI4/MM8_g
+ N_BLN<11>_XI20/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI4/MM5 N_XI20/XI4/NET34_XI20/XI4/MM5_d N_XI20/XI4/NET33_XI20/XI4/MM5_g
+ N_VDD_XI20/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI4/MM4 N_XI20/XI4/NET33_XI20/XI4/MM4_d N_XI20/XI4/NET34_XI20/XI4/MM4_g
+ N_VDD_XI20/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI4/MM10 N_XI20/XI4/NET35_XI20/XI4/MM10_d N_XI20/XI4/NET36_XI20/XI4/MM10_g
+ N_VDD_XI20/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI4/MM11 N_XI20/XI4/NET36_XI20/XI4/MM11_d N_XI20/XI4/NET35_XI20/XI4/MM11_g
+ N_VDD_XI20/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI5/MM2 N_XI20/XI5/NET34_XI20/XI5/MM2_d N_XI20/XI5/NET33_XI20/XI5/MM2_g
+ N_VSS_XI20/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI5/MM3 N_XI20/XI5/NET33_XI20/XI5/MM3_d N_WL<36>_XI20/XI5/MM3_g
+ N_BLN<10>_XI20/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI5/MM0 N_XI20/XI5/NET34_XI20/XI5/MM0_d N_WL<36>_XI20/XI5/MM0_g
+ N_BL<10>_XI20/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI5/MM1 N_XI20/XI5/NET33_XI20/XI5/MM1_d N_XI20/XI5/NET34_XI20/XI5/MM1_g
+ N_VSS_XI20/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI5/MM9 N_XI20/XI5/NET36_XI20/XI5/MM9_d N_WL<37>_XI20/XI5/MM9_g
+ N_BL<10>_XI20/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI5/MM6 N_XI20/XI5/NET35_XI20/XI5/MM6_d N_XI20/XI5/NET36_XI20/XI5/MM6_g
+ N_VSS_XI20/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI5/MM7 N_XI20/XI5/NET36_XI20/XI5/MM7_d N_XI20/XI5/NET35_XI20/XI5/MM7_g
+ N_VSS_XI20/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI5/MM8 N_XI20/XI5/NET35_XI20/XI5/MM8_d N_WL<37>_XI20/XI5/MM8_g
+ N_BLN<10>_XI20/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI5/MM5 N_XI20/XI5/NET34_XI20/XI5/MM5_d N_XI20/XI5/NET33_XI20/XI5/MM5_g
+ N_VDD_XI20/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI5/MM4 N_XI20/XI5/NET33_XI20/XI5/MM4_d N_XI20/XI5/NET34_XI20/XI5/MM4_g
+ N_VDD_XI20/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI5/MM10 N_XI20/XI5/NET35_XI20/XI5/MM10_d N_XI20/XI5/NET36_XI20/XI5/MM10_g
+ N_VDD_XI20/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI5/MM11 N_XI20/XI5/NET36_XI20/XI5/MM11_d N_XI20/XI5/NET35_XI20/XI5/MM11_g
+ N_VDD_XI20/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI6/MM2 N_XI20/XI6/NET34_XI20/XI6/MM2_d N_XI20/XI6/NET33_XI20/XI6/MM2_g
+ N_VSS_XI20/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM3 N_XI20/XI6/NET33_XI20/XI6/MM3_d N_WL<36>_XI20/XI6/MM3_g
+ N_BLN<9>_XI20/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM0 N_XI20/XI6/NET34_XI20/XI6/MM0_d N_WL<36>_XI20/XI6/MM0_g
+ N_BL<9>_XI20/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM1 N_XI20/XI6/NET33_XI20/XI6/MM1_d N_XI20/XI6/NET34_XI20/XI6/MM1_g
+ N_VSS_XI20/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM9 N_XI20/XI6/NET36_XI20/XI6/MM9_d N_WL<37>_XI20/XI6/MM9_g
+ N_BL<9>_XI20/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM6 N_XI20/XI6/NET35_XI20/XI6/MM6_d N_XI20/XI6/NET36_XI20/XI6/MM6_g
+ N_VSS_XI20/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM7 N_XI20/XI6/NET36_XI20/XI6/MM7_d N_XI20/XI6/NET35_XI20/XI6/MM7_g
+ N_VSS_XI20/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM8 N_XI20/XI6/NET35_XI20/XI6/MM8_d N_WL<37>_XI20/XI6/MM8_g
+ N_BLN<9>_XI20/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI6/MM5 N_XI20/XI6/NET34_XI20/XI6/MM5_d N_XI20/XI6/NET33_XI20/XI6/MM5_g
+ N_VDD_XI20/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI6/MM4 N_XI20/XI6/NET33_XI20/XI6/MM4_d N_XI20/XI6/NET34_XI20/XI6/MM4_g
+ N_VDD_XI20/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI6/MM10 N_XI20/XI6/NET35_XI20/XI6/MM10_d N_XI20/XI6/NET36_XI20/XI6/MM10_g
+ N_VDD_XI20/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI6/MM11 N_XI20/XI6/NET36_XI20/XI6/MM11_d N_XI20/XI6/NET35_XI20/XI6/MM11_g
+ N_VDD_XI20/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI7/MM2 N_XI20/XI7/NET34_XI20/XI7/MM2_d N_XI20/XI7/NET33_XI20/XI7/MM2_g
+ N_VSS_XI20/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM3 N_XI20/XI7/NET33_XI20/XI7/MM3_d N_WL<36>_XI20/XI7/MM3_g
+ N_BLN<8>_XI20/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM0 N_XI20/XI7/NET34_XI20/XI7/MM0_d N_WL<36>_XI20/XI7/MM0_g
+ N_BL<8>_XI20/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM1 N_XI20/XI7/NET33_XI20/XI7/MM1_d N_XI20/XI7/NET34_XI20/XI7/MM1_g
+ N_VSS_XI20/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM9 N_XI20/XI7/NET36_XI20/XI7/MM9_d N_WL<37>_XI20/XI7/MM9_g
+ N_BL<8>_XI20/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM6 N_XI20/XI7/NET35_XI20/XI7/MM6_d N_XI20/XI7/NET36_XI20/XI7/MM6_g
+ N_VSS_XI20/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM7 N_XI20/XI7/NET36_XI20/XI7/MM7_d N_XI20/XI7/NET35_XI20/XI7/MM7_g
+ N_VSS_XI20/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM8 N_XI20/XI7/NET35_XI20/XI7/MM8_d N_WL<37>_XI20/XI7/MM8_g
+ N_BLN<8>_XI20/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI7/MM5 N_XI20/XI7/NET34_XI20/XI7/MM5_d N_XI20/XI7/NET33_XI20/XI7/MM5_g
+ N_VDD_XI20/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI7/MM4 N_XI20/XI7/NET33_XI20/XI7/MM4_d N_XI20/XI7/NET34_XI20/XI7/MM4_g
+ N_VDD_XI20/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI7/MM10 N_XI20/XI7/NET35_XI20/XI7/MM10_d N_XI20/XI7/NET36_XI20/XI7/MM10_g
+ N_VDD_XI20/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI7/MM11 N_XI20/XI7/NET36_XI20/XI7/MM11_d N_XI20/XI7/NET35_XI20/XI7/MM11_g
+ N_VDD_XI20/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI8/MM2 N_XI20/XI8/NET34_XI20/XI8/MM2_d N_XI20/XI8/NET33_XI20/XI8/MM2_g
+ N_VSS_XI20/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM3 N_XI20/XI8/NET33_XI20/XI8/MM3_d N_WL<36>_XI20/XI8/MM3_g
+ N_BLN<7>_XI20/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM0 N_XI20/XI8/NET34_XI20/XI8/MM0_d N_WL<36>_XI20/XI8/MM0_g
+ N_BL<7>_XI20/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM1 N_XI20/XI8/NET33_XI20/XI8/MM1_d N_XI20/XI8/NET34_XI20/XI8/MM1_g
+ N_VSS_XI20/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM9 N_XI20/XI8/NET36_XI20/XI8/MM9_d N_WL<37>_XI20/XI8/MM9_g
+ N_BL<7>_XI20/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM6 N_XI20/XI8/NET35_XI20/XI8/MM6_d N_XI20/XI8/NET36_XI20/XI8/MM6_g
+ N_VSS_XI20/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM7 N_XI20/XI8/NET36_XI20/XI8/MM7_d N_XI20/XI8/NET35_XI20/XI8/MM7_g
+ N_VSS_XI20/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM8 N_XI20/XI8/NET35_XI20/XI8/MM8_d N_WL<37>_XI20/XI8/MM8_g
+ N_BLN<7>_XI20/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI8/MM5 N_XI20/XI8/NET34_XI20/XI8/MM5_d N_XI20/XI8/NET33_XI20/XI8/MM5_g
+ N_VDD_XI20/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI8/MM4 N_XI20/XI8/NET33_XI20/XI8/MM4_d N_XI20/XI8/NET34_XI20/XI8/MM4_g
+ N_VDD_XI20/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI8/MM10 N_XI20/XI8/NET35_XI20/XI8/MM10_d N_XI20/XI8/NET36_XI20/XI8/MM10_g
+ N_VDD_XI20/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI8/MM11 N_XI20/XI8/NET36_XI20/XI8/MM11_d N_XI20/XI8/NET35_XI20/XI8/MM11_g
+ N_VDD_XI20/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI9/MM2 N_XI20/XI9/NET34_XI20/XI9/MM2_d N_XI20/XI9/NET33_XI20/XI9/MM2_g
+ N_VSS_XI20/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM3 N_XI20/XI9/NET33_XI20/XI9/MM3_d N_WL<36>_XI20/XI9/MM3_g
+ N_BLN<6>_XI20/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM0 N_XI20/XI9/NET34_XI20/XI9/MM0_d N_WL<36>_XI20/XI9/MM0_g
+ N_BL<6>_XI20/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM1 N_XI20/XI9/NET33_XI20/XI9/MM1_d N_XI20/XI9/NET34_XI20/XI9/MM1_g
+ N_VSS_XI20/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM9 N_XI20/XI9/NET36_XI20/XI9/MM9_d N_WL<37>_XI20/XI9/MM9_g
+ N_BL<6>_XI20/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM6 N_XI20/XI9/NET35_XI20/XI9/MM6_d N_XI20/XI9/NET36_XI20/XI9/MM6_g
+ N_VSS_XI20/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM7 N_XI20/XI9/NET36_XI20/XI9/MM7_d N_XI20/XI9/NET35_XI20/XI9/MM7_g
+ N_VSS_XI20/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM8 N_XI20/XI9/NET35_XI20/XI9/MM8_d N_WL<37>_XI20/XI9/MM8_g
+ N_BLN<6>_XI20/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI9/MM5 N_XI20/XI9/NET34_XI20/XI9/MM5_d N_XI20/XI9/NET33_XI20/XI9/MM5_g
+ N_VDD_XI20/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI9/MM4 N_XI20/XI9/NET33_XI20/XI9/MM4_d N_XI20/XI9/NET34_XI20/XI9/MM4_g
+ N_VDD_XI20/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI9/MM10 N_XI20/XI9/NET35_XI20/XI9/MM10_d N_XI20/XI9/NET36_XI20/XI9/MM10_g
+ N_VDD_XI20/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI9/MM11 N_XI20/XI9/NET36_XI20/XI9/MM11_d N_XI20/XI9/NET35_XI20/XI9/MM11_g
+ N_VDD_XI20/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI10/MM2 N_XI20/XI10/NET34_XI20/XI10/MM2_d
+ N_XI20/XI10/NET33_XI20/XI10/MM2_g N_VSS_XI20/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI10/MM3 N_XI20/XI10/NET33_XI20/XI10/MM3_d N_WL<36>_XI20/XI10/MM3_g
+ N_BLN<5>_XI20/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI10/MM0 N_XI20/XI10/NET34_XI20/XI10/MM0_d N_WL<36>_XI20/XI10/MM0_g
+ N_BL<5>_XI20/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI10/MM1 N_XI20/XI10/NET33_XI20/XI10/MM1_d
+ N_XI20/XI10/NET34_XI20/XI10/MM1_g N_VSS_XI20/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI10/MM9 N_XI20/XI10/NET36_XI20/XI10/MM9_d N_WL<37>_XI20/XI10/MM9_g
+ N_BL<5>_XI20/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI10/MM6 N_XI20/XI10/NET35_XI20/XI10/MM6_d
+ N_XI20/XI10/NET36_XI20/XI10/MM6_g N_VSS_XI20/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI10/MM7 N_XI20/XI10/NET36_XI20/XI10/MM7_d
+ N_XI20/XI10/NET35_XI20/XI10/MM7_g N_VSS_XI20/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI10/MM8 N_XI20/XI10/NET35_XI20/XI10/MM8_d N_WL<37>_XI20/XI10/MM8_g
+ N_BLN<5>_XI20/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI10/MM5 N_XI20/XI10/NET34_XI20/XI10/MM5_d
+ N_XI20/XI10/NET33_XI20/XI10/MM5_g N_VDD_XI20/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI10/MM4 N_XI20/XI10/NET33_XI20/XI10/MM4_d
+ N_XI20/XI10/NET34_XI20/XI10/MM4_g N_VDD_XI20/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI10/MM10 N_XI20/XI10/NET35_XI20/XI10/MM10_d
+ N_XI20/XI10/NET36_XI20/XI10/MM10_g N_VDD_XI20/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI10/MM11 N_XI20/XI10/NET36_XI20/XI10/MM11_d
+ N_XI20/XI10/NET35_XI20/XI10/MM11_g N_VDD_XI20/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI11/MM2 N_XI20/XI11/NET34_XI20/XI11/MM2_d
+ N_XI20/XI11/NET33_XI20/XI11/MM2_g N_VSS_XI20/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI11/MM3 N_XI20/XI11/NET33_XI20/XI11/MM3_d N_WL<36>_XI20/XI11/MM3_g
+ N_BLN<4>_XI20/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI11/MM0 N_XI20/XI11/NET34_XI20/XI11/MM0_d N_WL<36>_XI20/XI11/MM0_g
+ N_BL<4>_XI20/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI11/MM1 N_XI20/XI11/NET33_XI20/XI11/MM1_d
+ N_XI20/XI11/NET34_XI20/XI11/MM1_g N_VSS_XI20/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI11/MM9 N_XI20/XI11/NET36_XI20/XI11/MM9_d N_WL<37>_XI20/XI11/MM9_g
+ N_BL<4>_XI20/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI11/MM6 N_XI20/XI11/NET35_XI20/XI11/MM6_d
+ N_XI20/XI11/NET36_XI20/XI11/MM6_g N_VSS_XI20/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI11/MM7 N_XI20/XI11/NET36_XI20/XI11/MM7_d
+ N_XI20/XI11/NET35_XI20/XI11/MM7_g N_VSS_XI20/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI11/MM8 N_XI20/XI11/NET35_XI20/XI11/MM8_d N_WL<37>_XI20/XI11/MM8_g
+ N_BLN<4>_XI20/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI11/MM5 N_XI20/XI11/NET34_XI20/XI11/MM5_d
+ N_XI20/XI11/NET33_XI20/XI11/MM5_g N_VDD_XI20/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI11/MM4 N_XI20/XI11/NET33_XI20/XI11/MM4_d
+ N_XI20/XI11/NET34_XI20/XI11/MM4_g N_VDD_XI20/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI11/MM10 N_XI20/XI11/NET35_XI20/XI11/MM10_d
+ N_XI20/XI11/NET36_XI20/XI11/MM10_g N_VDD_XI20/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI11/MM11 N_XI20/XI11/NET36_XI20/XI11/MM11_d
+ N_XI20/XI11/NET35_XI20/XI11/MM11_g N_VDD_XI20/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI12/MM2 N_XI20/XI12/NET34_XI20/XI12/MM2_d
+ N_XI20/XI12/NET33_XI20/XI12/MM2_g N_VSS_XI20/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI12/MM3 N_XI20/XI12/NET33_XI20/XI12/MM3_d N_WL<36>_XI20/XI12/MM3_g
+ N_BLN<3>_XI20/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI12/MM0 N_XI20/XI12/NET34_XI20/XI12/MM0_d N_WL<36>_XI20/XI12/MM0_g
+ N_BL<3>_XI20/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI12/MM1 N_XI20/XI12/NET33_XI20/XI12/MM1_d
+ N_XI20/XI12/NET34_XI20/XI12/MM1_g N_VSS_XI20/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI12/MM9 N_XI20/XI12/NET36_XI20/XI12/MM9_d N_WL<37>_XI20/XI12/MM9_g
+ N_BL<3>_XI20/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI12/MM6 N_XI20/XI12/NET35_XI20/XI12/MM6_d
+ N_XI20/XI12/NET36_XI20/XI12/MM6_g N_VSS_XI20/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI12/MM7 N_XI20/XI12/NET36_XI20/XI12/MM7_d
+ N_XI20/XI12/NET35_XI20/XI12/MM7_g N_VSS_XI20/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI12/MM8 N_XI20/XI12/NET35_XI20/XI12/MM8_d N_WL<37>_XI20/XI12/MM8_g
+ N_BLN<3>_XI20/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI12/MM5 N_XI20/XI12/NET34_XI20/XI12/MM5_d
+ N_XI20/XI12/NET33_XI20/XI12/MM5_g N_VDD_XI20/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI12/MM4 N_XI20/XI12/NET33_XI20/XI12/MM4_d
+ N_XI20/XI12/NET34_XI20/XI12/MM4_g N_VDD_XI20/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI12/MM10 N_XI20/XI12/NET35_XI20/XI12/MM10_d
+ N_XI20/XI12/NET36_XI20/XI12/MM10_g N_VDD_XI20/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI12/MM11 N_XI20/XI12/NET36_XI20/XI12/MM11_d
+ N_XI20/XI12/NET35_XI20/XI12/MM11_g N_VDD_XI20/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI13/MM2 N_XI20/XI13/NET34_XI20/XI13/MM2_d
+ N_XI20/XI13/NET33_XI20/XI13/MM2_g N_VSS_XI20/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI13/MM3 N_XI20/XI13/NET33_XI20/XI13/MM3_d N_WL<36>_XI20/XI13/MM3_g
+ N_BLN<2>_XI20/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI13/MM0 N_XI20/XI13/NET34_XI20/XI13/MM0_d N_WL<36>_XI20/XI13/MM0_g
+ N_BL<2>_XI20/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI13/MM1 N_XI20/XI13/NET33_XI20/XI13/MM1_d
+ N_XI20/XI13/NET34_XI20/XI13/MM1_g N_VSS_XI20/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI13/MM9 N_XI20/XI13/NET36_XI20/XI13/MM9_d N_WL<37>_XI20/XI13/MM9_g
+ N_BL<2>_XI20/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI13/MM6 N_XI20/XI13/NET35_XI20/XI13/MM6_d
+ N_XI20/XI13/NET36_XI20/XI13/MM6_g N_VSS_XI20/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI13/MM7 N_XI20/XI13/NET36_XI20/XI13/MM7_d
+ N_XI20/XI13/NET35_XI20/XI13/MM7_g N_VSS_XI20/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI13/MM8 N_XI20/XI13/NET35_XI20/XI13/MM8_d N_WL<37>_XI20/XI13/MM8_g
+ N_BLN<2>_XI20/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI13/MM5 N_XI20/XI13/NET34_XI20/XI13/MM5_d
+ N_XI20/XI13/NET33_XI20/XI13/MM5_g N_VDD_XI20/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI13/MM4 N_XI20/XI13/NET33_XI20/XI13/MM4_d
+ N_XI20/XI13/NET34_XI20/XI13/MM4_g N_VDD_XI20/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI13/MM10 N_XI20/XI13/NET35_XI20/XI13/MM10_d
+ N_XI20/XI13/NET36_XI20/XI13/MM10_g N_VDD_XI20/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI13/MM11 N_XI20/XI13/NET36_XI20/XI13/MM11_d
+ N_XI20/XI13/NET35_XI20/XI13/MM11_g N_VDD_XI20/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI14/MM2 N_XI20/XI14/NET34_XI20/XI14/MM2_d
+ N_XI20/XI14/NET33_XI20/XI14/MM2_g N_VSS_XI20/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI14/MM3 N_XI20/XI14/NET33_XI20/XI14/MM3_d N_WL<36>_XI20/XI14/MM3_g
+ N_BLN<1>_XI20/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI14/MM0 N_XI20/XI14/NET34_XI20/XI14/MM0_d N_WL<36>_XI20/XI14/MM0_g
+ N_BL<1>_XI20/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI14/MM1 N_XI20/XI14/NET33_XI20/XI14/MM1_d
+ N_XI20/XI14/NET34_XI20/XI14/MM1_g N_VSS_XI20/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI14/MM9 N_XI20/XI14/NET36_XI20/XI14/MM9_d N_WL<37>_XI20/XI14/MM9_g
+ N_BL<1>_XI20/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI14/MM6 N_XI20/XI14/NET35_XI20/XI14/MM6_d
+ N_XI20/XI14/NET36_XI20/XI14/MM6_g N_VSS_XI20/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI14/MM7 N_XI20/XI14/NET36_XI20/XI14/MM7_d
+ N_XI20/XI14/NET35_XI20/XI14/MM7_g N_VSS_XI20/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI14/MM8 N_XI20/XI14/NET35_XI20/XI14/MM8_d N_WL<37>_XI20/XI14/MM8_g
+ N_BLN<1>_XI20/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI14/MM5 N_XI20/XI14/NET34_XI20/XI14/MM5_d
+ N_XI20/XI14/NET33_XI20/XI14/MM5_g N_VDD_XI20/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI14/MM4 N_XI20/XI14/NET33_XI20/XI14/MM4_d
+ N_XI20/XI14/NET34_XI20/XI14/MM4_g N_VDD_XI20/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI14/MM10 N_XI20/XI14/NET35_XI20/XI14/MM10_d
+ N_XI20/XI14/NET36_XI20/XI14/MM10_g N_VDD_XI20/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI14/MM11 N_XI20/XI14/NET36_XI20/XI14/MM11_d
+ N_XI20/XI14/NET35_XI20/XI14/MM11_g N_VDD_XI20/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI15/MM2 N_XI20/XI15/NET34_XI20/XI15/MM2_d
+ N_XI20/XI15/NET33_XI20/XI15/MM2_g N_VSS_XI20/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI15/MM3 N_XI20/XI15/NET33_XI20/XI15/MM3_d N_WL<36>_XI20/XI15/MM3_g
+ N_BLN<0>_XI20/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI15/MM0 N_XI20/XI15/NET34_XI20/XI15/MM0_d N_WL<36>_XI20/XI15/MM0_g
+ N_BL<0>_XI20/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI15/MM1 N_XI20/XI15/NET33_XI20/XI15/MM1_d
+ N_XI20/XI15/NET34_XI20/XI15/MM1_g N_VSS_XI20/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI15/MM9 N_XI20/XI15/NET36_XI20/XI15/MM9_d N_WL<37>_XI20/XI15/MM9_g
+ N_BL<0>_XI20/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI15/MM6 N_XI20/XI15/NET35_XI20/XI15/MM6_d
+ N_XI20/XI15/NET36_XI20/XI15/MM6_g N_VSS_XI20/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI15/MM7 N_XI20/XI15/NET36_XI20/XI15/MM7_d
+ N_XI20/XI15/NET35_XI20/XI15/MM7_g N_VSS_XI20/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI20/XI15/MM8 N_XI20/XI15/NET35_XI20/XI15/MM8_d N_WL<37>_XI20/XI15/MM8_g
+ N_BLN<0>_XI20/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI20/XI15/MM5 N_XI20/XI15/NET34_XI20/XI15/MM5_d
+ N_XI20/XI15/NET33_XI20/XI15/MM5_g N_VDD_XI20/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI15/MM4 N_XI20/XI15/NET33_XI20/XI15/MM4_d
+ N_XI20/XI15/NET34_XI20/XI15/MM4_g N_VDD_XI20/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI15/MM10 N_XI20/XI15/NET35_XI20/XI15/MM10_d
+ N_XI20/XI15/NET36_XI20/XI15/MM10_g N_VDD_XI20/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI20/XI15/MM11 N_XI20/XI15/NET36_XI20/XI15/MM11_d
+ N_XI20/XI15/NET35_XI20/XI15/MM11_g N_VDD_XI20/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI0/MM2 N_XI21/XI0/NET34_XI21/XI0/MM2_d N_XI21/XI0/NET33_XI21/XI0/MM2_g
+ N_VSS_XI21/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI0/MM3 N_XI21/XI0/NET33_XI21/XI0/MM3_d N_WL<38>_XI21/XI0/MM3_g
+ N_BLN<15>_XI21/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI0/MM0 N_XI21/XI0/NET34_XI21/XI0/MM0_d N_WL<38>_XI21/XI0/MM0_g
+ N_BL<15>_XI21/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI0/MM1 N_XI21/XI0/NET33_XI21/XI0/MM1_d N_XI21/XI0/NET34_XI21/XI0/MM1_g
+ N_VSS_XI21/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI0/MM9 N_XI21/XI0/NET36_XI21/XI0/MM9_d N_WL<39>_XI21/XI0/MM9_g
+ N_BL<15>_XI21/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI0/MM6 N_XI21/XI0/NET35_XI21/XI0/MM6_d N_XI21/XI0/NET36_XI21/XI0/MM6_g
+ N_VSS_XI21/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI0/MM7 N_XI21/XI0/NET36_XI21/XI0/MM7_d N_XI21/XI0/NET35_XI21/XI0/MM7_g
+ N_VSS_XI21/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI0/MM8 N_XI21/XI0/NET35_XI21/XI0/MM8_d N_WL<39>_XI21/XI0/MM8_g
+ N_BLN<15>_XI21/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI0/MM5 N_XI21/XI0/NET34_XI21/XI0/MM5_d N_XI21/XI0/NET33_XI21/XI0/MM5_g
+ N_VDD_XI21/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI0/MM4 N_XI21/XI0/NET33_XI21/XI0/MM4_d N_XI21/XI0/NET34_XI21/XI0/MM4_g
+ N_VDD_XI21/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI0/MM10 N_XI21/XI0/NET35_XI21/XI0/MM10_d N_XI21/XI0/NET36_XI21/XI0/MM10_g
+ N_VDD_XI21/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI0/MM11 N_XI21/XI0/NET36_XI21/XI0/MM11_d N_XI21/XI0/NET35_XI21/XI0/MM11_g
+ N_VDD_XI21/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI1/MM2 N_XI21/XI1/NET34_XI21/XI1/MM2_d N_XI21/XI1/NET33_XI21/XI1/MM2_g
+ N_VSS_XI21/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI1/MM3 N_XI21/XI1/NET33_XI21/XI1/MM3_d N_WL<38>_XI21/XI1/MM3_g
+ N_BLN<14>_XI21/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI1/MM0 N_XI21/XI1/NET34_XI21/XI1/MM0_d N_WL<38>_XI21/XI1/MM0_g
+ N_BL<14>_XI21/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI1/MM1 N_XI21/XI1/NET33_XI21/XI1/MM1_d N_XI21/XI1/NET34_XI21/XI1/MM1_g
+ N_VSS_XI21/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI1/MM9 N_XI21/XI1/NET36_XI21/XI1/MM9_d N_WL<39>_XI21/XI1/MM9_g
+ N_BL<14>_XI21/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI1/MM6 N_XI21/XI1/NET35_XI21/XI1/MM6_d N_XI21/XI1/NET36_XI21/XI1/MM6_g
+ N_VSS_XI21/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI1/MM7 N_XI21/XI1/NET36_XI21/XI1/MM7_d N_XI21/XI1/NET35_XI21/XI1/MM7_g
+ N_VSS_XI21/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI1/MM8 N_XI21/XI1/NET35_XI21/XI1/MM8_d N_WL<39>_XI21/XI1/MM8_g
+ N_BLN<14>_XI21/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI1/MM5 N_XI21/XI1/NET34_XI21/XI1/MM5_d N_XI21/XI1/NET33_XI21/XI1/MM5_g
+ N_VDD_XI21/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI1/MM4 N_XI21/XI1/NET33_XI21/XI1/MM4_d N_XI21/XI1/NET34_XI21/XI1/MM4_g
+ N_VDD_XI21/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI1/MM10 N_XI21/XI1/NET35_XI21/XI1/MM10_d N_XI21/XI1/NET36_XI21/XI1/MM10_g
+ N_VDD_XI21/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI1/MM11 N_XI21/XI1/NET36_XI21/XI1/MM11_d N_XI21/XI1/NET35_XI21/XI1/MM11_g
+ N_VDD_XI21/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI2/MM2 N_XI21/XI2/NET34_XI21/XI2/MM2_d N_XI21/XI2/NET33_XI21/XI2/MM2_g
+ N_VSS_XI21/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI2/MM3 N_XI21/XI2/NET33_XI21/XI2/MM3_d N_WL<38>_XI21/XI2/MM3_g
+ N_BLN<13>_XI21/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI2/MM0 N_XI21/XI2/NET34_XI21/XI2/MM0_d N_WL<38>_XI21/XI2/MM0_g
+ N_BL<13>_XI21/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI2/MM1 N_XI21/XI2/NET33_XI21/XI2/MM1_d N_XI21/XI2/NET34_XI21/XI2/MM1_g
+ N_VSS_XI21/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI2/MM9 N_XI21/XI2/NET36_XI21/XI2/MM9_d N_WL<39>_XI21/XI2/MM9_g
+ N_BL<13>_XI21/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI2/MM6 N_XI21/XI2/NET35_XI21/XI2/MM6_d N_XI21/XI2/NET36_XI21/XI2/MM6_g
+ N_VSS_XI21/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI2/MM7 N_XI21/XI2/NET36_XI21/XI2/MM7_d N_XI21/XI2/NET35_XI21/XI2/MM7_g
+ N_VSS_XI21/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI2/MM8 N_XI21/XI2/NET35_XI21/XI2/MM8_d N_WL<39>_XI21/XI2/MM8_g
+ N_BLN<13>_XI21/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI2/MM5 N_XI21/XI2/NET34_XI21/XI2/MM5_d N_XI21/XI2/NET33_XI21/XI2/MM5_g
+ N_VDD_XI21/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI2/MM4 N_XI21/XI2/NET33_XI21/XI2/MM4_d N_XI21/XI2/NET34_XI21/XI2/MM4_g
+ N_VDD_XI21/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI2/MM10 N_XI21/XI2/NET35_XI21/XI2/MM10_d N_XI21/XI2/NET36_XI21/XI2/MM10_g
+ N_VDD_XI21/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI2/MM11 N_XI21/XI2/NET36_XI21/XI2/MM11_d N_XI21/XI2/NET35_XI21/XI2/MM11_g
+ N_VDD_XI21/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI3/MM2 N_XI21/XI3/NET34_XI21/XI3/MM2_d N_XI21/XI3/NET33_XI21/XI3/MM2_g
+ N_VSS_XI21/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI3/MM3 N_XI21/XI3/NET33_XI21/XI3/MM3_d N_WL<38>_XI21/XI3/MM3_g
+ N_BLN<12>_XI21/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI3/MM0 N_XI21/XI3/NET34_XI21/XI3/MM0_d N_WL<38>_XI21/XI3/MM0_g
+ N_BL<12>_XI21/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI3/MM1 N_XI21/XI3/NET33_XI21/XI3/MM1_d N_XI21/XI3/NET34_XI21/XI3/MM1_g
+ N_VSS_XI21/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI3/MM9 N_XI21/XI3/NET36_XI21/XI3/MM9_d N_WL<39>_XI21/XI3/MM9_g
+ N_BL<12>_XI21/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI3/MM6 N_XI21/XI3/NET35_XI21/XI3/MM6_d N_XI21/XI3/NET36_XI21/XI3/MM6_g
+ N_VSS_XI21/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI3/MM7 N_XI21/XI3/NET36_XI21/XI3/MM7_d N_XI21/XI3/NET35_XI21/XI3/MM7_g
+ N_VSS_XI21/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI3/MM8 N_XI21/XI3/NET35_XI21/XI3/MM8_d N_WL<39>_XI21/XI3/MM8_g
+ N_BLN<12>_XI21/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI3/MM5 N_XI21/XI3/NET34_XI21/XI3/MM5_d N_XI21/XI3/NET33_XI21/XI3/MM5_g
+ N_VDD_XI21/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI3/MM4 N_XI21/XI3/NET33_XI21/XI3/MM4_d N_XI21/XI3/NET34_XI21/XI3/MM4_g
+ N_VDD_XI21/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI3/MM10 N_XI21/XI3/NET35_XI21/XI3/MM10_d N_XI21/XI3/NET36_XI21/XI3/MM10_g
+ N_VDD_XI21/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI3/MM11 N_XI21/XI3/NET36_XI21/XI3/MM11_d N_XI21/XI3/NET35_XI21/XI3/MM11_g
+ N_VDD_XI21/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI4/MM2 N_XI21/XI4/NET34_XI21/XI4/MM2_d N_XI21/XI4/NET33_XI21/XI4/MM2_g
+ N_VSS_XI21/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI4/MM3 N_XI21/XI4/NET33_XI21/XI4/MM3_d N_WL<38>_XI21/XI4/MM3_g
+ N_BLN<11>_XI21/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI4/MM0 N_XI21/XI4/NET34_XI21/XI4/MM0_d N_WL<38>_XI21/XI4/MM0_g
+ N_BL<11>_XI21/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI4/MM1 N_XI21/XI4/NET33_XI21/XI4/MM1_d N_XI21/XI4/NET34_XI21/XI4/MM1_g
+ N_VSS_XI21/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI4/MM9 N_XI21/XI4/NET36_XI21/XI4/MM9_d N_WL<39>_XI21/XI4/MM9_g
+ N_BL<11>_XI21/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI4/MM6 N_XI21/XI4/NET35_XI21/XI4/MM6_d N_XI21/XI4/NET36_XI21/XI4/MM6_g
+ N_VSS_XI21/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI4/MM7 N_XI21/XI4/NET36_XI21/XI4/MM7_d N_XI21/XI4/NET35_XI21/XI4/MM7_g
+ N_VSS_XI21/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI4/MM8 N_XI21/XI4/NET35_XI21/XI4/MM8_d N_WL<39>_XI21/XI4/MM8_g
+ N_BLN<11>_XI21/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI4/MM5 N_XI21/XI4/NET34_XI21/XI4/MM5_d N_XI21/XI4/NET33_XI21/XI4/MM5_g
+ N_VDD_XI21/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI4/MM4 N_XI21/XI4/NET33_XI21/XI4/MM4_d N_XI21/XI4/NET34_XI21/XI4/MM4_g
+ N_VDD_XI21/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI4/MM10 N_XI21/XI4/NET35_XI21/XI4/MM10_d N_XI21/XI4/NET36_XI21/XI4/MM10_g
+ N_VDD_XI21/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI4/MM11 N_XI21/XI4/NET36_XI21/XI4/MM11_d N_XI21/XI4/NET35_XI21/XI4/MM11_g
+ N_VDD_XI21/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI5/MM2 N_XI21/XI5/NET34_XI21/XI5/MM2_d N_XI21/XI5/NET33_XI21/XI5/MM2_g
+ N_VSS_XI21/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI5/MM3 N_XI21/XI5/NET33_XI21/XI5/MM3_d N_WL<38>_XI21/XI5/MM3_g
+ N_BLN<10>_XI21/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI5/MM0 N_XI21/XI5/NET34_XI21/XI5/MM0_d N_WL<38>_XI21/XI5/MM0_g
+ N_BL<10>_XI21/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI5/MM1 N_XI21/XI5/NET33_XI21/XI5/MM1_d N_XI21/XI5/NET34_XI21/XI5/MM1_g
+ N_VSS_XI21/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI5/MM9 N_XI21/XI5/NET36_XI21/XI5/MM9_d N_WL<39>_XI21/XI5/MM9_g
+ N_BL<10>_XI21/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI5/MM6 N_XI21/XI5/NET35_XI21/XI5/MM6_d N_XI21/XI5/NET36_XI21/XI5/MM6_g
+ N_VSS_XI21/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI5/MM7 N_XI21/XI5/NET36_XI21/XI5/MM7_d N_XI21/XI5/NET35_XI21/XI5/MM7_g
+ N_VSS_XI21/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI5/MM8 N_XI21/XI5/NET35_XI21/XI5/MM8_d N_WL<39>_XI21/XI5/MM8_g
+ N_BLN<10>_XI21/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI5/MM5 N_XI21/XI5/NET34_XI21/XI5/MM5_d N_XI21/XI5/NET33_XI21/XI5/MM5_g
+ N_VDD_XI21/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI5/MM4 N_XI21/XI5/NET33_XI21/XI5/MM4_d N_XI21/XI5/NET34_XI21/XI5/MM4_g
+ N_VDD_XI21/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI5/MM10 N_XI21/XI5/NET35_XI21/XI5/MM10_d N_XI21/XI5/NET36_XI21/XI5/MM10_g
+ N_VDD_XI21/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI5/MM11 N_XI21/XI5/NET36_XI21/XI5/MM11_d N_XI21/XI5/NET35_XI21/XI5/MM11_g
+ N_VDD_XI21/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI6/MM2 N_XI21/XI6/NET34_XI21/XI6/MM2_d N_XI21/XI6/NET33_XI21/XI6/MM2_g
+ N_VSS_XI21/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM3 N_XI21/XI6/NET33_XI21/XI6/MM3_d N_WL<38>_XI21/XI6/MM3_g
+ N_BLN<9>_XI21/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM0 N_XI21/XI6/NET34_XI21/XI6/MM0_d N_WL<38>_XI21/XI6/MM0_g
+ N_BL<9>_XI21/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM1 N_XI21/XI6/NET33_XI21/XI6/MM1_d N_XI21/XI6/NET34_XI21/XI6/MM1_g
+ N_VSS_XI21/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM9 N_XI21/XI6/NET36_XI21/XI6/MM9_d N_WL<39>_XI21/XI6/MM9_g
+ N_BL<9>_XI21/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM6 N_XI21/XI6/NET35_XI21/XI6/MM6_d N_XI21/XI6/NET36_XI21/XI6/MM6_g
+ N_VSS_XI21/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM7 N_XI21/XI6/NET36_XI21/XI6/MM7_d N_XI21/XI6/NET35_XI21/XI6/MM7_g
+ N_VSS_XI21/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM8 N_XI21/XI6/NET35_XI21/XI6/MM8_d N_WL<39>_XI21/XI6/MM8_g
+ N_BLN<9>_XI21/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI6/MM5 N_XI21/XI6/NET34_XI21/XI6/MM5_d N_XI21/XI6/NET33_XI21/XI6/MM5_g
+ N_VDD_XI21/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI6/MM4 N_XI21/XI6/NET33_XI21/XI6/MM4_d N_XI21/XI6/NET34_XI21/XI6/MM4_g
+ N_VDD_XI21/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI6/MM10 N_XI21/XI6/NET35_XI21/XI6/MM10_d N_XI21/XI6/NET36_XI21/XI6/MM10_g
+ N_VDD_XI21/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI6/MM11 N_XI21/XI6/NET36_XI21/XI6/MM11_d N_XI21/XI6/NET35_XI21/XI6/MM11_g
+ N_VDD_XI21/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI7/MM2 N_XI21/XI7/NET34_XI21/XI7/MM2_d N_XI21/XI7/NET33_XI21/XI7/MM2_g
+ N_VSS_XI21/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM3 N_XI21/XI7/NET33_XI21/XI7/MM3_d N_WL<38>_XI21/XI7/MM3_g
+ N_BLN<8>_XI21/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM0 N_XI21/XI7/NET34_XI21/XI7/MM0_d N_WL<38>_XI21/XI7/MM0_g
+ N_BL<8>_XI21/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM1 N_XI21/XI7/NET33_XI21/XI7/MM1_d N_XI21/XI7/NET34_XI21/XI7/MM1_g
+ N_VSS_XI21/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM9 N_XI21/XI7/NET36_XI21/XI7/MM9_d N_WL<39>_XI21/XI7/MM9_g
+ N_BL<8>_XI21/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM6 N_XI21/XI7/NET35_XI21/XI7/MM6_d N_XI21/XI7/NET36_XI21/XI7/MM6_g
+ N_VSS_XI21/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM7 N_XI21/XI7/NET36_XI21/XI7/MM7_d N_XI21/XI7/NET35_XI21/XI7/MM7_g
+ N_VSS_XI21/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM8 N_XI21/XI7/NET35_XI21/XI7/MM8_d N_WL<39>_XI21/XI7/MM8_g
+ N_BLN<8>_XI21/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI7/MM5 N_XI21/XI7/NET34_XI21/XI7/MM5_d N_XI21/XI7/NET33_XI21/XI7/MM5_g
+ N_VDD_XI21/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI7/MM4 N_XI21/XI7/NET33_XI21/XI7/MM4_d N_XI21/XI7/NET34_XI21/XI7/MM4_g
+ N_VDD_XI21/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI7/MM10 N_XI21/XI7/NET35_XI21/XI7/MM10_d N_XI21/XI7/NET36_XI21/XI7/MM10_g
+ N_VDD_XI21/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI7/MM11 N_XI21/XI7/NET36_XI21/XI7/MM11_d N_XI21/XI7/NET35_XI21/XI7/MM11_g
+ N_VDD_XI21/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI8/MM2 N_XI21/XI8/NET34_XI21/XI8/MM2_d N_XI21/XI8/NET33_XI21/XI8/MM2_g
+ N_VSS_XI21/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM3 N_XI21/XI8/NET33_XI21/XI8/MM3_d N_WL<38>_XI21/XI8/MM3_g
+ N_BLN<7>_XI21/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM0 N_XI21/XI8/NET34_XI21/XI8/MM0_d N_WL<38>_XI21/XI8/MM0_g
+ N_BL<7>_XI21/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM1 N_XI21/XI8/NET33_XI21/XI8/MM1_d N_XI21/XI8/NET34_XI21/XI8/MM1_g
+ N_VSS_XI21/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM9 N_XI21/XI8/NET36_XI21/XI8/MM9_d N_WL<39>_XI21/XI8/MM9_g
+ N_BL<7>_XI21/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM6 N_XI21/XI8/NET35_XI21/XI8/MM6_d N_XI21/XI8/NET36_XI21/XI8/MM6_g
+ N_VSS_XI21/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM7 N_XI21/XI8/NET36_XI21/XI8/MM7_d N_XI21/XI8/NET35_XI21/XI8/MM7_g
+ N_VSS_XI21/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM8 N_XI21/XI8/NET35_XI21/XI8/MM8_d N_WL<39>_XI21/XI8/MM8_g
+ N_BLN<7>_XI21/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI8/MM5 N_XI21/XI8/NET34_XI21/XI8/MM5_d N_XI21/XI8/NET33_XI21/XI8/MM5_g
+ N_VDD_XI21/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI8/MM4 N_XI21/XI8/NET33_XI21/XI8/MM4_d N_XI21/XI8/NET34_XI21/XI8/MM4_g
+ N_VDD_XI21/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI8/MM10 N_XI21/XI8/NET35_XI21/XI8/MM10_d N_XI21/XI8/NET36_XI21/XI8/MM10_g
+ N_VDD_XI21/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI8/MM11 N_XI21/XI8/NET36_XI21/XI8/MM11_d N_XI21/XI8/NET35_XI21/XI8/MM11_g
+ N_VDD_XI21/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI9/MM2 N_XI21/XI9/NET34_XI21/XI9/MM2_d N_XI21/XI9/NET33_XI21/XI9/MM2_g
+ N_VSS_XI21/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM3 N_XI21/XI9/NET33_XI21/XI9/MM3_d N_WL<38>_XI21/XI9/MM3_g
+ N_BLN<6>_XI21/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM0 N_XI21/XI9/NET34_XI21/XI9/MM0_d N_WL<38>_XI21/XI9/MM0_g
+ N_BL<6>_XI21/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM1 N_XI21/XI9/NET33_XI21/XI9/MM1_d N_XI21/XI9/NET34_XI21/XI9/MM1_g
+ N_VSS_XI21/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM9 N_XI21/XI9/NET36_XI21/XI9/MM9_d N_WL<39>_XI21/XI9/MM9_g
+ N_BL<6>_XI21/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM6 N_XI21/XI9/NET35_XI21/XI9/MM6_d N_XI21/XI9/NET36_XI21/XI9/MM6_g
+ N_VSS_XI21/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM7 N_XI21/XI9/NET36_XI21/XI9/MM7_d N_XI21/XI9/NET35_XI21/XI9/MM7_g
+ N_VSS_XI21/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM8 N_XI21/XI9/NET35_XI21/XI9/MM8_d N_WL<39>_XI21/XI9/MM8_g
+ N_BLN<6>_XI21/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI9/MM5 N_XI21/XI9/NET34_XI21/XI9/MM5_d N_XI21/XI9/NET33_XI21/XI9/MM5_g
+ N_VDD_XI21/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI9/MM4 N_XI21/XI9/NET33_XI21/XI9/MM4_d N_XI21/XI9/NET34_XI21/XI9/MM4_g
+ N_VDD_XI21/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI9/MM10 N_XI21/XI9/NET35_XI21/XI9/MM10_d N_XI21/XI9/NET36_XI21/XI9/MM10_g
+ N_VDD_XI21/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI9/MM11 N_XI21/XI9/NET36_XI21/XI9/MM11_d N_XI21/XI9/NET35_XI21/XI9/MM11_g
+ N_VDD_XI21/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI10/MM2 N_XI21/XI10/NET34_XI21/XI10/MM2_d
+ N_XI21/XI10/NET33_XI21/XI10/MM2_g N_VSS_XI21/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI10/MM3 N_XI21/XI10/NET33_XI21/XI10/MM3_d N_WL<38>_XI21/XI10/MM3_g
+ N_BLN<5>_XI21/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI10/MM0 N_XI21/XI10/NET34_XI21/XI10/MM0_d N_WL<38>_XI21/XI10/MM0_g
+ N_BL<5>_XI21/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI10/MM1 N_XI21/XI10/NET33_XI21/XI10/MM1_d
+ N_XI21/XI10/NET34_XI21/XI10/MM1_g N_VSS_XI21/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI10/MM9 N_XI21/XI10/NET36_XI21/XI10/MM9_d N_WL<39>_XI21/XI10/MM9_g
+ N_BL<5>_XI21/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI10/MM6 N_XI21/XI10/NET35_XI21/XI10/MM6_d
+ N_XI21/XI10/NET36_XI21/XI10/MM6_g N_VSS_XI21/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI10/MM7 N_XI21/XI10/NET36_XI21/XI10/MM7_d
+ N_XI21/XI10/NET35_XI21/XI10/MM7_g N_VSS_XI21/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI10/MM8 N_XI21/XI10/NET35_XI21/XI10/MM8_d N_WL<39>_XI21/XI10/MM8_g
+ N_BLN<5>_XI21/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI10/MM5 N_XI21/XI10/NET34_XI21/XI10/MM5_d
+ N_XI21/XI10/NET33_XI21/XI10/MM5_g N_VDD_XI21/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI10/MM4 N_XI21/XI10/NET33_XI21/XI10/MM4_d
+ N_XI21/XI10/NET34_XI21/XI10/MM4_g N_VDD_XI21/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI10/MM10 N_XI21/XI10/NET35_XI21/XI10/MM10_d
+ N_XI21/XI10/NET36_XI21/XI10/MM10_g N_VDD_XI21/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI10/MM11 N_XI21/XI10/NET36_XI21/XI10/MM11_d
+ N_XI21/XI10/NET35_XI21/XI10/MM11_g N_VDD_XI21/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI11/MM2 N_XI21/XI11/NET34_XI21/XI11/MM2_d
+ N_XI21/XI11/NET33_XI21/XI11/MM2_g N_VSS_XI21/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI11/MM3 N_XI21/XI11/NET33_XI21/XI11/MM3_d N_WL<38>_XI21/XI11/MM3_g
+ N_BLN<4>_XI21/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI11/MM0 N_XI21/XI11/NET34_XI21/XI11/MM0_d N_WL<38>_XI21/XI11/MM0_g
+ N_BL<4>_XI21/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI11/MM1 N_XI21/XI11/NET33_XI21/XI11/MM1_d
+ N_XI21/XI11/NET34_XI21/XI11/MM1_g N_VSS_XI21/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI11/MM9 N_XI21/XI11/NET36_XI21/XI11/MM9_d N_WL<39>_XI21/XI11/MM9_g
+ N_BL<4>_XI21/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI11/MM6 N_XI21/XI11/NET35_XI21/XI11/MM6_d
+ N_XI21/XI11/NET36_XI21/XI11/MM6_g N_VSS_XI21/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI11/MM7 N_XI21/XI11/NET36_XI21/XI11/MM7_d
+ N_XI21/XI11/NET35_XI21/XI11/MM7_g N_VSS_XI21/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI11/MM8 N_XI21/XI11/NET35_XI21/XI11/MM8_d N_WL<39>_XI21/XI11/MM8_g
+ N_BLN<4>_XI21/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI11/MM5 N_XI21/XI11/NET34_XI21/XI11/MM5_d
+ N_XI21/XI11/NET33_XI21/XI11/MM5_g N_VDD_XI21/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI11/MM4 N_XI21/XI11/NET33_XI21/XI11/MM4_d
+ N_XI21/XI11/NET34_XI21/XI11/MM4_g N_VDD_XI21/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI11/MM10 N_XI21/XI11/NET35_XI21/XI11/MM10_d
+ N_XI21/XI11/NET36_XI21/XI11/MM10_g N_VDD_XI21/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI11/MM11 N_XI21/XI11/NET36_XI21/XI11/MM11_d
+ N_XI21/XI11/NET35_XI21/XI11/MM11_g N_VDD_XI21/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI12/MM2 N_XI21/XI12/NET34_XI21/XI12/MM2_d
+ N_XI21/XI12/NET33_XI21/XI12/MM2_g N_VSS_XI21/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI12/MM3 N_XI21/XI12/NET33_XI21/XI12/MM3_d N_WL<38>_XI21/XI12/MM3_g
+ N_BLN<3>_XI21/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI12/MM0 N_XI21/XI12/NET34_XI21/XI12/MM0_d N_WL<38>_XI21/XI12/MM0_g
+ N_BL<3>_XI21/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI12/MM1 N_XI21/XI12/NET33_XI21/XI12/MM1_d
+ N_XI21/XI12/NET34_XI21/XI12/MM1_g N_VSS_XI21/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI12/MM9 N_XI21/XI12/NET36_XI21/XI12/MM9_d N_WL<39>_XI21/XI12/MM9_g
+ N_BL<3>_XI21/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI12/MM6 N_XI21/XI12/NET35_XI21/XI12/MM6_d
+ N_XI21/XI12/NET36_XI21/XI12/MM6_g N_VSS_XI21/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI12/MM7 N_XI21/XI12/NET36_XI21/XI12/MM7_d
+ N_XI21/XI12/NET35_XI21/XI12/MM7_g N_VSS_XI21/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI12/MM8 N_XI21/XI12/NET35_XI21/XI12/MM8_d N_WL<39>_XI21/XI12/MM8_g
+ N_BLN<3>_XI21/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI12/MM5 N_XI21/XI12/NET34_XI21/XI12/MM5_d
+ N_XI21/XI12/NET33_XI21/XI12/MM5_g N_VDD_XI21/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI12/MM4 N_XI21/XI12/NET33_XI21/XI12/MM4_d
+ N_XI21/XI12/NET34_XI21/XI12/MM4_g N_VDD_XI21/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI12/MM10 N_XI21/XI12/NET35_XI21/XI12/MM10_d
+ N_XI21/XI12/NET36_XI21/XI12/MM10_g N_VDD_XI21/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI12/MM11 N_XI21/XI12/NET36_XI21/XI12/MM11_d
+ N_XI21/XI12/NET35_XI21/XI12/MM11_g N_VDD_XI21/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI13/MM2 N_XI21/XI13/NET34_XI21/XI13/MM2_d
+ N_XI21/XI13/NET33_XI21/XI13/MM2_g N_VSS_XI21/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI13/MM3 N_XI21/XI13/NET33_XI21/XI13/MM3_d N_WL<38>_XI21/XI13/MM3_g
+ N_BLN<2>_XI21/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI13/MM0 N_XI21/XI13/NET34_XI21/XI13/MM0_d N_WL<38>_XI21/XI13/MM0_g
+ N_BL<2>_XI21/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI13/MM1 N_XI21/XI13/NET33_XI21/XI13/MM1_d
+ N_XI21/XI13/NET34_XI21/XI13/MM1_g N_VSS_XI21/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI13/MM9 N_XI21/XI13/NET36_XI21/XI13/MM9_d N_WL<39>_XI21/XI13/MM9_g
+ N_BL<2>_XI21/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI13/MM6 N_XI21/XI13/NET35_XI21/XI13/MM6_d
+ N_XI21/XI13/NET36_XI21/XI13/MM6_g N_VSS_XI21/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI13/MM7 N_XI21/XI13/NET36_XI21/XI13/MM7_d
+ N_XI21/XI13/NET35_XI21/XI13/MM7_g N_VSS_XI21/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI13/MM8 N_XI21/XI13/NET35_XI21/XI13/MM8_d N_WL<39>_XI21/XI13/MM8_g
+ N_BLN<2>_XI21/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI13/MM5 N_XI21/XI13/NET34_XI21/XI13/MM5_d
+ N_XI21/XI13/NET33_XI21/XI13/MM5_g N_VDD_XI21/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI13/MM4 N_XI21/XI13/NET33_XI21/XI13/MM4_d
+ N_XI21/XI13/NET34_XI21/XI13/MM4_g N_VDD_XI21/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI13/MM10 N_XI21/XI13/NET35_XI21/XI13/MM10_d
+ N_XI21/XI13/NET36_XI21/XI13/MM10_g N_VDD_XI21/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI13/MM11 N_XI21/XI13/NET36_XI21/XI13/MM11_d
+ N_XI21/XI13/NET35_XI21/XI13/MM11_g N_VDD_XI21/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI14/MM2 N_XI21/XI14/NET34_XI21/XI14/MM2_d
+ N_XI21/XI14/NET33_XI21/XI14/MM2_g N_VSS_XI21/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI14/MM3 N_XI21/XI14/NET33_XI21/XI14/MM3_d N_WL<38>_XI21/XI14/MM3_g
+ N_BLN<1>_XI21/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI14/MM0 N_XI21/XI14/NET34_XI21/XI14/MM0_d N_WL<38>_XI21/XI14/MM0_g
+ N_BL<1>_XI21/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI14/MM1 N_XI21/XI14/NET33_XI21/XI14/MM1_d
+ N_XI21/XI14/NET34_XI21/XI14/MM1_g N_VSS_XI21/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI14/MM9 N_XI21/XI14/NET36_XI21/XI14/MM9_d N_WL<39>_XI21/XI14/MM9_g
+ N_BL<1>_XI21/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI14/MM6 N_XI21/XI14/NET35_XI21/XI14/MM6_d
+ N_XI21/XI14/NET36_XI21/XI14/MM6_g N_VSS_XI21/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI14/MM7 N_XI21/XI14/NET36_XI21/XI14/MM7_d
+ N_XI21/XI14/NET35_XI21/XI14/MM7_g N_VSS_XI21/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI14/MM8 N_XI21/XI14/NET35_XI21/XI14/MM8_d N_WL<39>_XI21/XI14/MM8_g
+ N_BLN<1>_XI21/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI14/MM5 N_XI21/XI14/NET34_XI21/XI14/MM5_d
+ N_XI21/XI14/NET33_XI21/XI14/MM5_g N_VDD_XI21/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI14/MM4 N_XI21/XI14/NET33_XI21/XI14/MM4_d
+ N_XI21/XI14/NET34_XI21/XI14/MM4_g N_VDD_XI21/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI14/MM10 N_XI21/XI14/NET35_XI21/XI14/MM10_d
+ N_XI21/XI14/NET36_XI21/XI14/MM10_g N_VDD_XI21/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI14/MM11 N_XI21/XI14/NET36_XI21/XI14/MM11_d
+ N_XI21/XI14/NET35_XI21/XI14/MM11_g N_VDD_XI21/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI15/MM2 N_XI21/XI15/NET34_XI21/XI15/MM2_d
+ N_XI21/XI15/NET33_XI21/XI15/MM2_g N_VSS_XI21/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI15/MM3 N_XI21/XI15/NET33_XI21/XI15/MM3_d N_WL<38>_XI21/XI15/MM3_g
+ N_BLN<0>_XI21/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI15/MM0 N_XI21/XI15/NET34_XI21/XI15/MM0_d N_WL<38>_XI21/XI15/MM0_g
+ N_BL<0>_XI21/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI15/MM1 N_XI21/XI15/NET33_XI21/XI15/MM1_d
+ N_XI21/XI15/NET34_XI21/XI15/MM1_g N_VSS_XI21/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI15/MM9 N_XI21/XI15/NET36_XI21/XI15/MM9_d N_WL<39>_XI21/XI15/MM9_g
+ N_BL<0>_XI21/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI15/MM6 N_XI21/XI15/NET35_XI21/XI15/MM6_d
+ N_XI21/XI15/NET36_XI21/XI15/MM6_g N_VSS_XI21/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI15/MM7 N_XI21/XI15/NET36_XI21/XI15/MM7_d
+ N_XI21/XI15/NET35_XI21/XI15/MM7_g N_VSS_XI21/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI21/XI15/MM8 N_XI21/XI15/NET35_XI21/XI15/MM8_d N_WL<39>_XI21/XI15/MM8_g
+ N_BLN<0>_XI21/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI21/XI15/MM5 N_XI21/XI15/NET34_XI21/XI15/MM5_d
+ N_XI21/XI15/NET33_XI21/XI15/MM5_g N_VDD_XI21/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI15/MM4 N_XI21/XI15/NET33_XI21/XI15/MM4_d
+ N_XI21/XI15/NET34_XI21/XI15/MM4_g N_VDD_XI21/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI15/MM10 N_XI21/XI15/NET35_XI21/XI15/MM10_d
+ N_XI21/XI15/NET36_XI21/XI15/MM10_g N_VDD_XI21/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI21/XI15/MM11 N_XI21/XI15/NET36_XI21/XI15/MM11_d
+ N_XI21/XI15/NET35_XI21/XI15/MM11_g N_VDD_XI21/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI0/MM2 N_XI22/XI0/NET34_XI22/XI0/MM2_d N_XI22/XI0/NET33_XI22/XI0/MM2_g
+ N_VSS_XI22/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI0/MM3 N_XI22/XI0/NET33_XI22/XI0/MM3_d N_WL<40>_XI22/XI0/MM3_g
+ N_BLN<15>_XI22/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI0/MM0 N_XI22/XI0/NET34_XI22/XI0/MM0_d N_WL<40>_XI22/XI0/MM0_g
+ N_BL<15>_XI22/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI0/MM1 N_XI22/XI0/NET33_XI22/XI0/MM1_d N_XI22/XI0/NET34_XI22/XI0/MM1_g
+ N_VSS_XI22/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI0/MM9 N_XI22/XI0/NET36_XI22/XI0/MM9_d N_WL<41>_XI22/XI0/MM9_g
+ N_BL<15>_XI22/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI0/MM6 N_XI22/XI0/NET35_XI22/XI0/MM6_d N_XI22/XI0/NET36_XI22/XI0/MM6_g
+ N_VSS_XI22/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI0/MM7 N_XI22/XI0/NET36_XI22/XI0/MM7_d N_XI22/XI0/NET35_XI22/XI0/MM7_g
+ N_VSS_XI22/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI0/MM8 N_XI22/XI0/NET35_XI22/XI0/MM8_d N_WL<41>_XI22/XI0/MM8_g
+ N_BLN<15>_XI22/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI0/MM5 N_XI22/XI0/NET34_XI22/XI0/MM5_d N_XI22/XI0/NET33_XI22/XI0/MM5_g
+ N_VDD_XI22/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI0/MM4 N_XI22/XI0/NET33_XI22/XI0/MM4_d N_XI22/XI0/NET34_XI22/XI0/MM4_g
+ N_VDD_XI22/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI0/MM10 N_XI22/XI0/NET35_XI22/XI0/MM10_d N_XI22/XI0/NET36_XI22/XI0/MM10_g
+ N_VDD_XI22/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI0/MM11 N_XI22/XI0/NET36_XI22/XI0/MM11_d N_XI22/XI0/NET35_XI22/XI0/MM11_g
+ N_VDD_XI22/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI1/MM2 N_XI22/XI1/NET34_XI22/XI1/MM2_d N_XI22/XI1/NET33_XI22/XI1/MM2_g
+ N_VSS_XI22/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI1/MM3 N_XI22/XI1/NET33_XI22/XI1/MM3_d N_WL<40>_XI22/XI1/MM3_g
+ N_BLN<14>_XI22/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI1/MM0 N_XI22/XI1/NET34_XI22/XI1/MM0_d N_WL<40>_XI22/XI1/MM0_g
+ N_BL<14>_XI22/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI1/MM1 N_XI22/XI1/NET33_XI22/XI1/MM1_d N_XI22/XI1/NET34_XI22/XI1/MM1_g
+ N_VSS_XI22/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI1/MM9 N_XI22/XI1/NET36_XI22/XI1/MM9_d N_WL<41>_XI22/XI1/MM9_g
+ N_BL<14>_XI22/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI1/MM6 N_XI22/XI1/NET35_XI22/XI1/MM6_d N_XI22/XI1/NET36_XI22/XI1/MM6_g
+ N_VSS_XI22/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI1/MM7 N_XI22/XI1/NET36_XI22/XI1/MM7_d N_XI22/XI1/NET35_XI22/XI1/MM7_g
+ N_VSS_XI22/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI1/MM8 N_XI22/XI1/NET35_XI22/XI1/MM8_d N_WL<41>_XI22/XI1/MM8_g
+ N_BLN<14>_XI22/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI1/MM5 N_XI22/XI1/NET34_XI22/XI1/MM5_d N_XI22/XI1/NET33_XI22/XI1/MM5_g
+ N_VDD_XI22/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI1/MM4 N_XI22/XI1/NET33_XI22/XI1/MM4_d N_XI22/XI1/NET34_XI22/XI1/MM4_g
+ N_VDD_XI22/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI1/MM10 N_XI22/XI1/NET35_XI22/XI1/MM10_d N_XI22/XI1/NET36_XI22/XI1/MM10_g
+ N_VDD_XI22/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI1/MM11 N_XI22/XI1/NET36_XI22/XI1/MM11_d N_XI22/XI1/NET35_XI22/XI1/MM11_g
+ N_VDD_XI22/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI2/MM2 N_XI22/XI2/NET34_XI22/XI2/MM2_d N_XI22/XI2/NET33_XI22/XI2/MM2_g
+ N_VSS_XI22/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI2/MM3 N_XI22/XI2/NET33_XI22/XI2/MM3_d N_WL<40>_XI22/XI2/MM3_g
+ N_BLN<13>_XI22/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI2/MM0 N_XI22/XI2/NET34_XI22/XI2/MM0_d N_WL<40>_XI22/XI2/MM0_g
+ N_BL<13>_XI22/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI2/MM1 N_XI22/XI2/NET33_XI22/XI2/MM1_d N_XI22/XI2/NET34_XI22/XI2/MM1_g
+ N_VSS_XI22/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI2/MM9 N_XI22/XI2/NET36_XI22/XI2/MM9_d N_WL<41>_XI22/XI2/MM9_g
+ N_BL<13>_XI22/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI2/MM6 N_XI22/XI2/NET35_XI22/XI2/MM6_d N_XI22/XI2/NET36_XI22/XI2/MM6_g
+ N_VSS_XI22/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI2/MM7 N_XI22/XI2/NET36_XI22/XI2/MM7_d N_XI22/XI2/NET35_XI22/XI2/MM7_g
+ N_VSS_XI22/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI2/MM8 N_XI22/XI2/NET35_XI22/XI2/MM8_d N_WL<41>_XI22/XI2/MM8_g
+ N_BLN<13>_XI22/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI2/MM5 N_XI22/XI2/NET34_XI22/XI2/MM5_d N_XI22/XI2/NET33_XI22/XI2/MM5_g
+ N_VDD_XI22/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI2/MM4 N_XI22/XI2/NET33_XI22/XI2/MM4_d N_XI22/XI2/NET34_XI22/XI2/MM4_g
+ N_VDD_XI22/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI2/MM10 N_XI22/XI2/NET35_XI22/XI2/MM10_d N_XI22/XI2/NET36_XI22/XI2/MM10_g
+ N_VDD_XI22/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI2/MM11 N_XI22/XI2/NET36_XI22/XI2/MM11_d N_XI22/XI2/NET35_XI22/XI2/MM11_g
+ N_VDD_XI22/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI3/MM2 N_XI22/XI3/NET34_XI22/XI3/MM2_d N_XI22/XI3/NET33_XI22/XI3/MM2_g
+ N_VSS_XI22/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI3/MM3 N_XI22/XI3/NET33_XI22/XI3/MM3_d N_WL<40>_XI22/XI3/MM3_g
+ N_BLN<12>_XI22/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI3/MM0 N_XI22/XI3/NET34_XI22/XI3/MM0_d N_WL<40>_XI22/XI3/MM0_g
+ N_BL<12>_XI22/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI3/MM1 N_XI22/XI3/NET33_XI22/XI3/MM1_d N_XI22/XI3/NET34_XI22/XI3/MM1_g
+ N_VSS_XI22/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI3/MM9 N_XI22/XI3/NET36_XI22/XI3/MM9_d N_WL<41>_XI22/XI3/MM9_g
+ N_BL<12>_XI22/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI3/MM6 N_XI22/XI3/NET35_XI22/XI3/MM6_d N_XI22/XI3/NET36_XI22/XI3/MM6_g
+ N_VSS_XI22/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI3/MM7 N_XI22/XI3/NET36_XI22/XI3/MM7_d N_XI22/XI3/NET35_XI22/XI3/MM7_g
+ N_VSS_XI22/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI3/MM8 N_XI22/XI3/NET35_XI22/XI3/MM8_d N_WL<41>_XI22/XI3/MM8_g
+ N_BLN<12>_XI22/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI3/MM5 N_XI22/XI3/NET34_XI22/XI3/MM5_d N_XI22/XI3/NET33_XI22/XI3/MM5_g
+ N_VDD_XI22/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI3/MM4 N_XI22/XI3/NET33_XI22/XI3/MM4_d N_XI22/XI3/NET34_XI22/XI3/MM4_g
+ N_VDD_XI22/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI3/MM10 N_XI22/XI3/NET35_XI22/XI3/MM10_d N_XI22/XI3/NET36_XI22/XI3/MM10_g
+ N_VDD_XI22/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI3/MM11 N_XI22/XI3/NET36_XI22/XI3/MM11_d N_XI22/XI3/NET35_XI22/XI3/MM11_g
+ N_VDD_XI22/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI4/MM2 N_XI22/XI4/NET34_XI22/XI4/MM2_d N_XI22/XI4/NET33_XI22/XI4/MM2_g
+ N_VSS_XI22/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI4/MM3 N_XI22/XI4/NET33_XI22/XI4/MM3_d N_WL<40>_XI22/XI4/MM3_g
+ N_BLN<11>_XI22/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI4/MM0 N_XI22/XI4/NET34_XI22/XI4/MM0_d N_WL<40>_XI22/XI4/MM0_g
+ N_BL<11>_XI22/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI4/MM1 N_XI22/XI4/NET33_XI22/XI4/MM1_d N_XI22/XI4/NET34_XI22/XI4/MM1_g
+ N_VSS_XI22/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI4/MM9 N_XI22/XI4/NET36_XI22/XI4/MM9_d N_WL<41>_XI22/XI4/MM9_g
+ N_BL<11>_XI22/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI4/MM6 N_XI22/XI4/NET35_XI22/XI4/MM6_d N_XI22/XI4/NET36_XI22/XI4/MM6_g
+ N_VSS_XI22/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI4/MM7 N_XI22/XI4/NET36_XI22/XI4/MM7_d N_XI22/XI4/NET35_XI22/XI4/MM7_g
+ N_VSS_XI22/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI4/MM8 N_XI22/XI4/NET35_XI22/XI4/MM8_d N_WL<41>_XI22/XI4/MM8_g
+ N_BLN<11>_XI22/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI4/MM5 N_XI22/XI4/NET34_XI22/XI4/MM5_d N_XI22/XI4/NET33_XI22/XI4/MM5_g
+ N_VDD_XI22/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI4/MM4 N_XI22/XI4/NET33_XI22/XI4/MM4_d N_XI22/XI4/NET34_XI22/XI4/MM4_g
+ N_VDD_XI22/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI4/MM10 N_XI22/XI4/NET35_XI22/XI4/MM10_d N_XI22/XI4/NET36_XI22/XI4/MM10_g
+ N_VDD_XI22/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI4/MM11 N_XI22/XI4/NET36_XI22/XI4/MM11_d N_XI22/XI4/NET35_XI22/XI4/MM11_g
+ N_VDD_XI22/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI5/MM2 N_XI22/XI5/NET34_XI22/XI5/MM2_d N_XI22/XI5/NET33_XI22/XI5/MM2_g
+ N_VSS_XI22/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI5/MM3 N_XI22/XI5/NET33_XI22/XI5/MM3_d N_WL<40>_XI22/XI5/MM3_g
+ N_BLN<10>_XI22/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI5/MM0 N_XI22/XI5/NET34_XI22/XI5/MM0_d N_WL<40>_XI22/XI5/MM0_g
+ N_BL<10>_XI22/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI5/MM1 N_XI22/XI5/NET33_XI22/XI5/MM1_d N_XI22/XI5/NET34_XI22/XI5/MM1_g
+ N_VSS_XI22/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI5/MM9 N_XI22/XI5/NET36_XI22/XI5/MM9_d N_WL<41>_XI22/XI5/MM9_g
+ N_BL<10>_XI22/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI5/MM6 N_XI22/XI5/NET35_XI22/XI5/MM6_d N_XI22/XI5/NET36_XI22/XI5/MM6_g
+ N_VSS_XI22/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI5/MM7 N_XI22/XI5/NET36_XI22/XI5/MM7_d N_XI22/XI5/NET35_XI22/XI5/MM7_g
+ N_VSS_XI22/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI5/MM8 N_XI22/XI5/NET35_XI22/XI5/MM8_d N_WL<41>_XI22/XI5/MM8_g
+ N_BLN<10>_XI22/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI5/MM5 N_XI22/XI5/NET34_XI22/XI5/MM5_d N_XI22/XI5/NET33_XI22/XI5/MM5_g
+ N_VDD_XI22/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI5/MM4 N_XI22/XI5/NET33_XI22/XI5/MM4_d N_XI22/XI5/NET34_XI22/XI5/MM4_g
+ N_VDD_XI22/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI5/MM10 N_XI22/XI5/NET35_XI22/XI5/MM10_d N_XI22/XI5/NET36_XI22/XI5/MM10_g
+ N_VDD_XI22/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI5/MM11 N_XI22/XI5/NET36_XI22/XI5/MM11_d N_XI22/XI5/NET35_XI22/XI5/MM11_g
+ N_VDD_XI22/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI6/MM2 N_XI22/XI6/NET34_XI22/XI6/MM2_d N_XI22/XI6/NET33_XI22/XI6/MM2_g
+ N_VSS_XI22/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM3 N_XI22/XI6/NET33_XI22/XI6/MM3_d N_WL<40>_XI22/XI6/MM3_g
+ N_BLN<9>_XI22/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM0 N_XI22/XI6/NET34_XI22/XI6/MM0_d N_WL<40>_XI22/XI6/MM0_g
+ N_BL<9>_XI22/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM1 N_XI22/XI6/NET33_XI22/XI6/MM1_d N_XI22/XI6/NET34_XI22/XI6/MM1_g
+ N_VSS_XI22/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM9 N_XI22/XI6/NET36_XI22/XI6/MM9_d N_WL<41>_XI22/XI6/MM9_g
+ N_BL<9>_XI22/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM6 N_XI22/XI6/NET35_XI22/XI6/MM6_d N_XI22/XI6/NET36_XI22/XI6/MM6_g
+ N_VSS_XI22/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM7 N_XI22/XI6/NET36_XI22/XI6/MM7_d N_XI22/XI6/NET35_XI22/XI6/MM7_g
+ N_VSS_XI22/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM8 N_XI22/XI6/NET35_XI22/XI6/MM8_d N_WL<41>_XI22/XI6/MM8_g
+ N_BLN<9>_XI22/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI6/MM5 N_XI22/XI6/NET34_XI22/XI6/MM5_d N_XI22/XI6/NET33_XI22/XI6/MM5_g
+ N_VDD_XI22/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI6/MM4 N_XI22/XI6/NET33_XI22/XI6/MM4_d N_XI22/XI6/NET34_XI22/XI6/MM4_g
+ N_VDD_XI22/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI6/MM10 N_XI22/XI6/NET35_XI22/XI6/MM10_d N_XI22/XI6/NET36_XI22/XI6/MM10_g
+ N_VDD_XI22/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI6/MM11 N_XI22/XI6/NET36_XI22/XI6/MM11_d N_XI22/XI6/NET35_XI22/XI6/MM11_g
+ N_VDD_XI22/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI7/MM2 N_XI22/XI7/NET34_XI22/XI7/MM2_d N_XI22/XI7/NET33_XI22/XI7/MM2_g
+ N_VSS_XI22/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM3 N_XI22/XI7/NET33_XI22/XI7/MM3_d N_WL<40>_XI22/XI7/MM3_g
+ N_BLN<8>_XI22/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM0 N_XI22/XI7/NET34_XI22/XI7/MM0_d N_WL<40>_XI22/XI7/MM0_g
+ N_BL<8>_XI22/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM1 N_XI22/XI7/NET33_XI22/XI7/MM1_d N_XI22/XI7/NET34_XI22/XI7/MM1_g
+ N_VSS_XI22/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM9 N_XI22/XI7/NET36_XI22/XI7/MM9_d N_WL<41>_XI22/XI7/MM9_g
+ N_BL<8>_XI22/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM6 N_XI22/XI7/NET35_XI22/XI7/MM6_d N_XI22/XI7/NET36_XI22/XI7/MM6_g
+ N_VSS_XI22/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM7 N_XI22/XI7/NET36_XI22/XI7/MM7_d N_XI22/XI7/NET35_XI22/XI7/MM7_g
+ N_VSS_XI22/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM8 N_XI22/XI7/NET35_XI22/XI7/MM8_d N_WL<41>_XI22/XI7/MM8_g
+ N_BLN<8>_XI22/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI7/MM5 N_XI22/XI7/NET34_XI22/XI7/MM5_d N_XI22/XI7/NET33_XI22/XI7/MM5_g
+ N_VDD_XI22/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI7/MM4 N_XI22/XI7/NET33_XI22/XI7/MM4_d N_XI22/XI7/NET34_XI22/XI7/MM4_g
+ N_VDD_XI22/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI7/MM10 N_XI22/XI7/NET35_XI22/XI7/MM10_d N_XI22/XI7/NET36_XI22/XI7/MM10_g
+ N_VDD_XI22/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI7/MM11 N_XI22/XI7/NET36_XI22/XI7/MM11_d N_XI22/XI7/NET35_XI22/XI7/MM11_g
+ N_VDD_XI22/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI8/MM2 N_XI22/XI8/NET34_XI22/XI8/MM2_d N_XI22/XI8/NET33_XI22/XI8/MM2_g
+ N_VSS_XI22/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM3 N_XI22/XI8/NET33_XI22/XI8/MM3_d N_WL<40>_XI22/XI8/MM3_g
+ N_BLN<7>_XI22/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM0 N_XI22/XI8/NET34_XI22/XI8/MM0_d N_WL<40>_XI22/XI8/MM0_g
+ N_BL<7>_XI22/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM1 N_XI22/XI8/NET33_XI22/XI8/MM1_d N_XI22/XI8/NET34_XI22/XI8/MM1_g
+ N_VSS_XI22/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM9 N_XI22/XI8/NET36_XI22/XI8/MM9_d N_WL<41>_XI22/XI8/MM9_g
+ N_BL<7>_XI22/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM6 N_XI22/XI8/NET35_XI22/XI8/MM6_d N_XI22/XI8/NET36_XI22/XI8/MM6_g
+ N_VSS_XI22/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM7 N_XI22/XI8/NET36_XI22/XI8/MM7_d N_XI22/XI8/NET35_XI22/XI8/MM7_g
+ N_VSS_XI22/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM8 N_XI22/XI8/NET35_XI22/XI8/MM8_d N_WL<41>_XI22/XI8/MM8_g
+ N_BLN<7>_XI22/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI8/MM5 N_XI22/XI8/NET34_XI22/XI8/MM5_d N_XI22/XI8/NET33_XI22/XI8/MM5_g
+ N_VDD_XI22/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI8/MM4 N_XI22/XI8/NET33_XI22/XI8/MM4_d N_XI22/XI8/NET34_XI22/XI8/MM4_g
+ N_VDD_XI22/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI8/MM10 N_XI22/XI8/NET35_XI22/XI8/MM10_d N_XI22/XI8/NET36_XI22/XI8/MM10_g
+ N_VDD_XI22/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI8/MM11 N_XI22/XI8/NET36_XI22/XI8/MM11_d N_XI22/XI8/NET35_XI22/XI8/MM11_g
+ N_VDD_XI22/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI9/MM2 N_XI22/XI9/NET34_XI22/XI9/MM2_d N_XI22/XI9/NET33_XI22/XI9/MM2_g
+ N_VSS_XI22/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM3 N_XI22/XI9/NET33_XI22/XI9/MM3_d N_WL<40>_XI22/XI9/MM3_g
+ N_BLN<6>_XI22/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM0 N_XI22/XI9/NET34_XI22/XI9/MM0_d N_WL<40>_XI22/XI9/MM0_g
+ N_BL<6>_XI22/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM1 N_XI22/XI9/NET33_XI22/XI9/MM1_d N_XI22/XI9/NET34_XI22/XI9/MM1_g
+ N_VSS_XI22/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM9 N_XI22/XI9/NET36_XI22/XI9/MM9_d N_WL<41>_XI22/XI9/MM9_g
+ N_BL<6>_XI22/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM6 N_XI22/XI9/NET35_XI22/XI9/MM6_d N_XI22/XI9/NET36_XI22/XI9/MM6_g
+ N_VSS_XI22/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM7 N_XI22/XI9/NET36_XI22/XI9/MM7_d N_XI22/XI9/NET35_XI22/XI9/MM7_g
+ N_VSS_XI22/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM8 N_XI22/XI9/NET35_XI22/XI9/MM8_d N_WL<41>_XI22/XI9/MM8_g
+ N_BLN<6>_XI22/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI9/MM5 N_XI22/XI9/NET34_XI22/XI9/MM5_d N_XI22/XI9/NET33_XI22/XI9/MM5_g
+ N_VDD_XI22/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI9/MM4 N_XI22/XI9/NET33_XI22/XI9/MM4_d N_XI22/XI9/NET34_XI22/XI9/MM4_g
+ N_VDD_XI22/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI9/MM10 N_XI22/XI9/NET35_XI22/XI9/MM10_d N_XI22/XI9/NET36_XI22/XI9/MM10_g
+ N_VDD_XI22/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI9/MM11 N_XI22/XI9/NET36_XI22/XI9/MM11_d N_XI22/XI9/NET35_XI22/XI9/MM11_g
+ N_VDD_XI22/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI10/MM2 N_XI22/XI10/NET34_XI22/XI10/MM2_d
+ N_XI22/XI10/NET33_XI22/XI10/MM2_g N_VSS_XI22/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI10/MM3 N_XI22/XI10/NET33_XI22/XI10/MM3_d N_WL<40>_XI22/XI10/MM3_g
+ N_BLN<5>_XI22/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI10/MM0 N_XI22/XI10/NET34_XI22/XI10/MM0_d N_WL<40>_XI22/XI10/MM0_g
+ N_BL<5>_XI22/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI10/MM1 N_XI22/XI10/NET33_XI22/XI10/MM1_d
+ N_XI22/XI10/NET34_XI22/XI10/MM1_g N_VSS_XI22/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI10/MM9 N_XI22/XI10/NET36_XI22/XI10/MM9_d N_WL<41>_XI22/XI10/MM9_g
+ N_BL<5>_XI22/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI10/MM6 N_XI22/XI10/NET35_XI22/XI10/MM6_d
+ N_XI22/XI10/NET36_XI22/XI10/MM6_g N_VSS_XI22/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI10/MM7 N_XI22/XI10/NET36_XI22/XI10/MM7_d
+ N_XI22/XI10/NET35_XI22/XI10/MM7_g N_VSS_XI22/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI10/MM8 N_XI22/XI10/NET35_XI22/XI10/MM8_d N_WL<41>_XI22/XI10/MM8_g
+ N_BLN<5>_XI22/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI10/MM5 N_XI22/XI10/NET34_XI22/XI10/MM5_d
+ N_XI22/XI10/NET33_XI22/XI10/MM5_g N_VDD_XI22/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI10/MM4 N_XI22/XI10/NET33_XI22/XI10/MM4_d
+ N_XI22/XI10/NET34_XI22/XI10/MM4_g N_VDD_XI22/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI10/MM10 N_XI22/XI10/NET35_XI22/XI10/MM10_d
+ N_XI22/XI10/NET36_XI22/XI10/MM10_g N_VDD_XI22/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI10/MM11 N_XI22/XI10/NET36_XI22/XI10/MM11_d
+ N_XI22/XI10/NET35_XI22/XI10/MM11_g N_VDD_XI22/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI11/MM2 N_XI22/XI11/NET34_XI22/XI11/MM2_d
+ N_XI22/XI11/NET33_XI22/XI11/MM2_g N_VSS_XI22/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI11/MM3 N_XI22/XI11/NET33_XI22/XI11/MM3_d N_WL<40>_XI22/XI11/MM3_g
+ N_BLN<4>_XI22/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI11/MM0 N_XI22/XI11/NET34_XI22/XI11/MM0_d N_WL<40>_XI22/XI11/MM0_g
+ N_BL<4>_XI22/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI11/MM1 N_XI22/XI11/NET33_XI22/XI11/MM1_d
+ N_XI22/XI11/NET34_XI22/XI11/MM1_g N_VSS_XI22/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI11/MM9 N_XI22/XI11/NET36_XI22/XI11/MM9_d N_WL<41>_XI22/XI11/MM9_g
+ N_BL<4>_XI22/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI11/MM6 N_XI22/XI11/NET35_XI22/XI11/MM6_d
+ N_XI22/XI11/NET36_XI22/XI11/MM6_g N_VSS_XI22/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI11/MM7 N_XI22/XI11/NET36_XI22/XI11/MM7_d
+ N_XI22/XI11/NET35_XI22/XI11/MM7_g N_VSS_XI22/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI11/MM8 N_XI22/XI11/NET35_XI22/XI11/MM8_d N_WL<41>_XI22/XI11/MM8_g
+ N_BLN<4>_XI22/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI11/MM5 N_XI22/XI11/NET34_XI22/XI11/MM5_d
+ N_XI22/XI11/NET33_XI22/XI11/MM5_g N_VDD_XI22/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI11/MM4 N_XI22/XI11/NET33_XI22/XI11/MM4_d
+ N_XI22/XI11/NET34_XI22/XI11/MM4_g N_VDD_XI22/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI11/MM10 N_XI22/XI11/NET35_XI22/XI11/MM10_d
+ N_XI22/XI11/NET36_XI22/XI11/MM10_g N_VDD_XI22/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI11/MM11 N_XI22/XI11/NET36_XI22/XI11/MM11_d
+ N_XI22/XI11/NET35_XI22/XI11/MM11_g N_VDD_XI22/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI12/MM2 N_XI22/XI12/NET34_XI22/XI12/MM2_d
+ N_XI22/XI12/NET33_XI22/XI12/MM2_g N_VSS_XI22/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI12/MM3 N_XI22/XI12/NET33_XI22/XI12/MM3_d N_WL<40>_XI22/XI12/MM3_g
+ N_BLN<3>_XI22/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI12/MM0 N_XI22/XI12/NET34_XI22/XI12/MM0_d N_WL<40>_XI22/XI12/MM0_g
+ N_BL<3>_XI22/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI12/MM1 N_XI22/XI12/NET33_XI22/XI12/MM1_d
+ N_XI22/XI12/NET34_XI22/XI12/MM1_g N_VSS_XI22/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI12/MM9 N_XI22/XI12/NET36_XI22/XI12/MM9_d N_WL<41>_XI22/XI12/MM9_g
+ N_BL<3>_XI22/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI12/MM6 N_XI22/XI12/NET35_XI22/XI12/MM6_d
+ N_XI22/XI12/NET36_XI22/XI12/MM6_g N_VSS_XI22/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI12/MM7 N_XI22/XI12/NET36_XI22/XI12/MM7_d
+ N_XI22/XI12/NET35_XI22/XI12/MM7_g N_VSS_XI22/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI12/MM8 N_XI22/XI12/NET35_XI22/XI12/MM8_d N_WL<41>_XI22/XI12/MM8_g
+ N_BLN<3>_XI22/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI12/MM5 N_XI22/XI12/NET34_XI22/XI12/MM5_d
+ N_XI22/XI12/NET33_XI22/XI12/MM5_g N_VDD_XI22/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI12/MM4 N_XI22/XI12/NET33_XI22/XI12/MM4_d
+ N_XI22/XI12/NET34_XI22/XI12/MM4_g N_VDD_XI22/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI12/MM10 N_XI22/XI12/NET35_XI22/XI12/MM10_d
+ N_XI22/XI12/NET36_XI22/XI12/MM10_g N_VDD_XI22/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI12/MM11 N_XI22/XI12/NET36_XI22/XI12/MM11_d
+ N_XI22/XI12/NET35_XI22/XI12/MM11_g N_VDD_XI22/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI13/MM2 N_XI22/XI13/NET34_XI22/XI13/MM2_d
+ N_XI22/XI13/NET33_XI22/XI13/MM2_g N_VSS_XI22/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI13/MM3 N_XI22/XI13/NET33_XI22/XI13/MM3_d N_WL<40>_XI22/XI13/MM3_g
+ N_BLN<2>_XI22/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI13/MM0 N_XI22/XI13/NET34_XI22/XI13/MM0_d N_WL<40>_XI22/XI13/MM0_g
+ N_BL<2>_XI22/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI13/MM1 N_XI22/XI13/NET33_XI22/XI13/MM1_d
+ N_XI22/XI13/NET34_XI22/XI13/MM1_g N_VSS_XI22/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI13/MM9 N_XI22/XI13/NET36_XI22/XI13/MM9_d N_WL<41>_XI22/XI13/MM9_g
+ N_BL<2>_XI22/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI13/MM6 N_XI22/XI13/NET35_XI22/XI13/MM6_d
+ N_XI22/XI13/NET36_XI22/XI13/MM6_g N_VSS_XI22/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI13/MM7 N_XI22/XI13/NET36_XI22/XI13/MM7_d
+ N_XI22/XI13/NET35_XI22/XI13/MM7_g N_VSS_XI22/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI13/MM8 N_XI22/XI13/NET35_XI22/XI13/MM8_d N_WL<41>_XI22/XI13/MM8_g
+ N_BLN<2>_XI22/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI13/MM5 N_XI22/XI13/NET34_XI22/XI13/MM5_d
+ N_XI22/XI13/NET33_XI22/XI13/MM5_g N_VDD_XI22/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI13/MM4 N_XI22/XI13/NET33_XI22/XI13/MM4_d
+ N_XI22/XI13/NET34_XI22/XI13/MM4_g N_VDD_XI22/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI13/MM10 N_XI22/XI13/NET35_XI22/XI13/MM10_d
+ N_XI22/XI13/NET36_XI22/XI13/MM10_g N_VDD_XI22/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI13/MM11 N_XI22/XI13/NET36_XI22/XI13/MM11_d
+ N_XI22/XI13/NET35_XI22/XI13/MM11_g N_VDD_XI22/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI14/MM2 N_XI22/XI14/NET34_XI22/XI14/MM2_d
+ N_XI22/XI14/NET33_XI22/XI14/MM2_g N_VSS_XI22/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI14/MM3 N_XI22/XI14/NET33_XI22/XI14/MM3_d N_WL<40>_XI22/XI14/MM3_g
+ N_BLN<1>_XI22/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI14/MM0 N_XI22/XI14/NET34_XI22/XI14/MM0_d N_WL<40>_XI22/XI14/MM0_g
+ N_BL<1>_XI22/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI14/MM1 N_XI22/XI14/NET33_XI22/XI14/MM1_d
+ N_XI22/XI14/NET34_XI22/XI14/MM1_g N_VSS_XI22/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI14/MM9 N_XI22/XI14/NET36_XI22/XI14/MM9_d N_WL<41>_XI22/XI14/MM9_g
+ N_BL<1>_XI22/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI14/MM6 N_XI22/XI14/NET35_XI22/XI14/MM6_d
+ N_XI22/XI14/NET36_XI22/XI14/MM6_g N_VSS_XI22/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI14/MM7 N_XI22/XI14/NET36_XI22/XI14/MM7_d
+ N_XI22/XI14/NET35_XI22/XI14/MM7_g N_VSS_XI22/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI14/MM8 N_XI22/XI14/NET35_XI22/XI14/MM8_d N_WL<41>_XI22/XI14/MM8_g
+ N_BLN<1>_XI22/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI14/MM5 N_XI22/XI14/NET34_XI22/XI14/MM5_d
+ N_XI22/XI14/NET33_XI22/XI14/MM5_g N_VDD_XI22/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI14/MM4 N_XI22/XI14/NET33_XI22/XI14/MM4_d
+ N_XI22/XI14/NET34_XI22/XI14/MM4_g N_VDD_XI22/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI14/MM10 N_XI22/XI14/NET35_XI22/XI14/MM10_d
+ N_XI22/XI14/NET36_XI22/XI14/MM10_g N_VDD_XI22/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI14/MM11 N_XI22/XI14/NET36_XI22/XI14/MM11_d
+ N_XI22/XI14/NET35_XI22/XI14/MM11_g N_VDD_XI22/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI15/MM2 N_XI22/XI15/NET34_XI22/XI15/MM2_d
+ N_XI22/XI15/NET33_XI22/XI15/MM2_g N_VSS_XI22/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI15/MM3 N_XI22/XI15/NET33_XI22/XI15/MM3_d N_WL<40>_XI22/XI15/MM3_g
+ N_BLN<0>_XI22/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI15/MM0 N_XI22/XI15/NET34_XI22/XI15/MM0_d N_WL<40>_XI22/XI15/MM0_g
+ N_BL<0>_XI22/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI15/MM1 N_XI22/XI15/NET33_XI22/XI15/MM1_d
+ N_XI22/XI15/NET34_XI22/XI15/MM1_g N_VSS_XI22/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI15/MM9 N_XI22/XI15/NET36_XI22/XI15/MM9_d N_WL<41>_XI22/XI15/MM9_g
+ N_BL<0>_XI22/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI15/MM6 N_XI22/XI15/NET35_XI22/XI15/MM6_d
+ N_XI22/XI15/NET36_XI22/XI15/MM6_g N_VSS_XI22/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI15/MM7 N_XI22/XI15/NET36_XI22/XI15/MM7_d
+ N_XI22/XI15/NET35_XI22/XI15/MM7_g N_VSS_XI22/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI22/XI15/MM8 N_XI22/XI15/NET35_XI22/XI15/MM8_d N_WL<41>_XI22/XI15/MM8_g
+ N_BLN<0>_XI22/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI22/XI15/MM5 N_XI22/XI15/NET34_XI22/XI15/MM5_d
+ N_XI22/XI15/NET33_XI22/XI15/MM5_g N_VDD_XI22/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI15/MM4 N_XI22/XI15/NET33_XI22/XI15/MM4_d
+ N_XI22/XI15/NET34_XI22/XI15/MM4_g N_VDD_XI22/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI15/MM10 N_XI22/XI15/NET35_XI22/XI15/MM10_d
+ N_XI22/XI15/NET36_XI22/XI15/MM10_g N_VDD_XI22/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI22/XI15/MM11 N_XI22/XI15/NET36_XI22/XI15/MM11_d
+ N_XI22/XI15/NET35_XI22/XI15/MM11_g N_VDD_XI22/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI0/MM2 N_XI23/XI0/NET34_XI23/XI0/MM2_d N_XI23/XI0/NET33_XI23/XI0/MM2_g
+ N_VSS_XI23/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI0/MM3 N_XI23/XI0/NET33_XI23/XI0/MM3_d N_WL<42>_XI23/XI0/MM3_g
+ N_BLN<15>_XI23/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI0/MM0 N_XI23/XI0/NET34_XI23/XI0/MM0_d N_WL<42>_XI23/XI0/MM0_g
+ N_BL<15>_XI23/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI0/MM1 N_XI23/XI0/NET33_XI23/XI0/MM1_d N_XI23/XI0/NET34_XI23/XI0/MM1_g
+ N_VSS_XI23/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI0/MM9 N_XI23/XI0/NET36_XI23/XI0/MM9_d N_WL<43>_XI23/XI0/MM9_g
+ N_BL<15>_XI23/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI0/MM6 N_XI23/XI0/NET35_XI23/XI0/MM6_d N_XI23/XI0/NET36_XI23/XI0/MM6_g
+ N_VSS_XI23/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI0/MM7 N_XI23/XI0/NET36_XI23/XI0/MM7_d N_XI23/XI0/NET35_XI23/XI0/MM7_g
+ N_VSS_XI23/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI0/MM8 N_XI23/XI0/NET35_XI23/XI0/MM8_d N_WL<43>_XI23/XI0/MM8_g
+ N_BLN<15>_XI23/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI0/MM5 N_XI23/XI0/NET34_XI23/XI0/MM5_d N_XI23/XI0/NET33_XI23/XI0/MM5_g
+ N_VDD_XI23/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI0/MM4 N_XI23/XI0/NET33_XI23/XI0/MM4_d N_XI23/XI0/NET34_XI23/XI0/MM4_g
+ N_VDD_XI23/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI0/MM10 N_XI23/XI0/NET35_XI23/XI0/MM10_d N_XI23/XI0/NET36_XI23/XI0/MM10_g
+ N_VDD_XI23/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI0/MM11 N_XI23/XI0/NET36_XI23/XI0/MM11_d N_XI23/XI0/NET35_XI23/XI0/MM11_g
+ N_VDD_XI23/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI1/MM2 N_XI23/XI1/NET34_XI23/XI1/MM2_d N_XI23/XI1/NET33_XI23/XI1/MM2_g
+ N_VSS_XI23/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI1/MM3 N_XI23/XI1/NET33_XI23/XI1/MM3_d N_WL<42>_XI23/XI1/MM3_g
+ N_BLN<14>_XI23/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI1/MM0 N_XI23/XI1/NET34_XI23/XI1/MM0_d N_WL<42>_XI23/XI1/MM0_g
+ N_BL<14>_XI23/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI1/MM1 N_XI23/XI1/NET33_XI23/XI1/MM1_d N_XI23/XI1/NET34_XI23/XI1/MM1_g
+ N_VSS_XI23/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI1/MM9 N_XI23/XI1/NET36_XI23/XI1/MM9_d N_WL<43>_XI23/XI1/MM9_g
+ N_BL<14>_XI23/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI1/MM6 N_XI23/XI1/NET35_XI23/XI1/MM6_d N_XI23/XI1/NET36_XI23/XI1/MM6_g
+ N_VSS_XI23/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI1/MM7 N_XI23/XI1/NET36_XI23/XI1/MM7_d N_XI23/XI1/NET35_XI23/XI1/MM7_g
+ N_VSS_XI23/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI1/MM8 N_XI23/XI1/NET35_XI23/XI1/MM8_d N_WL<43>_XI23/XI1/MM8_g
+ N_BLN<14>_XI23/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI1/MM5 N_XI23/XI1/NET34_XI23/XI1/MM5_d N_XI23/XI1/NET33_XI23/XI1/MM5_g
+ N_VDD_XI23/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI1/MM4 N_XI23/XI1/NET33_XI23/XI1/MM4_d N_XI23/XI1/NET34_XI23/XI1/MM4_g
+ N_VDD_XI23/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI1/MM10 N_XI23/XI1/NET35_XI23/XI1/MM10_d N_XI23/XI1/NET36_XI23/XI1/MM10_g
+ N_VDD_XI23/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI1/MM11 N_XI23/XI1/NET36_XI23/XI1/MM11_d N_XI23/XI1/NET35_XI23/XI1/MM11_g
+ N_VDD_XI23/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI2/MM2 N_XI23/XI2/NET34_XI23/XI2/MM2_d N_XI23/XI2/NET33_XI23/XI2/MM2_g
+ N_VSS_XI23/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI2/MM3 N_XI23/XI2/NET33_XI23/XI2/MM3_d N_WL<42>_XI23/XI2/MM3_g
+ N_BLN<13>_XI23/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI2/MM0 N_XI23/XI2/NET34_XI23/XI2/MM0_d N_WL<42>_XI23/XI2/MM0_g
+ N_BL<13>_XI23/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI2/MM1 N_XI23/XI2/NET33_XI23/XI2/MM1_d N_XI23/XI2/NET34_XI23/XI2/MM1_g
+ N_VSS_XI23/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI2/MM9 N_XI23/XI2/NET36_XI23/XI2/MM9_d N_WL<43>_XI23/XI2/MM9_g
+ N_BL<13>_XI23/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI2/MM6 N_XI23/XI2/NET35_XI23/XI2/MM6_d N_XI23/XI2/NET36_XI23/XI2/MM6_g
+ N_VSS_XI23/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI2/MM7 N_XI23/XI2/NET36_XI23/XI2/MM7_d N_XI23/XI2/NET35_XI23/XI2/MM7_g
+ N_VSS_XI23/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI2/MM8 N_XI23/XI2/NET35_XI23/XI2/MM8_d N_WL<43>_XI23/XI2/MM8_g
+ N_BLN<13>_XI23/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI2/MM5 N_XI23/XI2/NET34_XI23/XI2/MM5_d N_XI23/XI2/NET33_XI23/XI2/MM5_g
+ N_VDD_XI23/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI2/MM4 N_XI23/XI2/NET33_XI23/XI2/MM4_d N_XI23/XI2/NET34_XI23/XI2/MM4_g
+ N_VDD_XI23/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI2/MM10 N_XI23/XI2/NET35_XI23/XI2/MM10_d N_XI23/XI2/NET36_XI23/XI2/MM10_g
+ N_VDD_XI23/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI2/MM11 N_XI23/XI2/NET36_XI23/XI2/MM11_d N_XI23/XI2/NET35_XI23/XI2/MM11_g
+ N_VDD_XI23/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI3/MM2 N_XI23/XI3/NET34_XI23/XI3/MM2_d N_XI23/XI3/NET33_XI23/XI3/MM2_g
+ N_VSS_XI23/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI3/MM3 N_XI23/XI3/NET33_XI23/XI3/MM3_d N_WL<42>_XI23/XI3/MM3_g
+ N_BLN<12>_XI23/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI3/MM0 N_XI23/XI3/NET34_XI23/XI3/MM0_d N_WL<42>_XI23/XI3/MM0_g
+ N_BL<12>_XI23/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI3/MM1 N_XI23/XI3/NET33_XI23/XI3/MM1_d N_XI23/XI3/NET34_XI23/XI3/MM1_g
+ N_VSS_XI23/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI3/MM9 N_XI23/XI3/NET36_XI23/XI3/MM9_d N_WL<43>_XI23/XI3/MM9_g
+ N_BL<12>_XI23/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI3/MM6 N_XI23/XI3/NET35_XI23/XI3/MM6_d N_XI23/XI3/NET36_XI23/XI3/MM6_g
+ N_VSS_XI23/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI3/MM7 N_XI23/XI3/NET36_XI23/XI3/MM7_d N_XI23/XI3/NET35_XI23/XI3/MM7_g
+ N_VSS_XI23/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI3/MM8 N_XI23/XI3/NET35_XI23/XI3/MM8_d N_WL<43>_XI23/XI3/MM8_g
+ N_BLN<12>_XI23/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI3/MM5 N_XI23/XI3/NET34_XI23/XI3/MM5_d N_XI23/XI3/NET33_XI23/XI3/MM5_g
+ N_VDD_XI23/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI3/MM4 N_XI23/XI3/NET33_XI23/XI3/MM4_d N_XI23/XI3/NET34_XI23/XI3/MM4_g
+ N_VDD_XI23/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI3/MM10 N_XI23/XI3/NET35_XI23/XI3/MM10_d N_XI23/XI3/NET36_XI23/XI3/MM10_g
+ N_VDD_XI23/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI3/MM11 N_XI23/XI3/NET36_XI23/XI3/MM11_d N_XI23/XI3/NET35_XI23/XI3/MM11_g
+ N_VDD_XI23/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI4/MM2 N_XI23/XI4/NET34_XI23/XI4/MM2_d N_XI23/XI4/NET33_XI23/XI4/MM2_g
+ N_VSS_XI23/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI4/MM3 N_XI23/XI4/NET33_XI23/XI4/MM3_d N_WL<42>_XI23/XI4/MM3_g
+ N_BLN<11>_XI23/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI4/MM0 N_XI23/XI4/NET34_XI23/XI4/MM0_d N_WL<42>_XI23/XI4/MM0_g
+ N_BL<11>_XI23/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI4/MM1 N_XI23/XI4/NET33_XI23/XI4/MM1_d N_XI23/XI4/NET34_XI23/XI4/MM1_g
+ N_VSS_XI23/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI4/MM9 N_XI23/XI4/NET36_XI23/XI4/MM9_d N_WL<43>_XI23/XI4/MM9_g
+ N_BL<11>_XI23/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI4/MM6 N_XI23/XI4/NET35_XI23/XI4/MM6_d N_XI23/XI4/NET36_XI23/XI4/MM6_g
+ N_VSS_XI23/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI4/MM7 N_XI23/XI4/NET36_XI23/XI4/MM7_d N_XI23/XI4/NET35_XI23/XI4/MM7_g
+ N_VSS_XI23/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI4/MM8 N_XI23/XI4/NET35_XI23/XI4/MM8_d N_WL<43>_XI23/XI4/MM8_g
+ N_BLN<11>_XI23/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI4/MM5 N_XI23/XI4/NET34_XI23/XI4/MM5_d N_XI23/XI4/NET33_XI23/XI4/MM5_g
+ N_VDD_XI23/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI4/MM4 N_XI23/XI4/NET33_XI23/XI4/MM4_d N_XI23/XI4/NET34_XI23/XI4/MM4_g
+ N_VDD_XI23/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI4/MM10 N_XI23/XI4/NET35_XI23/XI4/MM10_d N_XI23/XI4/NET36_XI23/XI4/MM10_g
+ N_VDD_XI23/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI4/MM11 N_XI23/XI4/NET36_XI23/XI4/MM11_d N_XI23/XI4/NET35_XI23/XI4/MM11_g
+ N_VDD_XI23/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI5/MM2 N_XI23/XI5/NET34_XI23/XI5/MM2_d N_XI23/XI5/NET33_XI23/XI5/MM2_g
+ N_VSS_XI23/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI5/MM3 N_XI23/XI5/NET33_XI23/XI5/MM3_d N_WL<42>_XI23/XI5/MM3_g
+ N_BLN<10>_XI23/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI5/MM0 N_XI23/XI5/NET34_XI23/XI5/MM0_d N_WL<42>_XI23/XI5/MM0_g
+ N_BL<10>_XI23/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI5/MM1 N_XI23/XI5/NET33_XI23/XI5/MM1_d N_XI23/XI5/NET34_XI23/XI5/MM1_g
+ N_VSS_XI23/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI5/MM9 N_XI23/XI5/NET36_XI23/XI5/MM9_d N_WL<43>_XI23/XI5/MM9_g
+ N_BL<10>_XI23/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI5/MM6 N_XI23/XI5/NET35_XI23/XI5/MM6_d N_XI23/XI5/NET36_XI23/XI5/MM6_g
+ N_VSS_XI23/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI5/MM7 N_XI23/XI5/NET36_XI23/XI5/MM7_d N_XI23/XI5/NET35_XI23/XI5/MM7_g
+ N_VSS_XI23/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI5/MM8 N_XI23/XI5/NET35_XI23/XI5/MM8_d N_WL<43>_XI23/XI5/MM8_g
+ N_BLN<10>_XI23/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI5/MM5 N_XI23/XI5/NET34_XI23/XI5/MM5_d N_XI23/XI5/NET33_XI23/XI5/MM5_g
+ N_VDD_XI23/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI5/MM4 N_XI23/XI5/NET33_XI23/XI5/MM4_d N_XI23/XI5/NET34_XI23/XI5/MM4_g
+ N_VDD_XI23/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI5/MM10 N_XI23/XI5/NET35_XI23/XI5/MM10_d N_XI23/XI5/NET36_XI23/XI5/MM10_g
+ N_VDD_XI23/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI5/MM11 N_XI23/XI5/NET36_XI23/XI5/MM11_d N_XI23/XI5/NET35_XI23/XI5/MM11_g
+ N_VDD_XI23/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI6/MM2 N_XI23/XI6/NET34_XI23/XI6/MM2_d N_XI23/XI6/NET33_XI23/XI6/MM2_g
+ N_VSS_XI23/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM3 N_XI23/XI6/NET33_XI23/XI6/MM3_d N_WL<42>_XI23/XI6/MM3_g
+ N_BLN<9>_XI23/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM0 N_XI23/XI6/NET34_XI23/XI6/MM0_d N_WL<42>_XI23/XI6/MM0_g
+ N_BL<9>_XI23/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM1 N_XI23/XI6/NET33_XI23/XI6/MM1_d N_XI23/XI6/NET34_XI23/XI6/MM1_g
+ N_VSS_XI23/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM9 N_XI23/XI6/NET36_XI23/XI6/MM9_d N_WL<43>_XI23/XI6/MM9_g
+ N_BL<9>_XI23/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM6 N_XI23/XI6/NET35_XI23/XI6/MM6_d N_XI23/XI6/NET36_XI23/XI6/MM6_g
+ N_VSS_XI23/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM7 N_XI23/XI6/NET36_XI23/XI6/MM7_d N_XI23/XI6/NET35_XI23/XI6/MM7_g
+ N_VSS_XI23/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM8 N_XI23/XI6/NET35_XI23/XI6/MM8_d N_WL<43>_XI23/XI6/MM8_g
+ N_BLN<9>_XI23/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI6/MM5 N_XI23/XI6/NET34_XI23/XI6/MM5_d N_XI23/XI6/NET33_XI23/XI6/MM5_g
+ N_VDD_XI23/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI6/MM4 N_XI23/XI6/NET33_XI23/XI6/MM4_d N_XI23/XI6/NET34_XI23/XI6/MM4_g
+ N_VDD_XI23/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI6/MM10 N_XI23/XI6/NET35_XI23/XI6/MM10_d N_XI23/XI6/NET36_XI23/XI6/MM10_g
+ N_VDD_XI23/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI6/MM11 N_XI23/XI6/NET36_XI23/XI6/MM11_d N_XI23/XI6/NET35_XI23/XI6/MM11_g
+ N_VDD_XI23/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI7/MM2 N_XI23/XI7/NET34_XI23/XI7/MM2_d N_XI23/XI7/NET33_XI23/XI7/MM2_g
+ N_VSS_XI23/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM3 N_XI23/XI7/NET33_XI23/XI7/MM3_d N_WL<42>_XI23/XI7/MM3_g
+ N_BLN<8>_XI23/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM0 N_XI23/XI7/NET34_XI23/XI7/MM0_d N_WL<42>_XI23/XI7/MM0_g
+ N_BL<8>_XI23/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM1 N_XI23/XI7/NET33_XI23/XI7/MM1_d N_XI23/XI7/NET34_XI23/XI7/MM1_g
+ N_VSS_XI23/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM9 N_XI23/XI7/NET36_XI23/XI7/MM9_d N_WL<43>_XI23/XI7/MM9_g
+ N_BL<8>_XI23/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM6 N_XI23/XI7/NET35_XI23/XI7/MM6_d N_XI23/XI7/NET36_XI23/XI7/MM6_g
+ N_VSS_XI23/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM7 N_XI23/XI7/NET36_XI23/XI7/MM7_d N_XI23/XI7/NET35_XI23/XI7/MM7_g
+ N_VSS_XI23/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM8 N_XI23/XI7/NET35_XI23/XI7/MM8_d N_WL<43>_XI23/XI7/MM8_g
+ N_BLN<8>_XI23/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI7/MM5 N_XI23/XI7/NET34_XI23/XI7/MM5_d N_XI23/XI7/NET33_XI23/XI7/MM5_g
+ N_VDD_XI23/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI7/MM4 N_XI23/XI7/NET33_XI23/XI7/MM4_d N_XI23/XI7/NET34_XI23/XI7/MM4_g
+ N_VDD_XI23/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI7/MM10 N_XI23/XI7/NET35_XI23/XI7/MM10_d N_XI23/XI7/NET36_XI23/XI7/MM10_g
+ N_VDD_XI23/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI7/MM11 N_XI23/XI7/NET36_XI23/XI7/MM11_d N_XI23/XI7/NET35_XI23/XI7/MM11_g
+ N_VDD_XI23/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI8/MM2 N_XI23/XI8/NET34_XI23/XI8/MM2_d N_XI23/XI8/NET33_XI23/XI8/MM2_g
+ N_VSS_XI23/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM3 N_XI23/XI8/NET33_XI23/XI8/MM3_d N_WL<42>_XI23/XI8/MM3_g
+ N_BLN<7>_XI23/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM0 N_XI23/XI8/NET34_XI23/XI8/MM0_d N_WL<42>_XI23/XI8/MM0_g
+ N_BL<7>_XI23/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM1 N_XI23/XI8/NET33_XI23/XI8/MM1_d N_XI23/XI8/NET34_XI23/XI8/MM1_g
+ N_VSS_XI23/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM9 N_XI23/XI8/NET36_XI23/XI8/MM9_d N_WL<43>_XI23/XI8/MM9_g
+ N_BL<7>_XI23/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM6 N_XI23/XI8/NET35_XI23/XI8/MM6_d N_XI23/XI8/NET36_XI23/XI8/MM6_g
+ N_VSS_XI23/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM7 N_XI23/XI8/NET36_XI23/XI8/MM7_d N_XI23/XI8/NET35_XI23/XI8/MM7_g
+ N_VSS_XI23/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM8 N_XI23/XI8/NET35_XI23/XI8/MM8_d N_WL<43>_XI23/XI8/MM8_g
+ N_BLN<7>_XI23/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI8/MM5 N_XI23/XI8/NET34_XI23/XI8/MM5_d N_XI23/XI8/NET33_XI23/XI8/MM5_g
+ N_VDD_XI23/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI8/MM4 N_XI23/XI8/NET33_XI23/XI8/MM4_d N_XI23/XI8/NET34_XI23/XI8/MM4_g
+ N_VDD_XI23/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI8/MM10 N_XI23/XI8/NET35_XI23/XI8/MM10_d N_XI23/XI8/NET36_XI23/XI8/MM10_g
+ N_VDD_XI23/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI8/MM11 N_XI23/XI8/NET36_XI23/XI8/MM11_d N_XI23/XI8/NET35_XI23/XI8/MM11_g
+ N_VDD_XI23/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI9/MM2 N_XI23/XI9/NET34_XI23/XI9/MM2_d N_XI23/XI9/NET33_XI23/XI9/MM2_g
+ N_VSS_XI23/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM3 N_XI23/XI9/NET33_XI23/XI9/MM3_d N_WL<42>_XI23/XI9/MM3_g
+ N_BLN<6>_XI23/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM0 N_XI23/XI9/NET34_XI23/XI9/MM0_d N_WL<42>_XI23/XI9/MM0_g
+ N_BL<6>_XI23/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM1 N_XI23/XI9/NET33_XI23/XI9/MM1_d N_XI23/XI9/NET34_XI23/XI9/MM1_g
+ N_VSS_XI23/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM9 N_XI23/XI9/NET36_XI23/XI9/MM9_d N_WL<43>_XI23/XI9/MM9_g
+ N_BL<6>_XI23/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM6 N_XI23/XI9/NET35_XI23/XI9/MM6_d N_XI23/XI9/NET36_XI23/XI9/MM6_g
+ N_VSS_XI23/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM7 N_XI23/XI9/NET36_XI23/XI9/MM7_d N_XI23/XI9/NET35_XI23/XI9/MM7_g
+ N_VSS_XI23/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM8 N_XI23/XI9/NET35_XI23/XI9/MM8_d N_WL<43>_XI23/XI9/MM8_g
+ N_BLN<6>_XI23/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI9/MM5 N_XI23/XI9/NET34_XI23/XI9/MM5_d N_XI23/XI9/NET33_XI23/XI9/MM5_g
+ N_VDD_XI23/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI9/MM4 N_XI23/XI9/NET33_XI23/XI9/MM4_d N_XI23/XI9/NET34_XI23/XI9/MM4_g
+ N_VDD_XI23/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI9/MM10 N_XI23/XI9/NET35_XI23/XI9/MM10_d N_XI23/XI9/NET36_XI23/XI9/MM10_g
+ N_VDD_XI23/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI9/MM11 N_XI23/XI9/NET36_XI23/XI9/MM11_d N_XI23/XI9/NET35_XI23/XI9/MM11_g
+ N_VDD_XI23/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI10/MM2 N_XI23/XI10/NET34_XI23/XI10/MM2_d
+ N_XI23/XI10/NET33_XI23/XI10/MM2_g N_VSS_XI23/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI10/MM3 N_XI23/XI10/NET33_XI23/XI10/MM3_d N_WL<42>_XI23/XI10/MM3_g
+ N_BLN<5>_XI23/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI10/MM0 N_XI23/XI10/NET34_XI23/XI10/MM0_d N_WL<42>_XI23/XI10/MM0_g
+ N_BL<5>_XI23/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI10/MM1 N_XI23/XI10/NET33_XI23/XI10/MM1_d
+ N_XI23/XI10/NET34_XI23/XI10/MM1_g N_VSS_XI23/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI10/MM9 N_XI23/XI10/NET36_XI23/XI10/MM9_d N_WL<43>_XI23/XI10/MM9_g
+ N_BL<5>_XI23/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI10/MM6 N_XI23/XI10/NET35_XI23/XI10/MM6_d
+ N_XI23/XI10/NET36_XI23/XI10/MM6_g N_VSS_XI23/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI10/MM7 N_XI23/XI10/NET36_XI23/XI10/MM7_d
+ N_XI23/XI10/NET35_XI23/XI10/MM7_g N_VSS_XI23/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI10/MM8 N_XI23/XI10/NET35_XI23/XI10/MM8_d N_WL<43>_XI23/XI10/MM8_g
+ N_BLN<5>_XI23/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI10/MM5 N_XI23/XI10/NET34_XI23/XI10/MM5_d
+ N_XI23/XI10/NET33_XI23/XI10/MM5_g N_VDD_XI23/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI10/MM4 N_XI23/XI10/NET33_XI23/XI10/MM4_d
+ N_XI23/XI10/NET34_XI23/XI10/MM4_g N_VDD_XI23/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI10/MM10 N_XI23/XI10/NET35_XI23/XI10/MM10_d
+ N_XI23/XI10/NET36_XI23/XI10/MM10_g N_VDD_XI23/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI10/MM11 N_XI23/XI10/NET36_XI23/XI10/MM11_d
+ N_XI23/XI10/NET35_XI23/XI10/MM11_g N_VDD_XI23/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI11/MM2 N_XI23/XI11/NET34_XI23/XI11/MM2_d
+ N_XI23/XI11/NET33_XI23/XI11/MM2_g N_VSS_XI23/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI11/MM3 N_XI23/XI11/NET33_XI23/XI11/MM3_d N_WL<42>_XI23/XI11/MM3_g
+ N_BLN<4>_XI23/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI11/MM0 N_XI23/XI11/NET34_XI23/XI11/MM0_d N_WL<42>_XI23/XI11/MM0_g
+ N_BL<4>_XI23/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI11/MM1 N_XI23/XI11/NET33_XI23/XI11/MM1_d
+ N_XI23/XI11/NET34_XI23/XI11/MM1_g N_VSS_XI23/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI11/MM9 N_XI23/XI11/NET36_XI23/XI11/MM9_d N_WL<43>_XI23/XI11/MM9_g
+ N_BL<4>_XI23/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI11/MM6 N_XI23/XI11/NET35_XI23/XI11/MM6_d
+ N_XI23/XI11/NET36_XI23/XI11/MM6_g N_VSS_XI23/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI11/MM7 N_XI23/XI11/NET36_XI23/XI11/MM7_d
+ N_XI23/XI11/NET35_XI23/XI11/MM7_g N_VSS_XI23/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI11/MM8 N_XI23/XI11/NET35_XI23/XI11/MM8_d N_WL<43>_XI23/XI11/MM8_g
+ N_BLN<4>_XI23/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI11/MM5 N_XI23/XI11/NET34_XI23/XI11/MM5_d
+ N_XI23/XI11/NET33_XI23/XI11/MM5_g N_VDD_XI23/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI11/MM4 N_XI23/XI11/NET33_XI23/XI11/MM4_d
+ N_XI23/XI11/NET34_XI23/XI11/MM4_g N_VDD_XI23/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI11/MM10 N_XI23/XI11/NET35_XI23/XI11/MM10_d
+ N_XI23/XI11/NET36_XI23/XI11/MM10_g N_VDD_XI23/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI11/MM11 N_XI23/XI11/NET36_XI23/XI11/MM11_d
+ N_XI23/XI11/NET35_XI23/XI11/MM11_g N_VDD_XI23/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI12/MM2 N_XI23/XI12/NET34_XI23/XI12/MM2_d
+ N_XI23/XI12/NET33_XI23/XI12/MM2_g N_VSS_XI23/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI12/MM3 N_XI23/XI12/NET33_XI23/XI12/MM3_d N_WL<42>_XI23/XI12/MM3_g
+ N_BLN<3>_XI23/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI12/MM0 N_XI23/XI12/NET34_XI23/XI12/MM0_d N_WL<42>_XI23/XI12/MM0_g
+ N_BL<3>_XI23/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI12/MM1 N_XI23/XI12/NET33_XI23/XI12/MM1_d
+ N_XI23/XI12/NET34_XI23/XI12/MM1_g N_VSS_XI23/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI12/MM9 N_XI23/XI12/NET36_XI23/XI12/MM9_d N_WL<43>_XI23/XI12/MM9_g
+ N_BL<3>_XI23/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI12/MM6 N_XI23/XI12/NET35_XI23/XI12/MM6_d
+ N_XI23/XI12/NET36_XI23/XI12/MM6_g N_VSS_XI23/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI12/MM7 N_XI23/XI12/NET36_XI23/XI12/MM7_d
+ N_XI23/XI12/NET35_XI23/XI12/MM7_g N_VSS_XI23/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI12/MM8 N_XI23/XI12/NET35_XI23/XI12/MM8_d N_WL<43>_XI23/XI12/MM8_g
+ N_BLN<3>_XI23/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI12/MM5 N_XI23/XI12/NET34_XI23/XI12/MM5_d
+ N_XI23/XI12/NET33_XI23/XI12/MM5_g N_VDD_XI23/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI12/MM4 N_XI23/XI12/NET33_XI23/XI12/MM4_d
+ N_XI23/XI12/NET34_XI23/XI12/MM4_g N_VDD_XI23/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI12/MM10 N_XI23/XI12/NET35_XI23/XI12/MM10_d
+ N_XI23/XI12/NET36_XI23/XI12/MM10_g N_VDD_XI23/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI12/MM11 N_XI23/XI12/NET36_XI23/XI12/MM11_d
+ N_XI23/XI12/NET35_XI23/XI12/MM11_g N_VDD_XI23/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI13/MM2 N_XI23/XI13/NET34_XI23/XI13/MM2_d
+ N_XI23/XI13/NET33_XI23/XI13/MM2_g N_VSS_XI23/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI13/MM3 N_XI23/XI13/NET33_XI23/XI13/MM3_d N_WL<42>_XI23/XI13/MM3_g
+ N_BLN<2>_XI23/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI13/MM0 N_XI23/XI13/NET34_XI23/XI13/MM0_d N_WL<42>_XI23/XI13/MM0_g
+ N_BL<2>_XI23/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI13/MM1 N_XI23/XI13/NET33_XI23/XI13/MM1_d
+ N_XI23/XI13/NET34_XI23/XI13/MM1_g N_VSS_XI23/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI13/MM9 N_XI23/XI13/NET36_XI23/XI13/MM9_d N_WL<43>_XI23/XI13/MM9_g
+ N_BL<2>_XI23/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI13/MM6 N_XI23/XI13/NET35_XI23/XI13/MM6_d
+ N_XI23/XI13/NET36_XI23/XI13/MM6_g N_VSS_XI23/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI13/MM7 N_XI23/XI13/NET36_XI23/XI13/MM7_d
+ N_XI23/XI13/NET35_XI23/XI13/MM7_g N_VSS_XI23/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI13/MM8 N_XI23/XI13/NET35_XI23/XI13/MM8_d N_WL<43>_XI23/XI13/MM8_g
+ N_BLN<2>_XI23/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI13/MM5 N_XI23/XI13/NET34_XI23/XI13/MM5_d
+ N_XI23/XI13/NET33_XI23/XI13/MM5_g N_VDD_XI23/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI13/MM4 N_XI23/XI13/NET33_XI23/XI13/MM4_d
+ N_XI23/XI13/NET34_XI23/XI13/MM4_g N_VDD_XI23/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI13/MM10 N_XI23/XI13/NET35_XI23/XI13/MM10_d
+ N_XI23/XI13/NET36_XI23/XI13/MM10_g N_VDD_XI23/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI13/MM11 N_XI23/XI13/NET36_XI23/XI13/MM11_d
+ N_XI23/XI13/NET35_XI23/XI13/MM11_g N_VDD_XI23/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI14/MM2 N_XI23/XI14/NET34_XI23/XI14/MM2_d
+ N_XI23/XI14/NET33_XI23/XI14/MM2_g N_VSS_XI23/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI14/MM3 N_XI23/XI14/NET33_XI23/XI14/MM3_d N_WL<42>_XI23/XI14/MM3_g
+ N_BLN<1>_XI23/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI14/MM0 N_XI23/XI14/NET34_XI23/XI14/MM0_d N_WL<42>_XI23/XI14/MM0_g
+ N_BL<1>_XI23/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI14/MM1 N_XI23/XI14/NET33_XI23/XI14/MM1_d
+ N_XI23/XI14/NET34_XI23/XI14/MM1_g N_VSS_XI23/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI14/MM9 N_XI23/XI14/NET36_XI23/XI14/MM9_d N_WL<43>_XI23/XI14/MM9_g
+ N_BL<1>_XI23/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI14/MM6 N_XI23/XI14/NET35_XI23/XI14/MM6_d
+ N_XI23/XI14/NET36_XI23/XI14/MM6_g N_VSS_XI23/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI14/MM7 N_XI23/XI14/NET36_XI23/XI14/MM7_d
+ N_XI23/XI14/NET35_XI23/XI14/MM7_g N_VSS_XI23/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI14/MM8 N_XI23/XI14/NET35_XI23/XI14/MM8_d N_WL<43>_XI23/XI14/MM8_g
+ N_BLN<1>_XI23/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI14/MM5 N_XI23/XI14/NET34_XI23/XI14/MM5_d
+ N_XI23/XI14/NET33_XI23/XI14/MM5_g N_VDD_XI23/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI14/MM4 N_XI23/XI14/NET33_XI23/XI14/MM4_d
+ N_XI23/XI14/NET34_XI23/XI14/MM4_g N_VDD_XI23/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI14/MM10 N_XI23/XI14/NET35_XI23/XI14/MM10_d
+ N_XI23/XI14/NET36_XI23/XI14/MM10_g N_VDD_XI23/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI14/MM11 N_XI23/XI14/NET36_XI23/XI14/MM11_d
+ N_XI23/XI14/NET35_XI23/XI14/MM11_g N_VDD_XI23/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI15/MM2 N_XI23/XI15/NET34_XI23/XI15/MM2_d
+ N_XI23/XI15/NET33_XI23/XI15/MM2_g N_VSS_XI23/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI15/MM3 N_XI23/XI15/NET33_XI23/XI15/MM3_d N_WL<42>_XI23/XI15/MM3_g
+ N_BLN<0>_XI23/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI15/MM0 N_XI23/XI15/NET34_XI23/XI15/MM0_d N_WL<42>_XI23/XI15/MM0_g
+ N_BL<0>_XI23/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI15/MM1 N_XI23/XI15/NET33_XI23/XI15/MM1_d
+ N_XI23/XI15/NET34_XI23/XI15/MM1_g N_VSS_XI23/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI15/MM9 N_XI23/XI15/NET36_XI23/XI15/MM9_d N_WL<43>_XI23/XI15/MM9_g
+ N_BL<0>_XI23/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI15/MM6 N_XI23/XI15/NET35_XI23/XI15/MM6_d
+ N_XI23/XI15/NET36_XI23/XI15/MM6_g N_VSS_XI23/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI15/MM7 N_XI23/XI15/NET36_XI23/XI15/MM7_d
+ N_XI23/XI15/NET35_XI23/XI15/MM7_g N_VSS_XI23/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI23/XI15/MM8 N_XI23/XI15/NET35_XI23/XI15/MM8_d N_WL<43>_XI23/XI15/MM8_g
+ N_BLN<0>_XI23/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI23/XI15/MM5 N_XI23/XI15/NET34_XI23/XI15/MM5_d
+ N_XI23/XI15/NET33_XI23/XI15/MM5_g N_VDD_XI23/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI15/MM4 N_XI23/XI15/NET33_XI23/XI15/MM4_d
+ N_XI23/XI15/NET34_XI23/XI15/MM4_g N_VDD_XI23/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI15/MM10 N_XI23/XI15/NET35_XI23/XI15/MM10_d
+ N_XI23/XI15/NET36_XI23/XI15/MM10_g N_VDD_XI23/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI23/XI15/MM11 N_XI23/XI15/NET36_XI23/XI15/MM11_d
+ N_XI23/XI15/NET35_XI23/XI15/MM11_g N_VDD_XI23/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI0/MM2 N_XI24/XI0/NET34_XI24/XI0/MM2_d N_XI24/XI0/NET33_XI24/XI0/MM2_g
+ N_VSS_XI24/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI0/MM3 N_XI24/XI0/NET33_XI24/XI0/MM3_d N_WL<44>_XI24/XI0/MM3_g
+ N_BLN<15>_XI24/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI0/MM0 N_XI24/XI0/NET34_XI24/XI0/MM0_d N_WL<44>_XI24/XI0/MM0_g
+ N_BL<15>_XI24/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI0/MM1 N_XI24/XI0/NET33_XI24/XI0/MM1_d N_XI24/XI0/NET34_XI24/XI0/MM1_g
+ N_VSS_XI24/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI0/MM9 N_XI24/XI0/NET36_XI24/XI0/MM9_d N_WL<45>_XI24/XI0/MM9_g
+ N_BL<15>_XI24/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI0/MM6 N_XI24/XI0/NET35_XI24/XI0/MM6_d N_XI24/XI0/NET36_XI24/XI0/MM6_g
+ N_VSS_XI24/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI0/MM7 N_XI24/XI0/NET36_XI24/XI0/MM7_d N_XI24/XI0/NET35_XI24/XI0/MM7_g
+ N_VSS_XI24/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI0/MM8 N_XI24/XI0/NET35_XI24/XI0/MM8_d N_WL<45>_XI24/XI0/MM8_g
+ N_BLN<15>_XI24/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI0/MM5 N_XI24/XI0/NET34_XI24/XI0/MM5_d N_XI24/XI0/NET33_XI24/XI0/MM5_g
+ N_VDD_XI24/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI0/MM4 N_XI24/XI0/NET33_XI24/XI0/MM4_d N_XI24/XI0/NET34_XI24/XI0/MM4_g
+ N_VDD_XI24/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI0/MM10 N_XI24/XI0/NET35_XI24/XI0/MM10_d N_XI24/XI0/NET36_XI24/XI0/MM10_g
+ N_VDD_XI24/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI0/MM11 N_XI24/XI0/NET36_XI24/XI0/MM11_d N_XI24/XI0/NET35_XI24/XI0/MM11_g
+ N_VDD_XI24/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI1/MM2 N_XI24/XI1/NET34_XI24/XI1/MM2_d N_XI24/XI1/NET33_XI24/XI1/MM2_g
+ N_VSS_XI24/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI1/MM3 N_XI24/XI1/NET33_XI24/XI1/MM3_d N_WL<44>_XI24/XI1/MM3_g
+ N_BLN<14>_XI24/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI1/MM0 N_XI24/XI1/NET34_XI24/XI1/MM0_d N_WL<44>_XI24/XI1/MM0_g
+ N_BL<14>_XI24/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI1/MM1 N_XI24/XI1/NET33_XI24/XI1/MM1_d N_XI24/XI1/NET34_XI24/XI1/MM1_g
+ N_VSS_XI24/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI1/MM9 N_XI24/XI1/NET36_XI24/XI1/MM9_d N_WL<45>_XI24/XI1/MM9_g
+ N_BL<14>_XI24/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI1/MM6 N_XI24/XI1/NET35_XI24/XI1/MM6_d N_XI24/XI1/NET36_XI24/XI1/MM6_g
+ N_VSS_XI24/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI1/MM7 N_XI24/XI1/NET36_XI24/XI1/MM7_d N_XI24/XI1/NET35_XI24/XI1/MM7_g
+ N_VSS_XI24/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI1/MM8 N_XI24/XI1/NET35_XI24/XI1/MM8_d N_WL<45>_XI24/XI1/MM8_g
+ N_BLN<14>_XI24/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI1/MM5 N_XI24/XI1/NET34_XI24/XI1/MM5_d N_XI24/XI1/NET33_XI24/XI1/MM5_g
+ N_VDD_XI24/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI1/MM4 N_XI24/XI1/NET33_XI24/XI1/MM4_d N_XI24/XI1/NET34_XI24/XI1/MM4_g
+ N_VDD_XI24/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI1/MM10 N_XI24/XI1/NET35_XI24/XI1/MM10_d N_XI24/XI1/NET36_XI24/XI1/MM10_g
+ N_VDD_XI24/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI1/MM11 N_XI24/XI1/NET36_XI24/XI1/MM11_d N_XI24/XI1/NET35_XI24/XI1/MM11_g
+ N_VDD_XI24/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI2/MM2 N_XI24/XI2/NET34_XI24/XI2/MM2_d N_XI24/XI2/NET33_XI24/XI2/MM2_g
+ N_VSS_XI24/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI2/MM3 N_XI24/XI2/NET33_XI24/XI2/MM3_d N_WL<44>_XI24/XI2/MM3_g
+ N_BLN<13>_XI24/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI2/MM0 N_XI24/XI2/NET34_XI24/XI2/MM0_d N_WL<44>_XI24/XI2/MM0_g
+ N_BL<13>_XI24/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI2/MM1 N_XI24/XI2/NET33_XI24/XI2/MM1_d N_XI24/XI2/NET34_XI24/XI2/MM1_g
+ N_VSS_XI24/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI2/MM9 N_XI24/XI2/NET36_XI24/XI2/MM9_d N_WL<45>_XI24/XI2/MM9_g
+ N_BL<13>_XI24/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI2/MM6 N_XI24/XI2/NET35_XI24/XI2/MM6_d N_XI24/XI2/NET36_XI24/XI2/MM6_g
+ N_VSS_XI24/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI2/MM7 N_XI24/XI2/NET36_XI24/XI2/MM7_d N_XI24/XI2/NET35_XI24/XI2/MM7_g
+ N_VSS_XI24/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI2/MM8 N_XI24/XI2/NET35_XI24/XI2/MM8_d N_WL<45>_XI24/XI2/MM8_g
+ N_BLN<13>_XI24/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI2/MM5 N_XI24/XI2/NET34_XI24/XI2/MM5_d N_XI24/XI2/NET33_XI24/XI2/MM5_g
+ N_VDD_XI24/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI2/MM4 N_XI24/XI2/NET33_XI24/XI2/MM4_d N_XI24/XI2/NET34_XI24/XI2/MM4_g
+ N_VDD_XI24/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI2/MM10 N_XI24/XI2/NET35_XI24/XI2/MM10_d N_XI24/XI2/NET36_XI24/XI2/MM10_g
+ N_VDD_XI24/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI2/MM11 N_XI24/XI2/NET36_XI24/XI2/MM11_d N_XI24/XI2/NET35_XI24/XI2/MM11_g
+ N_VDD_XI24/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI3/MM2 N_XI24/XI3/NET34_XI24/XI3/MM2_d N_XI24/XI3/NET33_XI24/XI3/MM2_g
+ N_VSS_XI24/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI3/MM3 N_XI24/XI3/NET33_XI24/XI3/MM3_d N_WL<44>_XI24/XI3/MM3_g
+ N_BLN<12>_XI24/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI3/MM0 N_XI24/XI3/NET34_XI24/XI3/MM0_d N_WL<44>_XI24/XI3/MM0_g
+ N_BL<12>_XI24/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI3/MM1 N_XI24/XI3/NET33_XI24/XI3/MM1_d N_XI24/XI3/NET34_XI24/XI3/MM1_g
+ N_VSS_XI24/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI3/MM9 N_XI24/XI3/NET36_XI24/XI3/MM9_d N_WL<45>_XI24/XI3/MM9_g
+ N_BL<12>_XI24/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI3/MM6 N_XI24/XI3/NET35_XI24/XI3/MM6_d N_XI24/XI3/NET36_XI24/XI3/MM6_g
+ N_VSS_XI24/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI3/MM7 N_XI24/XI3/NET36_XI24/XI3/MM7_d N_XI24/XI3/NET35_XI24/XI3/MM7_g
+ N_VSS_XI24/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI3/MM8 N_XI24/XI3/NET35_XI24/XI3/MM8_d N_WL<45>_XI24/XI3/MM8_g
+ N_BLN<12>_XI24/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI3/MM5 N_XI24/XI3/NET34_XI24/XI3/MM5_d N_XI24/XI3/NET33_XI24/XI3/MM5_g
+ N_VDD_XI24/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI3/MM4 N_XI24/XI3/NET33_XI24/XI3/MM4_d N_XI24/XI3/NET34_XI24/XI3/MM4_g
+ N_VDD_XI24/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI3/MM10 N_XI24/XI3/NET35_XI24/XI3/MM10_d N_XI24/XI3/NET36_XI24/XI3/MM10_g
+ N_VDD_XI24/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI3/MM11 N_XI24/XI3/NET36_XI24/XI3/MM11_d N_XI24/XI3/NET35_XI24/XI3/MM11_g
+ N_VDD_XI24/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI4/MM2 N_XI24/XI4/NET34_XI24/XI4/MM2_d N_XI24/XI4/NET33_XI24/XI4/MM2_g
+ N_VSS_XI24/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI4/MM3 N_XI24/XI4/NET33_XI24/XI4/MM3_d N_WL<44>_XI24/XI4/MM3_g
+ N_BLN<11>_XI24/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI4/MM0 N_XI24/XI4/NET34_XI24/XI4/MM0_d N_WL<44>_XI24/XI4/MM0_g
+ N_BL<11>_XI24/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI4/MM1 N_XI24/XI4/NET33_XI24/XI4/MM1_d N_XI24/XI4/NET34_XI24/XI4/MM1_g
+ N_VSS_XI24/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI4/MM9 N_XI24/XI4/NET36_XI24/XI4/MM9_d N_WL<45>_XI24/XI4/MM9_g
+ N_BL<11>_XI24/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI4/MM6 N_XI24/XI4/NET35_XI24/XI4/MM6_d N_XI24/XI4/NET36_XI24/XI4/MM6_g
+ N_VSS_XI24/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI4/MM7 N_XI24/XI4/NET36_XI24/XI4/MM7_d N_XI24/XI4/NET35_XI24/XI4/MM7_g
+ N_VSS_XI24/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI4/MM8 N_XI24/XI4/NET35_XI24/XI4/MM8_d N_WL<45>_XI24/XI4/MM8_g
+ N_BLN<11>_XI24/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI4/MM5 N_XI24/XI4/NET34_XI24/XI4/MM5_d N_XI24/XI4/NET33_XI24/XI4/MM5_g
+ N_VDD_XI24/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI4/MM4 N_XI24/XI4/NET33_XI24/XI4/MM4_d N_XI24/XI4/NET34_XI24/XI4/MM4_g
+ N_VDD_XI24/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI4/MM10 N_XI24/XI4/NET35_XI24/XI4/MM10_d N_XI24/XI4/NET36_XI24/XI4/MM10_g
+ N_VDD_XI24/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI4/MM11 N_XI24/XI4/NET36_XI24/XI4/MM11_d N_XI24/XI4/NET35_XI24/XI4/MM11_g
+ N_VDD_XI24/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI5/MM2 N_XI24/XI5/NET34_XI24/XI5/MM2_d N_XI24/XI5/NET33_XI24/XI5/MM2_g
+ N_VSS_XI24/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI5/MM3 N_XI24/XI5/NET33_XI24/XI5/MM3_d N_WL<44>_XI24/XI5/MM3_g
+ N_BLN<10>_XI24/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI5/MM0 N_XI24/XI5/NET34_XI24/XI5/MM0_d N_WL<44>_XI24/XI5/MM0_g
+ N_BL<10>_XI24/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI5/MM1 N_XI24/XI5/NET33_XI24/XI5/MM1_d N_XI24/XI5/NET34_XI24/XI5/MM1_g
+ N_VSS_XI24/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI5/MM9 N_XI24/XI5/NET36_XI24/XI5/MM9_d N_WL<45>_XI24/XI5/MM9_g
+ N_BL<10>_XI24/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI5/MM6 N_XI24/XI5/NET35_XI24/XI5/MM6_d N_XI24/XI5/NET36_XI24/XI5/MM6_g
+ N_VSS_XI24/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI5/MM7 N_XI24/XI5/NET36_XI24/XI5/MM7_d N_XI24/XI5/NET35_XI24/XI5/MM7_g
+ N_VSS_XI24/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI5/MM8 N_XI24/XI5/NET35_XI24/XI5/MM8_d N_WL<45>_XI24/XI5/MM8_g
+ N_BLN<10>_XI24/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI5/MM5 N_XI24/XI5/NET34_XI24/XI5/MM5_d N_XI24/XI5/NET33_XI24/XI5/MM5_g
+ N_VDD_XI24/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI5/MM4 N_XI24/XI5/NET33_XI24/XI5/MM4_d N_XI24/XI5/NET34_XI24/XI5/MM4_g
+ N_VDD_XI24/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI5/MM10 N_XI24/XI5/NET35_XI24/XI5/MM10_d N_XI24/XI5/NET36_XI24/XI5/MM10_g
+ N_VDD_XI24/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI5/MM11 N_XI24/XI5/NET36_XI24/XI5/MM11_d N_XI24/XI5/NET35_XI24/XI5/MM11_g
+ N_VDD_XI24/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI6/MM2 N_XI24/XI6/NET34_XI24/XI6/MM2_d N_XI24/XI6/NET33_XI24/XI6/MM2_g
+ N_VSS_XI24/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM3 N_XI24/XI6/NET33_XI24/XI6/MM3_d N_WL<44>_XI24/XI6/MM3_g
+ N_BLN<9>_XI24/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM0 N_XI24/XI6/NET34_XI24/XI6/MM0_d N_WL<44>_XI24/XI6/MM0_g
+ N_BL<9>_XI24/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM1 N_XI24/XI6/NET33_XI24/XI6/MM1_d N_XI24/XI6/NET34_XI24/XI6/MM1_g
+ N_VSS_XI24/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM9 N_XI24/XI6/NET36_XI24/XI6/MM9_d N_WL<45>_XI24/XI6/MM9_g
+ N_BL<9>_XI24/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM6 N_XI24/XI6/NET35_XI24/XI6/MM6_d N_XI24/XI6/NET36_XI24/XI6/MM6_g
+ N_VSS_XI24/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM7 N_XI24/XI6/NET36_XI24/XI6/MM7_d N_XI24/XI6/NET35_XI24/XI6/MM7_g
+ N_VSS_XI24/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM8 N_XI24/XI6/NET35_XI24/XI6/MM8_d N_WL<45>_XI24/XI6/MM8_g
+ N_BLN<9>_XI24/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI6/MM5 N_XI24/XI6/NET34_XI24/XI6/MM5_d N_XI24/XI6/NET33_XI24/XI6/MM5_g
+ N_VDD_XI24/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI6/MM4 N_XI24/XI6/NET33_XI24/XI6/MM4_d N_XI24/XI6/NET34_XI24/XI6/MM4_g
+ N_VDD_XI24/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI6/MM10 N_XI24/XI6/NET35_XI24/XI6/MM10_d N_XI24/XI6/NET36_XI24/XI6/MM10_g
+ N_VDD_XI24/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI6/MM11 N_XI24/XI6/NET36_XI24/XI6/MM11_d N_XI24/XI6/NET35_XI24/XI6/MM11_g
+ N_VDD_XI24/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI7/MM2 N_XI24/XI7/NET34_XI24/XI7/MM2_d N_XI24/XI7/NET33_XI24/XI7/MM2_g
+ N_VSS_XI24/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM3 N_XI24/XI7/NET33_XI24/XI7/MM3_d N_WL<44>_XI24/XI7/MM3_g
+ N_BLN<8>_XI24/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM0 N_XI24/XI7/NET34_XI24/XI7/MM0_d N_WL<44>_XI24/XI7/MM0_g
+ N_BL<8>_XI24/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM1 N_XI24/XI7/NET33_XI24/XI7/MM1_d N_XI24/XI7/NET34_XI24/XI7/MM1_g
+ N_VSS_XI24/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM9 N_XI24/XI7/NET36_XI24/XI7/MM9_d N_WL<45>_XI24/XI7/MM9_g
+ N_BL<8>_XI24/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM6 N_XI24/XI7/NET35_XI24/XI7/MM6_d N_XI24/XI7/NET36_XI24/XI7/MM6_g
+ N_VSS_XI24/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM7 N_XI24/XI7/NET36_XI24/XI7/MM7_d N_XI24/XI7/NET35_XI24/XI7/MM7_g
+ N_VSS_XI24/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM8 N_XI24/XI7/NET35_XI24/XI7/MM8_d N_WL<45>_XI24/XI7/MM8_g
+ N_BLN<8>_XI24/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI7/MM5 N_XI24/XI7/NET34_XI24/XI7/MM5_d N_XI24/XI7/NET33_XI24/XI7/MM5_g
+ N_VDD_XI24/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI7/MM4 N_XI24/XI7/NET33_XI24/XI7/MM4_d N_XI24/XI7/NET34_XI24/XI7/MM4_g
+ N_VDD_XI24/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI7/MM10 N_XI24/XI7/NET35_XI24/XI7/MM10_d N_XI24/XI7/NET36_XI24/XI7/MM10_g
+ N_VDD_XI24/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI7/MM11 N_XI24/XI7/NET36_XI24/XI7/MM11_d N_XI24/XI7/NET35_XI24/XI7/MM11_g
+ N_VDD_XI24/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI8/MM2 N_XI24/XI8/NET34_XI24/XI8/MM2_d N_XI24/XI8/NET33_XI24/XI8/MM2_g
+ N_VSS_XI24/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM3 N_XI24/XI8/NET33_XI24/XI8/MM3_d N_WL<44>_XI24/XI8/MM3_g
+ N_BLN<7>_XI24/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM0 N_XI24/XI8/NET34_XI24/XI8/MM0_d N_WL<44>_XI24/XI8/MM0_g
+ N_BL<7>_XI24/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM1 N_XI24/XI8/NET33_XI24/XI8/MM1_d N_XI24/XI8/NET34_XI24/XI8/MM1_g
+ N_VSS_XI24/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM9 N_XI24/XI8/NET36_XI24/XI8/MM9_d N_WL<45>_XI24/XI8/MM9_g
+ N_BL<7>_XI24/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM6 N_XI24/XI8/NET35_XI24/XI8/MM6_d N_XI24/XI8/NET36_XI24/XI8/MM6_g
+ N_VSS_XI24/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM7 N_XI24/XI8/NET36_XI24/XI8/MM7_d N_XI24/XI8/NET35_XI24/XI8/MM7_g
+ N_VSS_XI24/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM8 N_XI24/XI8/NET35_XI24/XI8/MM8_d N_WL<45>_XI24/XI8/MM8_g
+ N_BLN<7>_XI24/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI8/MM5 N_XI24/XI8/NET34_XI24/XI8/MM5_d N_XI24/XI8/NET33_XI24/XI8/MM5_g
+ N_VDD_XI24/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI8/MM4 N_XI24/XI8/NET33_XI24/XI8/MM4_d N_XI24/XI8/NET34_XI24/XI8/MM4_g
+ N_VDD_XI24/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI8/MM10 N_XI24/XI8/NET35_XI24/XI8/MM10_d N_XI24/XI8/NET36_XI24/XI8/MM10_g
+ N_VDD_XI24/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI8/MM11 N_XI24/XI8/NET36_XI24/XI8/MM11_d N_XI24/XI8/NET35_XI24/XI8/MM11_g
+ N_VDD_XI24/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI9/MM2 N_XI24/XI9/NET34_XI24/XI9/MM2_d N_XI24/XI9/NET33_XI24/XI9/MM2_g
+ N_VSS_XI24/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM3 N_XI24/XI9/NET33_XI24/XI9/MM3_d N_WL<44>_XI24/XI9/MM3_g
+ N_BLN<6>_XI24/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM0 N_XI24/XI9/NET34_XI24/XI9/MM0_d N_WL<44>_XI24/XI9/MM0_g
+ N_BL<6>_XI24/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM1 N_XI24/XI9/NET33_XI24/XI9/MM1_d N_XI24/XI9/NET34_XI24/XI9/MM1_g
+ N_VSS_XI24/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM9 N_XI24/XI9/NET36_XI24/XI9/MM9_d N_WL<45>_XI24/XI9/MM9_g
+ N_BL<6>_XI24/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM6 N_XI24/XI9/NET35_XI24/XI9/MM6_d N_XI24/XI9/NET36_XI24/XI9/MM6_g
+ N_VSS_XI24/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM7 N_XI24/XI9/NET36_XI24/XI9/MM7_d N_XI24/XI9/NET35_XI24/XI9/MM7_g
+ N_VSS_XI24/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM8 N_XI24/XI9/NET35_XI24/XI9/MM8_d N_WL<45>_XI24/XI9/MM8_g
+ N_BLN<6>_XI24/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI9/MM5 N_XI24/XI9/NET34_XI24/XI9/MM5_d N_XI24/XI9/NET33_XI24/XI9/MM5_g
+ N_VDD_XI24/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI9/MM4 N_XI24/XI9/NET33_XI24/XI9/MM4_d N_XI24/XI9/NET34_XI24/XI9/MM4_g
+ N_VDD_XI24/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI9/MM10 N_XI24/XI9/NET35_XI24/XI9/MM10_d N_XI24/XI9/NET36_XI24/XI9/MM10_g
+ N_VDD_XI24/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI9/MM11 N_XI24/XI9/NET36_XI24/XI9/MM11_d N_XI24/XI9/NET35_XI24/XI9/MM11_g
+ N_VDD_XI24/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI10/MM2 N_XI24/XI10/NET34_XI24/XI10/MM2_d
+ N_XI24/XI10/NET33_XI24/XI10/MM2_g N_VSS_XI24/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI10/MM3 N_XI24/XI10/NET33_XI24/XI10/MM3_d N_WL<44>_XI24/XI10/MM3_g
+ N_BLN<5>_XI24/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI10/MM0 N_XI24/XI10/NET34_XI24/XI10/MM0_d N_WL<44>_XI24/XI10/MM0_g
+ N_BL<5>_XI24/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI10/MM1 N_XI24/XI10/NET33_XI24/XI10/MM1_d
+ N_XI24/XI10/NET34_XI24/XI10/MM1_g N_VSS_XI24/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI10/MM9 N_XI24/XI10/NET36_XI24/XI10/MM9_d N_WL<45>_XI24/XI10/MM9_g
+ N_BL<5>_XI24/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI10/MM6 N_XI24/XI10/NET35_XI24/XI10/MM6_d
+ N_XI24/XI10/NET36_XI24/XI10/MM6_g N_VSS_XI24/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI10/MM7 N_XI24/XI10/NET36_XI24/XI10/MM7_d
+ N_XI24/XI10/NET35_XI24/XI10/MM7_g N_VSS_XI24/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI10/MM8 N_XI24/XI10/NET35_XI24/XI10/MM8_d N_WL<45>_XI24/XI10/MM8_g
+ N_BLN<5>_XI24/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI10/MM5 N_XI24/XI10/NET34_XI24/XI10/MM5_d
+ N_XI24/XI10/NET33_XI24/XI10/MM5_g N_VDD_XI24/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI10/MM4 N_XI24/XI10/NET33_XI24/XI10/MM4_d
+ N_XI24/XI10/NET34_XI24/XI10/MM4_g N_VDD_XI24/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI10/MM10 N_XI24/XI10/NET35_XI24/XI10/MM10_d
+ N_XI24/XI10/NET36_XI24/XI10/MM10_g N_VDD_XI24/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI10/MM11 N_XI24/XI10/NET36_XI24/XI10/MM11_d
+ N_XI24/XI10/NET35_XI24/XI10/MM11_g N_VDD_XI24/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI11/MM2 N_XI24/XI11/NET34_XI24/XI11/MM2_d
+ N_XI24/XI11/NET33_XI24/XI11/MM2_g N_VSS_XI24/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI11/MM3 N_XI24/XI11/NET33_XI24/XI11/MM3_d N_WL<44>_XI24/XI11/MM3_g
+ N_BLN<4>_XI24/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI11/MM0 N_XI24/XI11/NET34_XI24/XI11/MM0_d N_WL<44>_XI24/XI11/MM0_g
+ N_BL<4>_XI24/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI11/MM1 N_XI24/XI11/NET33_XI24/XI11/MM1_d
+ N_XI24/XI11/NET34_XI24/XI11/MM1_g N_VSS_XI24/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI11/MM9 N_XI24/XI11/NET36_XI24/XI11/MM9_d N_WL<45>_XI24/XI11/MM9_g
+ N_BL<4>_XI24/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI11/MM6 N_XI24/XI11/NET35_XI24/XI11/MM6_d
+ N_XI24/XI11/NET36_XI24/XI11/MM6_g N_VSS_XI24/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI11/MM7 N_XI24/XI11/NET36_XI24/XI11/MM7_d
+ N_XI24/XI11/NET35_XI24/XI11/MM7_g N_VSS_XI24/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI11/MM8 N_XI24/XI11/NET35_XI24/XI11/MM8_d N_WL<45>_XI24/XI11/MM8_g
+ N_BLN<4>_XI24/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI11/MM5 N_XI24/XI11/NET34_XI24/XI11/MM5_d
+ N_XI24/XI11/NET33_XI24/XI11/MM5_g N_VDD_XI24/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI11/MM4 N_XI24/XI11/NET33_XI24/XI11/MM4_d
+ N_XI24/XI11/NET34_XI24/XI11/MM4_g N_VDD_XI24/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI11/MM10 N_XI24/XI11/NET35_XI24/XI11/MM10_d
+ N_XI24/XI11/NET36_XI24/XI11/MM10_g N_VDD_XI24/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI11/MM11 N_XI24/XI11/NET36_XI24/XI11/MM11_d
+ N_XI24/XI11/NET35_XI24/XI11/MM11_g N_VDD_XI24/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI12/MM2 N_XI24/XI12/NET34_XI24/XI12/MM2_d
+ N_XI24/XI12/NET33_XI24/XI12/MM2_g N_VSS_XI24/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI12/MM3 N_XI24/XI12/NET33_XI24/XI12/MM3_d N_WL<44>_XI24/XI12/MM3_g
+ N_BLN<3>_XI24/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI12/MM0 N_XI24/XI12/NET34_XI24/XI12/MM0_d N_WL<44>_XI24/XI12/MM0_g
+ N_BL<3>_XI24/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI12/MM1 N_XI24/XI12/NET33_XI24/XI12/MM1_d
+ N_XI24/XI12/NET34_XI24/XI12/MM1_g N_VSS_XI24/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI12/MM9 N_XI24/XI12/NET36_XI24/XI12/MM9_d N_WL<45>_XI24/XI12/MM9_g
+ N_BL<3>_XI24/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI12/MM6 N_XI24/XI12/NET35_XI24/XI12/MM6_d
+ N_XI24/XI12/NET36_XI24/XI12/MM6_g N_VSS_XI24/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI12/MM7 N_XI24/XI12/NET36_XI24/XI12/MM7_d
+ N_XI24/XI12/NET35_XI24/XI12/MM7_g N_VSS_XI24/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI12/MM8 N_XI24/XI12/NET35_XI24/XI12/MM8_d N_WL<45>_XI24/XI12/MM8_g
+ N_BLN<3>_XI24/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI12/MM5 N_XI24/XI12/NET34_XI24/XI12/MM5_d
+ N_XI24/XI12/NET33_XI24/XI12/MM5_g N_VDD_XI24/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI12/MM4 N_XI24/XI12/NET33_XI24/XI12/MM4_d
+ N_XI24/XI12/NET34_XI24/XI12/MM4_g N_VDD_XI24/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI12/MM10 N_XI24/XI12/NET35_XI24/XI12/MM10_d
+ N_XI24/XI12/NET36_XI24/XI12/MM10_g N_VDD_XI24/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI12/MM11 N_XI24/XI12/NET36_XI24/XI12/MM11_d
+ N_XI24/XI12/NET35_XI24/XI12/MM11_g N_VDD_XI24/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI13/MM2 N_XI24/XI13/NET34_XI24/XI13/MM2_d
+ N_XI24/XI13/NET33_XI24/XI13/MM2_g N_VSS_XI24/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI13/MM3 N_XI24/XI13/NET33_XI24/XI13/MM3_d N_WL<44>_XI24/XI13/MM3_g
+ N_BLN<2>_XI24/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI13/MM0 N_XI24/XI13/NET34_XI24/XI13/MM0_d N_WL<44>_XI24/XI13/MM0_g
+ N_BL<2>_XI24/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI13/MM1 N_XI24/XI13/NET33_XI24/XI13/MM1_d
+ N_XI24/XI13/NET34_XI24/XI13/MM1_g N_VSS_XI24/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI13/MM9 N_XI24/XI13/NET36_XI24/XI13/MM9_d N_WL<45>_XI24/XI13/MM9_g
+ N_BL<2>_XI24/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI13/MM6 N_XI24/XI13/NET35_XI24/XI13/MM6_d
+ N_XI24/XI13/NET36_XI24/XI13/MM6_g N_VSS_XI24/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI13/MM7 N_XI24/XI13/NET36_XI24/XI13/MM7_d
+ N_XI24/XI13/NET35_XI24/XI13/MM7_g N_VSS_XI24/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI13/MM8 N_XI24/XI13/NET35_XI24/XI13/MM8_d N_WL<45>_XI24/XI13/MM8_g
+ N_BLN<2>_XI24/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI13/MM5 N_XI24/XI13/NET34_XI24/XI13/MM5_d
+ N_XI24/XI13/NET33_XI24/XI13/MM5_g N_VDD_XI24/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI13/MM4 N_XI24/XI13/NET33_XI24/XI13/MM4_d
+ N_XI24/XI13/NET34_XI24/XI13/MM4_g N_VDD_XI24/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI13/MM10 N_XI24/XI13/NET35_XI24/XI13/MM10_d
+ N_XI24/XI13/NET36_XI24/XI13/MM10_g N_VDD_XI24/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI13/MM11 N_XI24/XI13/NET36_XI24/XI13/MM11_d
+ N_XI24/XI13/NET35_XI24/XI13/MM11_g N_VDD_XI24/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI14/MM2 N_XI24/XI14/NET34_XI24/XI14/MM2_d
+ N_XI24/XI14/NET33_XI24/XI14/MM2_g N_VSS_XI24/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI14/MM3 N_XI24/XI14/NET33_XI24/XI14/MM3_d N_WL<44>_XI24/XI14/MM3_g
+ N_BLN<1>_XI24/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI14/MM0 N_XI24/XI14/NET34_XI24/XI14/MM0_d N_WL<44>_XI24/XI14/MM0_g
+ N_BL<1>_XI24/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI14/MM1 N_XI24/XI14/NET33_XI24/XI14/MM1_d
+ N_XI24/XI14/NET34_XI24/XI14/MM1_g N_VSS_XI24/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI14/MM9 N_XI24/XI14/NET36_XI24/XI14/MM9_d N_WL<45>_XI24/XI14/MM9_g
+ N_BL<1>_XI24/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI14/MM6 N_XI24/XI14/NET35_XI24/XI14/MM6_d
+ N_XI24/XI14/NET36_XI24/XI14/MM6_g N_VSS_XI24/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI14/MM7 N_XI24/XI14/NET36_XI24/XI14/MM7_d
+ N_XI24/XI14/NET35_XI24/XI14/MM7_g N_VSS_XI24/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI14/MM8 N_XI24/XI14/NET35_XI24/XI14/MM8_d N_WL<45>_XI24/XI14/MM8_g
+ N_BLN<1>_XI24/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI14/MM5 N_XI24/XI14/NET34_XI24/XI14/MM5_d
+ N_XI24/XI14/NET33_XI24/XI14/MM5_g N_VDD_XI24/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI14/MM4 N_XI24/XI14/NET33_XI24/XI14/MM4_d
+ N_XI24/XI14/NET34_XI24/XI14/MM4_g N_VDD_XI24/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI14/MM10 N_XI24/XI14/NET35_XI24/XI14/MM10_d
+ N_XI24/XI14/NET36_XI24/XI14/MM10_g N_VDD_XI24/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI14/MM11 N_XI24/XI14/NET36_XI24/XI14/MM11_d
+ N_XI24/XI14/NET35_XI24/XI14/MM11_g N_VDD_XI24/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI15/MM2 N_XI24/XI15/NET34_XI24/XI15/MM2_d
+ N_XI24/XI15/NET33_XI24/XI15/MM2_g N_VSS_XI24/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI15/MM3 N_XI24/XI15/NET33_XI24/XI15/MM3_d N_WL<44>_XI24/XI15/MM3_g
+ N_BLN<0>_XI24/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI15/MM0 N_XI24/XI15/NET34_XI24/XI15/MM0_d N_WL<44>_XI24/XI15/MM0_g
+ N_BL<0>_XI24/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI15/MM1 N_XI24/XI15/NET33_XI24/XI15/MM1_d
+ N_XI24/XI15/NET34_XI24/XI15/MM1_g N_VSS_XI24/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI15/MM9 N_XI24/XI15/NET36_XI24/XI15/MM9_d N_WL<45>_XI24/XI15/MM9_g
+ N_BL<0>_XI24/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI15/MM6 N_XI24/XI15/NET35_XI24/XI15/MM6_d
+ N_XI24/XI15/NET36_XI24/XI15/MM6_g N_VSS_XI24/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI15/MM7 N_XI24/XI15/NET36_XI24/XI15/MM7_d
+ N_XI24/XI15/NET35_XI24/XI15/MM7_g N_VSS_XI24/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI24/XI15/MM8 N_XI24/XI15/NET35_XI24/XI15/MM8_d N_WL<45>_XI24/XI15/MM8_g
+ N_BLN<0>_XI24/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI24/XI15/MM5 N_XI24/XI15/NET34_XI24/XI15/MM5_d
+ N_XI24/XI15/NET33_XI24/XI15/MM5_g N_VDD_XI24/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI15/MM4 N_XI24/XI15/NET33_XI24/XI15/MM4_d
+ N_XI24/XI15/NET34_XI24/XI15/MM4_g N_VDD_XI24/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI15/MM10 N_XI24/XI15/NET35_XI24/XI15/MM10_d
+ N_XI24/XI15/NET36_XI24/XI15/MM10_g N_VDD_XI24/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI24/XI15/MM11 N_XI24/XI15/NET36_XI24/XI15/MM11_d
+ N_XI24/XI15/NET35_XI24/XI15/MM11_g N_VDD_XI24/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI0/MM2 N_XI25/XI0/NET34_XI25/XI0/MM2_d N_XI25/XI0/NET33_XI25/XI0/MM2_g
+ N_VSS_XI25/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI0/MM3 N_XI25/XI0/NET33_XI25/XI0/MM3_d N_WL<46>_XI25/XI0/MM3_g
+ N_BLN<15>_XI25/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI0/MM0 N_XI25/XI0/NET34_XI25/XI0/MM0_d N_WL<46>_XI25/XI0/MM0_g
+ N_BL<15>_XI25/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI0/MM1 N_XI25/XI0/NET33_XI25/XI0/MM1_d N_XI25/XI0/NET34_XI25/XI0/MM1_g
+ N_VSS_XI25/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI0/MM9 N_XI25/XI0/NET36_XI25/XI0/MM9_d N_WL<47>_XI25/XI0/MM9_g
+ N_BL<15>_XI25/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI0/MM6 N_XI25/XI0/NET35_XI25/XI0/MM6_d N_XI25/XI0/NET36_XI25/XI0/MM6_g
+ N_VSS_XI25/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI0/MM7 N_XI25/XI0/NET36_XI25/XI0/MM7_d N_XI25/XI0/NET35_XI25/XI0/MM7_g
+ N_VSS_XI25/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI0/MM8 N_XI25/XI0/NET35_XI25/XI0/MM8_d N_WL<47>_XI25/XI0/MM8_g
+ N_BLN<15>_XI25/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI0/MM5 N_XI25/XI0/NET34_XI25/XI0/MM5_d N_XI25/XI0/NET33_XI25/XI0/MM5_g
+ N_VDD_XI25/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI0/MM4 N_XI25/XI0/NET33_XI25/XI0/MM4_d N_XI25/XI0/NET34_XI25/XI0/MM4_g
+ N_VDD_XI25/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI0/MM10 N_XI25/XI0/NET35_XI25/XI0/MM10_d N_XI25/XI0/NET36_XI25/XI0/MM10_g
+ N_VDD_XI25/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI0/MM11 N_XI25/XI0/NET36_XI25/XI0/MM11_d N_XI25/XI0/NET35_XI25/XI0/MM11_g
+ N_VDD_XI25/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI1/MM2 N_XI25/XI1/NET34_XI25/XI1/MM2_d N_XI25/XI1/NET33_XI25/XI1/MM2_g
+ N_VSS_XI25/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI1/MM3 N_XI25/XI1/NET33_XI25/XI1/MM3_d N_WL<46>_XI25/XI1/MM3_g
+ N_BLN<14>_XI25/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI1/MM0 N_XI25/XI1/NET34_XI25/XI1/MM0_d N_WL<46>_XI25/XI1/MM0_g
+ N_BL<14>_XI25/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI1/MM1 N_XI25/XI1/NET33_XI25/XI1/MM1_d N_XI25/XI1/NET34_XI25/XI1/MM1_g
+ N_VSS_XI25/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI1/MM9 N_XI25/XI1/NET36_XI25/XI1/MM9_d N_WL<47>_XI25/XI1/MM9_g
+ N_BL<14>_XI25/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI1/MM6 N_XI25/XI1/NET35_XI25/XI1/MM6_d N_XI25/XI1/NET36_XI25/XI1/MM6_g
+ N_VSS_XI25/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI1/MM7 N_XI25/XI1/NET36_XI25/XI1/MM7_d N_XI25/XI1/NET35_XI25/XI1/MM7_g
+ N_VSS_XI25/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI1/MM8 N_XI25/XI1/NET35_XI25/XI1/MM8_d N_WL<47>_XI25/XI1/MM8_g
+ N_BLN<14>_XI25/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI1/MM5 N_XI25/XI1/NET34_XI25/XI1/MM5_d N_XI25/XI1/NET33_XI25/XI1/MM5_g
+ N_VDD_XI25/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI1/MM4 N_XI25/XI1/NET33_XI25/XI1/MM4_d N_XI25/XI1/NET34_XI25/XI1/MM4_g
+ N_VDD_XI25/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI1/MM10 N_XI25/XI1/NET35_XI25/XI1/MM10_d N_XI25/XI1/NET36_XI25/XI1/MM10_g
+ N_VDD_XI25/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI1/MM11 N_XI25/XI1/NET36_XI25/XI1/MM11_d N_XI25/XI1/NET35_XI25/XI1/MM11_g
+ N_VDD_XI25/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI2/MM2 N_XI25/XI2/NET34_XI25/XI2/MM2_d N_XI25/XI2/NET33_XI25/XI2/MM2_g
+ N_VSS_XI25/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI2/MM3 N_XI25/XI2/NET33_XI25/XI2/MM3_d N_WL<46>_XI25/XI2/MM3_g
+ N_BLN<13>_XI25/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI2/MM0 N_XI25/XI2/NET34_XI25/XI2/MM0_d N_WL<46>_XI25/XI2/MM0_g
+ N_BL<13>_XI25/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI2/MM1 N_XI25/XI2/NET33_XI25/XI2/MM1_d N_XI25/XI2/NET34_XI25/XI2/MM1_g
+ N_VSS_XI25/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI2/MM9 N_XI25/XI2/NET36_XI25/XI2/MM9_d N_WL<47>_XI25/XI2/MM9_g
+ N_BL<13>_XI25/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI2/MM6 N_XI25/XI2/NET35_XI25/XI2/MM6_d N_XI25/XI2/NET36_XI25/XI2/MM6_g
+ N_VSS_XI25/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI2/MM7 N_XI25/XI2/NET36_XI25/XI2/MM7_d N_XI25/XI2/NET35_XI25/XI2/MM7_g
+ N_VSS_XI25/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI2/MM8 N_XI25/XI2/NET35_XI25/XI2/MM8_d N_WL<47>_XI25/XI2/MM8_g
+ N_BLN<13>_XI25/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI2/MM5 N_XI25/XI2/NET34_XI25/XI2/MM5_d N_XI25/XI2/NET33_XI25/XI2/MM5_g
+ N_VDD_XI25/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI2/MM4 N_XI25/XI2/NET33_XI25/XI2/MM4_d N_XI25/XI2/NET34_XI25/XI2/MM4_g
+ N_VDD_XI25/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI2/MM10 N_XI25/XI2/NET35_XI25/XI2/MM10_d N_XI25/XI2/NET36_XI25/XI2/MM10_g
+ N_VDD_XI25/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI2/MM11 N_XI25/XI2/NET36_XI25/XI2/MM11_d N_XI25/XI2/NET35_XI25/XI2/MM11_g
+ N_VDD_XI25/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI3/MM2 N_XI25/XI3/NET34_XI25/XI3/MM2_d N_XI25/XI3/NET33_XI25/XI3/MM2_g
+ N_VSS_XI25/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI3/MM3 N_XI25/XI3/NET33_XI25/XI3/MM3_d N_WL<46>_XI25/XI3/MM3_g
+ N_BLN<12>_XI25/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI3/MM0 N_XI25/XI3/NET34_XI25/XI3/MM0_d N_WL<46>_XI25/XI3/MM0_g
+ N_BL<12>_XI25/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI3/MM1 N_XI25/XI3/NET33_XI25/XI3/MM1_d N_XI25/XI3/NET34_XI25/XI3/MM1_g
+ N_VSS_XI25/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI3/MM9 N_XI25/XI3/NET36_XI25/XI3/MM9_d N_WL<47>_XI25/XI3/MM9_g
+ N_BL<12>_XI25/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI3/MM6 N_XI25/XI3/NET35_XI25/XI3/MM6_d N_XI25/XI3/NET36_XI25/XI3/MM6_g
+ N_VSS_XI25/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI3/MM7 N_XI25/XI3/NET36_XI25/XI3/MM7_d N_XI25/XI3/NET35_XI25/XI3/MM7_g
+ N_VSS_XI25/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI3/MM8 N_XI25/XI3/NET35_XI25/XI3/MM8_d N_WL<47>_XI25/XI3/MM8_g
+ N_BLN<12>_XI25/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI3/MM5 N_XI25/XI3/NET34_XI25/XI3/MM5_d N_XI25/XI3/NET33_XI25/XI3/MM5_g
+ N_VDD_XI25/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI3/MM4 N_XI25/XI3/NET33_XI25/XI3/MM4_d N_XI25/XI3/NET34_XI25/XI3/MM4_g
+ N_VDD_XI25/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI3/MM10 N_XI25/XI3/NET35_XI25/XI3/MM10_d N_XI25/XI3/NET36_XI25/XI3/MM10_g
+ N_VDD_XI25/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI3/MM11 N_XI25/XI3/NET36_XI25/XI3/MM11_d N_XI25/XI3/NET35_XI25/XI3/MM11_g
+ N_VDD_XI25/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI4/MM2 N_XI25/XI4/NET34_XI25/XI4/MM2_d N_XI25/XI4/NET33_XI25/XI4/MM2_g
+ N_VSS_XI25/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI4/MM3 N_XI25/XI4/NET33_XI25/XI4/MM3_d N_WL<46>_XI25/XI4/MM3_g
+ N_BLN<11>_XI25/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI4/MM0 N_XI25/XI4/NET34_XI25/XI4/MM0_d N_WL<46>_XI25/XI4/MM0_g
+ N_BL<11>_XI25/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI4/MM1 N_XI25/XI4/NET33_XI25/XI4/MM1_d N_XI25/XI4/NET34_XI25/XI4/MM1_g
+ N_VSS_XI25/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI4/MM9 N_XI25/XI4/NET36_XI25/XI4/MM9_d N_WL<47>_XI25/XI4/MM9_g
+ N_BL<11>_XI25/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI4/MM6 N_XI25/XI4/NET35_XI25/XI4/MM6_d N_XI25/XI4/NET36_XI25/XI4/MM6_g
+ N_VSS_XI25/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI4/MM7 N_XI25/XI4/NET36_XI25/XI4/MM7_d N_XI25/XI4/NET35_XI25/XI4/MM7_g
+ N_VSS_XI25/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI4/MM8 N_XI25/XI4/NET35_XI25/XI4/MM8_d N_WL<47>_XI25/XI4/MM8_g
+ N_BLN<11>_XI25/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI4/MM5 N_XI25/XI4/NET34_XI25/XI4/MM5_d N_XI25/XI4/NET33_XI25/XI4/MM5_g
+ N_VDD_XI25/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI4/MM4 N_XI25/XI4/NET33_XI25/XI4/MM4_d N_XI25/XI4/NET34_XI25/XI4/MM4_g
+ N_VDD_XI25/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI4/MM10 N_XI25/XI4/NET35_XI25/XI4/MM10_d N_XI25/XI4/NET36_XI25/XI4/MM10_g
+ N_VDD_XI25/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI4/MM11 N_XI25/XI4/NET36_XI25/XI4/MM11_d N_XI25/XI4/NET35_XI25/XI4/MM11_g
+ N_VDD_XI25/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI5/MM2 N_XI25/XI5/NET34_XI25/XI5/MM2_d N_XI25/XI5/NET33_XI25/XI5/MM2_g
+ N_VSS_XI25/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI5/MM3 N_XI25/XI5/NET33_XI25/XI5/MM3_d N_WL<46>_XI25/XI5/MM3_g
+ N_BLN<10>_XI25/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI5/MM0 N_XI25/XI5/NET34_XI25/XI5/MM0_d N_WL<46>_XI25/XI5/MM0_g
+ N_BL<10>_XI25/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI5/MM1 N_XI25/XI5/NET33_XI25/XI5/MM1_d N_XI25/XI5/NET34_XI25/XI5/MM1_g
+ N_VSS_XI25/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI5/MM9 N_XI25/XI5/NET36_XI25/XI5/MM9_d N_WL<47>_XI25/XI5/MM9_g
+ N_BL<10>_XI25/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI5/MM6 N_XI25/XI5/NET35_XI25/XI5/MM6_d N_XI25/XI5/NET36_XI25/XI5/MM6_g
+ N_VSS_XI25/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI5/MM7 N_XI25/XI5/NET36_XI25/XI5/MM7_d N_XI25/XI5/NET35_XI25/XI5/MM7_g
+ N_VSS_XI25/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI5/MM8 N_XI25/XI5/NET35_XI25/XI5/MM8_d N_WL<47>_XI25/XI5/MM8_g
+ N_BLN<10>_XI25/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI5/MM5 N_XI25/XI5/NET34_XI25/XI5/MM5_d N_XI25/XI5/NET33_XI25/XI5/MM5_g
+ N_VDD_XI25/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI5/MM4 N_XI25/XI5/NET33_XI25/XI5/MM4_d N_XI25/XI5/NET34_XI25/XI5/MM4_g
+ N_VDD_XI25/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI5/MM10 N_XI25/XI5/NET35_XI25/XI5/MM10_d N_XI25/XI5/NET36_XI25/XI5/MM10_g
+ N_VDD_XI25/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI5/MM11 N_XI25/XI5/NET36_XI25/XI5/MM11_d N_XI25/XI5/NET35_XI25/XI5/MM11_g
+ N_VDD_XI25/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI6/MM2 N_XI25/XI6/NET34_XI25/XI6/MM2_d N_XI25/XI6/NET33_XI25/XI6/MM2_g
+ N_VSS_XI25/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM3 N_XI25/XI6/NET33_XI25/XI6/MM3_d N_WL<46>_XI25/XI6/MM3_g
+ N_BLN<9>_XI25/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM0 N_XI25/XI6/NET34_XI25/XI6/MM0_d N_WL<46>_XI25/XI6/MM0_g
+ N_BL<9>_XI25/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM1 N_XI25/XI6/NET33_XI25/XI6/MM1_d N_XI25/XI6/NET34_XI25/XI6/MM1_g
+ N_VSS_XI25/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM9 N_XI25/XI6/NET36_XI25/XI6/MM9_d N_WL<47>_XI25/XI6/MM9_g
+ N_BL<9>_XI25/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM6 N_XI25/XI6/NET35_XI25/XI6/MM6_d N_XI25/XI6/NET36_XI25/XI6/MM6_g
+ N_VSS_XI25/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM7 N_XI25/XI6/NET36_XI25/XI6/MM7_d N_XI25/XI6/NET35_XI25/XI6/MM7_g
+ N_VSS_XI25/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM8 N_XI25/XI6/NET35_XI25/XI6/MM8_d N_WL<47>_XI25/XI6/MM8_g
+ N_BLN<9>_XI25/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI6/MM5 N_XI25/XI6/NET34_XI25/XI6/MM5_d N_XI25/XI6/NET33_XI25/XI6/MM5_g
+ N_VDD_XI25/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI6/MM4 N_XI25/XI6/NET33_XI25/XI6/MM4_d N_XI25/XI6/NET34_XI25/XI6/MM4_g
+ N_VDD_XI25/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI6/MM10 N_XI25/XI6/NET35_XI25/XI6/MM10_d N_XI25/XI6/NET36_XI25/XI6/MM10_g
+ N_VDD_XI25/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI6/MM11 N_XI25/XI6/NET36_XI25/XI6/MM11_d N_XI25/XI6/NET35_XI25/XI6/MM11_g
+ N_VDD_XI25/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI7/MM2 N_XI25/XI7/NET34_XI25/XI7/MM2_d N_XI25/XI7/NET33_XI25/XI7/MM2_g
+ N_VSS_XI25/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM3 N_XI25/XI7/NET33_XI25/XI7/MM3_d N_WL<46>_XI25/XI7/MM3_g
+ N_BLN<8>_XI25/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM0 N_XI25/XI7/NET34_XI25/XI7/MM0_d N_WL<46>_XI25/XI7/MM0_g
+ N_BL<8>_XI25/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM1 N_XI25/XI7/NET33_XI25/XI7/MM1_d N_XI25/XI7/NET34_XI25/XI7/MM1_g
+ N_VSS_XI25/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM9 N_XI25/XI7/NET36_XI25/XI7/MM9_d N_WL<47>_XI25/XI7/MM9_g
+ N_BL<8>_XI25/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM6 N_XI25/XI7/NET35_XI25/XI7/MM6_d N_XI25/XI7/NET36_XI25/XI7/MM6_g
+ N_VSS_XI25/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM7 N_XI25/XI7/NET36_XI25/XI7/MM7_d N_XI25/XI7/NET35_XI25/XI7/MM7_g
+ N_VSS_XI25/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM8 N_XI25/XI7/NET35_XI25/XI7/MM8_d N_WL<47>_XI25/XI7/MM8_g
+ N_BLN<8>_XI25/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI7/MM5 N_XI25/XI7/NET34_XI25/XI7/MM5_d N_XI25/XI7/NET33_XI25/XI7/MM5_g
+ N_VDD_XI25/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI7/MM4 N_XI25/XI7/NET33_XI25/XI7/MM4_d N_XI25/XI7/NET34_XI25/XI7/MM4_g
+ N_VDD_XI25/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI7/MM10 N_XI25/XI7/NET35_XI25/XI7/MM10_d N_XI25/XI7/NET36_XI25/XI7/MM10_g
+ N_VDD_XI25/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI7/MM11 N_XI25/XI7/NET36_XI25/XI7/MM11_d N_XI25/XI7/NET35_XI25/XI7/MM11_g
+ N_VDD_XI25/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI8/MM2 N_XI25/XI8/NET34_XI25/XI8/MM2_d N_XI25/XI8/NET33_XI25/XI8/MM2_g
+ N_VSS_XI25/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM3 N_XI25/XI8/NET33_XI25/XI8/MM3_d N_WL<46>_XI25/XI8/MM3_g
+ N_BLN<7>_XI25/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM0 N_XI25/XI8/NET34_XI25/XI8/MM0_d N_WL<46>_XI25/XI8/MM0_g
+ N_BL<7>_XI25/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM1 N_XI25/XI8/NET33_XI25/XI8/MM1_d N_XI25/XI8/NET34_XI25/XI8/MM1_g
+ N_VSS_XI25/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM9 N_XI25/XI8/NET36_XI25/XI8/MM9_d N_WL<47>_XI25/XI8/MM9_g
+ N_BL<7>_XI25/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM6 N_XI25/XI8/NET35_XI25/XI8/MM6_d N_XI25/XI8/NET36_XI25/XI8/MM6_g
+ N_VSS_XI25/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM7 N_XI25/XI8/NET36_XI25/XI8/MM7_d N_XI25/XI8/NET35_XI25/XI8/MM7_g
+ N_VSS_XI25/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM8 N_XI25/XI8/NET35_XI25/XI8/MM8_d N_WL<47>_XI25/XI8/MM8_g
+ N_BLN<7>_XI25/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI8/MM5 N_XI25/XI8/NET34_XI25/XI8/MM5_d N_XI25/XI8/NET33_XI25/XI8/MM5_g
+ N_VDD_XI25/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI8/MM4 N_XI25/XI8/NET33_XI25/XI8/MM4_d N_XI25/XI8/NET34_XI25/XI8/MM4_g
+ N_VDD_XI25/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI8/MM10 N_XI25/XI8/NET35_XI25/XI8/MM10_d N_XI25/XI8/NET36_XI25/XI8/MM10_g
+ N_VDD_XI25/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI8/MM11 N_XI25/XI8/NET36_XI25/XI8/MM11_d N_XI25/XI8/NET35_XI25/XI8/MM11_g
+ N_VDD_XI25/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI9/MM2 N_XI25/XI9/NET34_XI25/XI9/MM2_d N_XI25/XI9/NET33_XI25/XI9/MM2_g
+ N_VSS_XI25/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM3 N_XI25/XI9/NET33_XI25/XI9/MM3_d N_WL<46>_XI25/XI9/MM3_g
+ N_BLN<6>_XI25/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM0 N_XI25/XI9/NET34_XI25/XI9/MM0_d N_WL<46>_XI25/XI9/MM0_g
+ N_BL<6>_XI25/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM1 N_XI25/XI9/NET33_XI25/XI9/MM1_d N_XI25/XI9/NET34_XI25/XI9/MM1_g
+ N_VSS_XI25/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM9 N_XI25/XI9/NET36_XI25/XI9/MM9_d N_WL<47>_XI25/XI9/MM9_g
+ N_BL<6>_XI25/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM6 N_XI25/XI9/NET35_XI25/XI9/MM6_d N_XI25/XI9/NET36_XI25/XI9/MM6_g
+ N_VSS_XI25/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM7 N_XI25/XI9/NET36_XI25/XI9/MM7_d N_XI25/XI9/NET35_XI25/XI9/MM7_g
+ N_VSS_XI25/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM8 N_XI25/XI9/NET35_XI25/XI9/MM8_d N_WL<47>_XI25/XI9/MM8_g
+ N_BLN<6>_XI25/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI9/MM5 N_XI25/XI9/NET34_XI25/XI9/MM5_d N_XI25/XI9/NET33_XI25/XI9/MM5_g
+ N_VDD_XI25/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI9/MM4 N_XI25/XI9/NET33_XI25/XI9/MM4_d N_XI25/XI9/NET34_XI25/XI9/MM4_g
+ N_VDD_XI25/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI9/MM10 N_XI25/XI9/NET35_XI25/XI9/MM10_d N_XI25/XI9/NET36_XI25/XI9/MM10_g
+ N_VDD_XI25/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI9/MM11 N_XI25/XI9/NET36_XI25/XI9/MM11_d N_XI25/XI9/NET35_XI25/XI9/MM11_g
+ N_VDD_XI25/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI10/MM2 N_XI25/XI10/NET34_XI25/XI10/MM2_d
+ N_XI25/XI10/NET33_XI25/XI10/MM2_g N_VSS_XI25/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI10/MM3 N_XI25/XI10/NET33_XI25/XI10/MM3_d N_WL<46>_XI25/XI10/MM3_g
+ N_BLN<5>_XI25/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI10/MM0 N_XI25/XI10/NET34_XI25/XI10/MM0_d N_WL<46>_XI25/XI10/MM0_g
+ N_BL<5>_XI25/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI10/MM1 N_XI25/XI10/NET33_XI25/XI10/MM1_d
+ N_XI25/XI10/NET34_XI25/XI10/MM1_g N_VSS_XI25/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI10/MM9 N_XI25/XI10/NET36_XI25/XI10/MM9_d N_WL<47>_XI25/XI10/MM9_g
+ N_BL<5>_XI25/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI10/MM6 N_XI25/XI10/NET35_XI25/XI10/MM6_d
+ N_XI25/XI10/NET36_XI25/XI10/MM6_g N_VSS_XI25/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI10/MM7 N_XI25/XI10/NET36_XI25/XI10/MM7_d
+ N_XI25/XI10/NET35_XI25/XI10/MM7_g N_VSS_XI25/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI10/MM8 N_XI25/XI10/NET35_XI25/XI10/MM8_d N_WL<47>_XI25/XI10/MM8_g
+ N_BLN<5>_XI25/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI10/MM5 N_XI25/XI10/NET34_XI25/XI10/MM5_d
+ N_XI25/XI10/NET33_XI25/XI10/MM5_g N_VDD_XI25/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI10/MM4 N_XI25/XI10/NET33_XI25/XI10/MM4_d
+ N_XI25/XI10/NET34_XI25/XI10/MM4_g N_VDD_XI25/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI10/MM10 N_XI25/XI10/NET35_XI25/XI10/MM10_d
+ N_XI25/XI10/NET36_XI25/XI10/MM10_g N_VDD_XI25/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI10/MM11 N_XI25/XI10/NET36_XI25/XI10/MM11_d
+ N_XI25/XI10/NET35_XI25/XI10/MM11_g N_VDD_XI25/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI11/MM2 N_XI25/XI11/NET34_XI25/XI11/MM2_d
+ N_XI25/XI11/NET33_XI25/XI11/MM2_g N_VSS_XI25/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI11/MM3 N_XI25/XI11/NET33_XI25/XI11/MM3_d N_WL<46>_XI25/XI11/MM3_g
+ N_BLN<4>_XI25/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI11/MM0 N_XI25/XI11/NET34_XI25/XI11/MM0_d N_WL<46>_XI25/XI11/MM0_g
+ N_BL<4>_XI25/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI11/MM1 N_XI25/XI11/NET33_XI25/XI11/MM1_d
+ N_XI25/XI11/NET34_XI25/XI11/MM1_g N_VSS_XI25/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI11/MM9 N_XI25/XI11/NET36_XI25/XI11/MM9_d N_WL<47>_XI25/XI11/MM9_g
+ N_BL<4>_XI25/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI11/MM6 N_XI25/XI11/NET35_XI25/XI11/MM6_d
+ N_XI25/XI11/NET36_XI25/XI11/MM6_g N_VSS_XI25/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI11/MM7 N_XI25/XI11/NET36_XI25/XI11/MM7_d
+ N_XI25/XI11/NET35_XI25/XI11/MM7_g N_VSS_XI25/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI11/MM8 N_XI25/XI11/NET35_XI25/XI11/MM8_d N_WL<47>_XI25/XI11/MM8_g
+ N_BLN<4>_XI25/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI11/MM5 N_XI25/XI11/NET34_XI25/XI11/MM5_d
+ N_XI25/XI11/NET33_XI25/XI11/MM5_g N_VDD_XI25/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI11/MM4 N_XI25/XI11/NET33_XI25/XI11/MM4_d
+ N_XI25/XI11/NET34_XI25/XI11/MM4_g N_VDD_XI25/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI11/MM10 N_XI25/XI11/NET35_XI25/XI11/MM10_d
+ N_XI25/XI11/NET36_XI25/XI11/MM10_g N_VDD_XI25/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI11/MM11 N_XI25/XI11/NET36_XI25/XI11/MM11_d
+ N_XI25/XI11/NET35_XI25/XI11/MM11_g N_VDD_XI25/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI12/MM2 N_XI25/XI12/NET34_XI25/XI12/MM2_d
+ N_XI25/XI12/NET33_XI25/XI12/MM2_g N_VSS_XI25/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI12/MM3 N_XI25/XI12/NET33_XI25/XI12/MM3_d N_WL<46>_XI25/XI12/MM3_g
+ N_BLN<3>_XI25/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI12/MM0 N_XI25/XI12/NET34_XI25/XI12/MM0_d N_WL<46>_XI25/XI12/MM0_g
+ N_BL<3>_XI25/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI12/MM1 N_XI25/XI12/NET33_XI25/XI12/MM1_d
+ N_XI25/XI12/NET34_XI25/XI12/MM1_g N_VSS_XI25/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI12/MM9 N_XI25/XI12/NET36_XI25/XI12/MM9_d N_WL<47>_XI25/XI12/MM9_g
+ N_BL<3>_XI25/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI12/MM6 N_XI25/XI12/NET35_XI25/XI12/MM6_d
+ N_XI25/XI12/NET36_XI25/XI12/MM6_g N_VSS_XI25/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI12/MM7 N_XI25/XI12/NET36_XI25/XI12/MM7_d
+ N_XI25/XI12/NET35_XI25/XI12/MM7_g N_VSS_XI25/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI12/MM8 N_XI25/XI12/NET35_XI25/XI12/MM8_d N_WL<47>_XI25/XI12/MM8_g
+ N_BLN<3>_XI25/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI12/MM5 N_XI25/XI12/NET34_XI25/XI12/MM5_d
+ N_XI25/XI12/NET33_XI25/XI12/MM5_g N_VDD_XI25/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI12/MM4 N_XI25/XI12/NET33_XI25/XI12/MM4_d
+ N_XI25/XI12/NET34_XI25/XI12/MM4_g N_VDD_XI25/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI12/MM10 N_XI25/XI12/NET35_XI25/XI12/MM10_d
+ N_XI25/XI12/NET36_XI25/XI12/MM10_g N_VDD_XI25/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI12/MM11 N_XI25/XI12/NET36_XI25/XI12/MM11_d
+ N_XI25/XI12/NET35_XI25/XI12/MM11_g N_VDD_XI25/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI13/MM2 N_XI25/XI13/NET34_XI25/XI13/MM2_d
+ N_XI25/XI13/NET33_XI25/XI13/MM2_g N_VSS_XI25/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI13/MM3 N_XI25/XI13/NET33_XI25/XI13/MM3_d N_WL<46>_XI25/XI13/MM3_g
+ N_BLN<2>_XI25/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI13/MM0 N_XI25/XI13/NET34_XI25/XI13/MM0_d N_WL<46>_XI25/XI13/MM0_g
+ N_BL<2>_XI25/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI13/MM1 N_XI25/XI13/NET33_XI25/XI13/MM1_d
+ N_XI25/XI13/NET34_XI25/XI13/MM1_g N_VSS_XI25/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI13/MM9 N_XI25/XI13/NET36_XI25/XI13/MM9_d N_WL<47>_XI25/XI13/MM9_g
+ N_BL<2>_XI25/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI13/MM6 N_XI25/XI13/NET35_XI25/XI13/MM6_d
+ N_XI25/XI13/NET36_XI25/XI13/MM6_g N_VSS_XI25/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI13/MM7 N_XI25/XI13/NET36_XI25/XI13/MM7_d
+ N_XI25/XI13/NET35_XI25/XI13/MM7_g N_VSS_XI25/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI13/MM8 N_XI25/XI13/NET35_XI25/XI13/MM8_d N_WL<47>_XI25/XI13/MM8_g
+ N_BLN<2>_XI25/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI13/MM5 N_XI25/XI13/NET34_XI25/XI13/MM5_d
+ N_XI25/XI13/NET33_XI25/XI13/MM5_g N_VDD_XI25/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI13/MM4 N_XI25/XI13/NET33_XI25/XI13/MM4_d
+ N_XI25/XI13/NET34_XI25/XI13/MM4_g N_VDD_XI25/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI13/MM10 N_XI25/XI13/NET35_XI25/XI13/MM10_d
+ N_XI25/XI13/NET36_XI25/XI13/MM10_g N_VDD_XI25/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI13/MM11 N_XI25/XI13/NET36_XI25/XI13/MM11_d
+ N_XI25/XI13/NET35_XI25/XI13/MM11_g N_VDD_XI25/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI14/MM2 N_XI25/XI14/NET34_XI25/XI14/MM2_d
+ N_XI25/XI14/NET33_XI25/XI14/MM2_g N_VSS_XI25/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI14/MM3 N_XI25/XI14/NET33_XI25/XI14/MM3_d N_WL<46>_XI25/XI14/MM3_g
+ N_BLN<1>_XI25/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI14/MM0 N_XI25/XI14/NET34_XI25/XI14/MM0_d N_WL<46>_XI25/XI14/MM0_g
+ N_BL<1>_XI25/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI14/MM1 N_XI25/XI14/NET33_XI25/XI14/MM1_d
+ N_XI25/XI14/NET34_XI25/XI14/MM1_g N_VSS_XI25/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI14/MM9 N_XI25/XI14/NET36_XI25/XI14/MM9_d N_WL<47>_XI25/XI14/MM9_g
+ N_BL<1>_XI25/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI14/MM6 N_XI25/XI14/NET35_XI25/XI14/MM6_d
+ N_XI25/XI14/NET36_XI25/XI14/MM6_g N_VSS_XI25/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI14/MM7 N_XI25/XI14/NET36_XI25/XI14/MM7_d
+ N_XI25/XI14/NET35_XI25/XI14/MM7_g N_VSS_XI25/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI14/MM8 N_XI25/XI14/NET35_XI25/XI14/MM8_d N_WL<47>_XI25/XI14/MM8_g
+ N_BLN<1>_XI25/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI14/MM5 N_XI25/XI14/NET34_XI25/XI14/MM5_d
+ N_XI25/XI14/NET33_XI25/XI14/MM5_g N_VDD_XI25/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI14/MM4 N_XI25/XI14/NET33_XI25/XI14/MM4_d
+ N_XI25/XI14/NET34_XI25/XI14/MM4_g N_VDD_XI25/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI14/MM10 N_XI25/XI14/NET35_XI25/XI14/MM10_d
+ N_XI25/XI14/NET36_XI25/XI14/MM10_g N_VDD_XI25/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI14/MM11 N_XI25/XI14/NET36_XI25/XI14/MM11_d
+ N_XI25/XI14/NET35_XI25/XI14/MM11_g N_VDD_XI25/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI15/MM2 N_XI25/XI15/NET34_XI25/XI15/MM2_d
+ N_XI25/XI15/NET33_XI25/XI15/MM2_g N_VSS_XI25/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI15/MM3 N_XI25/XI15/NET33_XI25/XI15/MM3_d N_WL<46>_XI25/XI15/MM3_g
+ N_BLN<0>_XI25/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI15/MM0 N_XI25/XI15/NET34_XI25/XI15/MM0_d N_WL<46>_XI25/XI15/MM0_g
+ N_BL<0>_XI25/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI15/MM1 N_XI25/XI15/NET33_XI25/XI15/MM1_d
+ N_XI25/XI15/NET34_XI25/XI15/MM1_g N_VSS_XI25/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI15/MM9 N_XI25/XI15/NET36_XI25/XI15/MM9_d N_WL<47>_XI25/XI15/MM9_g
+ N_BL<0>_XI25/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI15/MM6 N_XI25/XI15/NET35_XI25/XI15/MM6_d
+ N_XI25/XI15/NET36_XI25/XI15/MM6_g N_VSS_XI25/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI15/MM7 N_XI25/XI15/NET36_XI25/XI15/MM7_d
+ N_XI25/XI15/NET35_XI25/XI15/MM7_g N_VSS_XI25/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI25/XI15/MM8 N_XI25/XI15/NET35_XI25/XI15/MM8_d N_WL<47>_XI25/XI15/MM8_g
+ N_BLN<0>_XI25/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI25/XI15/MM5 N_XI25/XI15/NET34_XI25/XI15/MM5_d
+ N_XI25/XI15/NET33_XI25/XI15/MM5_g N_VDD_XI25/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI15/MM4 N_XI25/XI15/NET33_XI25/XI15/MM4_d
+ N_XI25/XI15/NET34_XI25/XI15/MM4_g N_VDD_XI25/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI15/MM10 N_XI25/XI15/NET35_XI25/XI15/MM10_d
+ N_XI25/XI15/NET36_XI25/XI15/MM10_g N_VDD_XI25/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI25/XI15/MM11 N_XI25/XI15/NET36_XI25/XI15/MM11_d
+ N_XI25/XI15/NET35_XI25/XI15/MM11_g N_VDD_XI25/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI0/MM2 N_XI26/XI0/NET34_XI26/XI0/MM2_d N_XI26/XI0/NET33_XI26/XI0/MM2_g
+ N_VSS_XI26/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI0/MM3 N_XI26/XI0/NET33_XI26/XI0/MM3_d N_WL<48>_XI26/XI0/MM3_g
+ N_BLN<15>_XI26/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI0/MM0 N_XI26/XI0/NET34_XI26/XI0/MM0_d N_WL<48>_XI26/XI0/MM0_g
+ N_BL<15>_XI26/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI0/MM1 N_XI26/XI0/NET33_XI26/XI0/MM1_d N_XI26/XI0/NET34_XI26/XI0/MM1_g
+ N_VSS_XI26/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI0/MM9 N_XI26/XI0/NET36_XI26/XI0/MM9_d N_WL<49>_XI26/XI0/MM9_g
+ N_BL<15>_XI26/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI0/MM6 N_XI26/XI0/NET35_XI26/XI0/MM6_d N_XI26/XI0/NET36_XI26/XI0/MM6_g
+ N_VSS_XI26/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI0/MM7 N_XI26/XI0/NET36_XI26/XI0/MM7_d N_XI26/XI0/NET35_XI26/XI0/MM7_g
+ N_VSS_XI26/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI0/MM8 N_XI26/XI0/NET35_XI26/XI0/MM8_d N_WL<49>_XI26/XI0/MM8_g
+ N_BLN<15>_XI26/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI0/MM5 N_XI26/XI0/NET34_XI26/XI0/MM5_d N_XI26/XI0/NET33_XI26/XI0/MM5_g
+ N_VDD_XI26/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI0/MM4 N_XI26/XI0/NET33_XI26/XI0/MM4_d N_XI26/XI0/NET34_XI26/XI0/MM4_g
+ N_VDD_XI26/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI0/MM10 N_XI26/XI0/NET35_XI26/XI0/MM10_d N_XI26/XI0/NET36_XI26/XI0/MM10_g
+ N_VDD_XI26/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI0/MM11 N_XI26/XI0/NET36_XI26/XI0/MM11_d N_XI26/XI0/NET35_XI26/XI0/MM11_g
+ N_VDD_XI26/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI1/MM2 N_XI26/XI1/NET34_XI26/XI1/MM2_d N_XI26/XI1/NET33_XI26/XI1/MM2_g
+ N_VSS_XI26/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI1/MM3 N_XI26/XI1/NET33_XI26/XI1/MM3_d N_WL<48>_XI26/XI1/MM3_g
+ N_BLN<14>_XI26/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI1/MM0 N_XI26/XI1/NET34_XI26/XI1/MM0_d N_WL<48>_XI26/XI1/MM0_g
+ N_BL<14>_XI26/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI1/MM1 N_XI26/XI1/NET33_XI26/XI1/MM1_d N_XI26/XI1/NET34_XI26/XI1/MM1_g
+ N_VSS_XI26/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI1/MM9 N_XI26/XI1/NET36_XI26/XI1/MM9_d N_WL<49>_XI26/XI1/MM9_g
+ N_BL<14>_XI26/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI1/MM6 N_XI26/XI1/NET35_XI26/XI1/MM6_d N_XI26/XI1/NET36_XI26/XI1/MM6_g
+ N_VSS_XI26/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI1/MM7 N_XI26/XI1/NET36_XI26/XI1/MM7_d N_XI26/XI1/NET35_XI26/XI1/MM7_g
+ N_VSS_XI26/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI1/MM8 N_XI26/XI1/NET35_XI26/XI1/MM8_d N_WL<49>_XI26/XI1/MM8_g
+ N_BLN<14>_XI26/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI1/MM5 N_XI26/XI1/NET34_XI26/XI1/MM5_d N_XI26/XI1/NET33_XI26/XI1/MM5_g
+ N_VDD_XI26/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI1/MM4 N_XI26/XI1/NET33_XI26/XI1/MM4_d N_XI26/XI1/NET34_XI26/XI1/MM4_g
+ N_VDD_XI26/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI1/MM10 N_XI26/XI1/NET35_XI26/XI1/MM10_d N_XI26/XI1/NET36_XI26/XI1/MM10_g
+ N_VDD_XI26/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI1/MM11 N_XI26/XI1/NET36_XI26/XI1/MM11_d N_XI26/XI1/NET35_XI26/XI1/MM11_g
+ N_VDD_XI26/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI2/MM2 N_XI26/XI2/NET34_XI26/XI2/MM2_d N_XI26/XI2/NET33_XI26/XI2/MM2_g
+ N_VSS_XI26/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI2/MM3 N_XI26/XI2/NET33_XI26/XI2/MM3_d N_WL<48>_XI26/XI2/MM3_g
+ N_BLN<13>_XI26/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI2/MM0 N_XI26/XI2/NET34_XI26/XI2/MM0_d N_WL<48>_XI26/XI2/MM0_g
+ N_BL<13>_XI26/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI2/MM1 N_XI26/XI2/NET33_XI26/XI2/MM1_d N_XI26/XI2/NET34_XI26/XI2/MM1_g
+ N_VSS_XI26/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI2/MM9 N_XI26/XI2/NET36_XI26/XI2/MM9_d N_WL<49>_XI26/XI2/MM9_g
+ N_BL<13>_XI26/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI2/MM6 N_XI26/XI2/NET35_XI26/XI2/MM6_d N_XI26/XI2/NET36_XI26/XI2/MM6_g
+ N_VSS_XI26/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI2/MM7 N_XI26/XI2/NET36_XI26/XI2/MM7_d N_XI26/XI2/NET35_XI26/XI2/MM7_g
+ N_VSS_XI26/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI2/MM8 N_XI26/XI2/NET35_XI26/XI2/MM8_d N_WL<49>_XI26/XI2/MM8_g
+ N_BLN<13>_XI26/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI2/MM5 N_XI26/XI2/NET34_XI26/XI2/MM5_d N_XI26/XI2/NET33_XI26/XI2/MM5_g
+ N_VDD_XI26/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI2/MM4 N_XI26/XI2/NET33_XI26/XI2/MM4_d N_XI26/XI2/NET34_XI26/XI2/MM4_g
+ N_VDD_XI26/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI2/MM10 N_XI26/XI2/NET35_XI26/XI2/MM10_d N_XI26/XI2/NET36_XI26/XI2/MM10_g
+ N_VDD_XI26/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI2/MM11 N_XI26/XI2/NET36_XI26/XI2/MM11_d N_XI26/XI2/NET35_XI26/XI2/MM11_g
+ N_VDD_XI26/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI3/MM2 N_XI26/XI3/NET34_XI26/XI3/MM2_d N_XI26/XI3/NET33_XI26/XI3/MM2_g
+ N_VSS_XI26/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI3/MM3 N_XI26/XI3/NET33_XI26/XI3/MM3_d N_WL<48>_XI26/XI3/MM3_g
+ N_BLN<12>_XI26/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI3/MM0 N_XI26/XI3/NET34_XI26/XI3/MM0_d N_WL<48>_XI26/XI3/MM0_g
+ N_BL<12>_XI26/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI3/MM1 N_XI26/XI3/NET33_XI26/XI3/MM1_d N_XI26/XI3/NET34_XI26/XI3/MM1_g
+ N_VSS_XI26/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI3/MM9 N_XI26/XI3/NET36_XI26/XI3/MM9_d N_WL<49>_XI26/XI3/MM9_g
+ N_BL<12>_XI26/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI3/MM6 N_XI26/XI3/NET35_XI26/XI3/MM6_d N_XI26/XI3/NET36_XI26/XI3/MM6_g
+ N_VSS_XI26/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI3/MM7 N_XI26/XI3/NET36_XI26/XI3/MM7_d N_XI26/XI3/NET35_XI26/XI3/MM7_g
+ N_VSS_XI26/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI3/MM8 N_XI26/XI3/NET35_XI26/XI3/MM8_d N_WL<49>_XI26/XI3/MM8_g
+ N_BLN<12>_XI26/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI3/MM5 N_XI26/XI3/NET34_XI26/XI3/MM5_d N_XI26/XI3/NET33_XI26/XI3/MM5_g
+ N_VDD_XI26/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI3/MM4 N_XI26/XI3/NET33_XI26/XI3/MM4_d N_XI26/XI3/NET34_XI26/XI3/MM4_g
+ N_VDD_XI26/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI3/MM10 N_XI26/XI3/NET35_XI26/XI3/MM10_d N_XI26/XI3/NET36_XI26/XI3/MM10_g
+ N_VDD_XI26/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI3/MM11 N_XI26/XI3/NET36_XI26/XI3/MM11_d N_XI26/XI3/NET35_XI26/XI3/MM11_g
+ N_VDD_XI26/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI4/MM2 N_XI26/XI4/NET34_XI26/XI4/MM2_d N_XI26/XI4/NET33_XI26/XI4/MM2_g
+ N_VSS_XI26/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI4/MM3 N_XI26/XI4/NET33_XI26/XI4/MM3_d N_WL<48>_XI26/XI4/MM3_g
+ N_BLN<11>_XI26/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI4/MM0 N_XI26/XI4/NET34_XI26/XI4/MM0_d N_WL<48>_XI26/XI4/MM0_g
+ N_BL<11>_XI26/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI4/MM1 N_XI26/XI4/NET33_XI26/XI4/MM1_d N_XI26/XI4/NET34_XI26/XI4/MM1_g
+ N_VSS_XI26/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI4/MM9 N_XI26/XI4/NET36_XI26/XI4/MM9_d N_WL<49>_XI26/XI4/MM9_g
+ N_BL<11>_XI26/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI4/MM6 N_XI26/XI4/NET35_XI26/XI4/MM6_d N_XI26/XI4/NET36_XI26/XI4/MM6_g
+ N_VSS_XI26/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI4/MM7 N_XI26/XI4/NET36_XI26/XI4/MM7_d N_XI26/XI4/NET35_XI26/XI4/MM7_g
+ N_VSS_XI26/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI4/MM8 N_XI26/XI4/NET35_XI26/XI4/MM8_d N_WL<49>_XI26/XI4/MM8_g
+ N_BLN<11>_XI26/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI4/MM5 N_XI26/XI4/NET34_XI26/XI4/MM5_d N_XI26/XI4/NET33_XI26/XI4/MM5_g
+ N_VDD_XI26/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI4/MM4 N_XI26/XI4/NET33_XI26/XI4/MM4_d N_XI26/XI4/NET34_XI26/XI4/MM4_g
+ N_VDD_XI26/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI4/MM10 N_XI26/XI4/NET35_XI26/XI4/MM10_d N_XI26/XI4/NET36_XI26/XI4/MM10_g
+ N_VDD_XI26/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI4/MM11 N_XI26/XI4/NET36_XI26/XI4/MM11_d N_XI26/XI4/NET35_XI26/XI4/MM11_g
+ N_VDD_XI26/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI5/MM2 N_XI26/XI5/NET34_XI26/XI5/MM2_d N_XI26/XI5/NET33_XI26/XI5/MM2_g
+ N_VSS_XI26/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI5/MM3 N_XI26/XI5/NET33_XI26/XI5/MM3_d N_WL<48>_XI26/XI5/MM3_g
+ N_BLN<10>_XI26/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI5/MM0 N_XI26/XI5/NET34_XI26/XI5/MM0_d N_WL<48>_XI26/XI5/MM0_g
+ N_BL<10>_XI26/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI5/MM1 N_XI26/XI5/NET33_XI26/XI5/MM1_d N_XI26/XI5/NET34_XI26/XI5/MM1_g
+ N_VSS_XI26/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI5/MM9 N_XI26/XI5/NET36_XI26/XI5/MM9_d N_WL<49>_XI26/XI5/MM9_g
+ N_BL<10>_XI26/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI5/MM6 N_XI26/XI5/NET35_XI26/XI5/MM6_d N_XI26/XI5/NET36_XI26/XI5/MM6_g
+ N_VSS_XI26/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI5/MM7 N_XI26/XI5/NET36_XI26/XI5/MM7_d N_XI26/XI5/NET35_XI26/XI5/MM7_g
+ N_VSS_XI26/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI5/MM8 N_XI26/XI5/NET35_XI26/XI5/MM8_d N_WL<49>_XI26/XI5/MM8_g
+ N_BLN<10>_XI26/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI5/MM5 N_XI26/XI5/NET34_XI26/XI5/MM5_d N_XI26/XI5/NET33_XI26/XI5/MM5_g
+ N_VDD_XI26/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI5/MM4 N_XI26/XI5/NET33_XI26/XI5/MM4_d N_XI26/XI5/NET34_XI26/XI5/MM4_g
+ N_VDD_XI26/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI5/MM10 N_XI26/XI5/NET35_XI26/XI5/MM10_d N_XI26/XI5/NET36_XI26/XI5/MM10_g
+ N_VDD_XI26/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI5/MM11 N_XI26/XI5/NET36_XI26/XI5/MM11_d N_XI26/XI5/NET35_XI26/XI5/MM11_g
+ N_VDD_XI26/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI6/MM2 N_XI26/XI6/NET34_XI26/XI6/MM2_d N_XI26/XI6/NET33_XI26/XI6/MM2_g
+ N_VSS_XI26/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM3 N_XI26/XI6/NET33_XI26/XI6/MM3_d N_WL<48>_XI26/XI6/MM3_g
+ N_BLN<9>_XI26/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM0 N_XI26/XI6/NET34_XI26/XI6/MM0_d N_WL<48>_XI26/XI6/MM0_g
+ N_BL<9>_XI26/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM1 N_XI26/XI6/NET33_XI26/XI6/MM1_d N_XI26/XI6/NET34_XI26/XI6/MM1_g
+ N_VSS_XI26/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM9 N_XI26/XI6/NET36_XI26/XI6/MM9_d N_WL<49>_XI26/XI6/MM9_g
+ N_BL<9>_XI26/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM6 N_XI26/XI6/NET35_XI26/XI6/MM6_d N_XI26/XI6/NET36_XI26/XI6/MM6_g
+ N_VSS_XI26/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM7 N_XI26/XI6/NET36_XI26/XI6/MM7_d N_XI26/XI6/NET35_XI26/XI6/MM7_g
+ N_VSS_XI26/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM8 N_XI26/XI6/NET35_XI26/XI6/MM8_d N_WL<49>_XI26/XI6/MM8_g
+ N_BLN<9>_XI26/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI6/MM5 N_XI26/XI6/NET34_XI26/XI6/MM5_d N_XI26/XI6/NET33_XI26/XI6/MM5_g
+ N_VDD_XI26/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI6/MM4 N_XI26/XI6/NET33_XI26/XI6/MM4_d N_XI26/XI6/NET34_XI26/XI6/MM4_g
+ N_VDD_XI26/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI6/MM10 N_XI26/XI6/NET35_XI26/XI6/MM10_d N_XI26/XI6/NET36_XI26/XI6/MM10_g
+ N_VDD_XI26/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI6/MM11 N_XI26/XI6/NET36_XI26/XI6/MM11_d N_XI26/XI6/NET35_XI26/XI6/MM11_g
+ N_VDD_XI26/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI7/MM2 N_XI26/XI7/NET34_XI26/XI7/MM2_d N_XI26/XI7/NET33_XI26/XI7/MM2_g
+ N_VSS_XI26/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM3 N_XI26/XI7/NET33_XI26/XI7/MM3_d N_WL<48>_XI26/XI7/MM3_g
+ N_BLN<8>_XI26/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM0 N_XI26/XI7/NET34_XI26/XI7/MM0_d N_WL<48>_XI26/XI7/MM0_g
+ N_BL<8>_XI26/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM1 N_XI26/XI7/NET33_XI26/XI7/MM1_d N_XI26/XI7/NET34_XI26/XI7/MM1_g
+ N_VSS_XI26/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM9 N_XI26/XI7/NET36_XI26/XI7/MM9_d N_WL<49>_XI26/XI7/MM9_g
+ N_BL<8>_XI26/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM6 N_XI26/XI7/NET35_XI26/XI7/MM6_d N_XI26/XI7/NET36_XI26/XI7/MM6_g
+ N_VSS_XI26/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM7 N_XI26/XI7/NET36_XI26/XI7/MM7_d N_XI26/XI7/NET35_XI26/XI7/MM7_g
+ N_VSS_XI26/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM8 N_XI26/XI7/NET35_XI26/XI7/MM8_d N_WL<49>_XI26/XI7/MM8_g
+ N_BLN<8>_XI26/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI7/MM5 N_XI26/XI7/NET34_XI26/XI7/MM5_d N_XI26/XI7/NET33_XI26/XI7/MM5_g
+ N_VDD_XI26/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI7/MM4 N_XI26/XI7/NET33_XI26/XI7/MM4_d N_XI26/XI7/NET34_XI26/XI7/MM4_g
+ N_VDD_XI26/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI7/MM10 N_XI26/XI7/NET35_XI26/XI7/MM10_d N_XI26/XI7/NET36_XI26/XI7/MM10_g
+ N_VDD_XI26/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI7/MM11 N_XI26/XI7/NET36_XI26/XI7/MM11_d N_XI26/XI7/NET35_XI26/XI7/MM11_g
+ N_VDD_XI26/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI8/MM2 N_XI26/XI8/NET34_XI26/XI8/MM2_d N_XI26/XI8/NET33_XI26/XI8/MM2_g
+ N_VSS_XI26/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM3 N_XI26/XI8/NET33_XI26/XI8/MM3_d N_WL<48>_XI26/XI8/MM3_g
+ N_BLN<7>_XI26/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM0 N_XI26/XI8/NET34_XI26/XI8/MM0_d N_WL<48>_XI26/XI8/MM0_g
+ N_BL<7>_XI26/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM1 N_XI26/XI8/NET33_XI26/XI8/MM1_d N_XI26/XI8/NET34_XI26/XI8/MM1_g
+ N_VSS_XI26/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM9 N_XI26/XI8/NET36_XI26/XI8/MM9_d N_WL<49>_XI26/XI8/MM9_g
+ N_BL<7>_XI26/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM6 N_XI26/XI8/NET35_XI26/XI8/MM6_d N_XI26/XI8/NET36_XI26/XI8/MM6_g
+ N_VSS_XI26/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM7 N_XI26/XI8/NET36_XI26/XI8/MM7_d N_XI26/XI8/NET35_XI26/XI8/MM7_g
+ N_VSS_XI26/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM8 N_XI26/XI8/NET35_XI26/XI8/MM8_d N_WL<49>_XI26/XI8/MM8_g
+ N_BLN<7>_XI26/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI8/MM5 N_XI26/XI8/NET34_XI26/XI8/MM5_d N_XI26/XI8/NET33_XI26/XI8/MM5_g
+ N_VDD_XI26/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI8/MM4 N_XI26/XI8/NET33_XI26/XI8/MM4_d N_XI26/XI8/NET34_XI26/XI8/MM4_g
+ N_VDD_XI26/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI8/MM10 N_XI26/XI8/NET35_XI26/XI8/MM10_d N_XI26/XI8/NET36_XI26/XI8/MM10_g
+ N_VDD_XI26/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI8/MM11 N_XI26/XI8/NET36_XI26/XI8/MM11_d N_XI26/XI8/NET35_XI26/XI8/MM11_g
+ N_VDD_XI26/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI9/MM2 N_XI26/XI9/NET34_XI26/XI9/MM2_d N_XI26/XI9/NET33_XI26/XI9/MM2_g
+ N_VSS_XI26/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM3 N_XI26/XI9/NET33_XI26/XI9/MM3_d N_WL<48>_XI26/XI9/MM3_g
+ N_BLN<6>_XI26/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM0 N_XI26/XI9/NET34_XI26/XI9/MM0_d N_WL<48>_XI26/XI9/MM0_g
+ N_BL<6>_XI26/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM1 N_XI26/XI9/NET33_XI26/XI9/MM1_d N_XI26/XI9/NET34_XI26/XI9/MM1_g
+ N_VSS_XI26/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM9 N_XI26/XI9/NET36_XI26/XI9/MM9_d N_WL<49>_XI26/XI9/MM9_g
+ N_BL<6>_XI26/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM6 N_XI26/XI9/NET35_XI26/XI9/MM6_d N_XI26/XI9/NET36_XI26/XI9/MM6_g
+ N_VSS_XI26/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM7 N_XI26/XI9/NET36_XI26/XI9/MM7_d N_XI26/XI9/NET35_XI26/XI9/MM7_g
+ N_VSS_XI26/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM8 N_XI26/XI9/NET35_XI26/XI9/MM8_d N_WL<49>_XI26/XI9/MM8_g
+ N_BLN<6>_XI26/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI9/MM5 N_XI26/XI9/NET34_XI26/XI9/MM5_d N_XI26/XI9/NET33_XI26/XI9/MM5_g
+ N_VDD_XI26/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI9/MM4 N_XI26/XI9/NET33_XI26/XI9/MM4_d N_XI26/XI9/NET34_XI26/XI9/MM4_g
+ N_VDD_XI26/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI9/MM10 N_XI26/XI9/NET35_XI26/XI9/MM10_d N_XI26/XI9/NET36_XI26/XI9/MM10_g
+ N_VDD_XI26/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI9/MM11 N_XI26/XI9/NET36_XI26/XI9/MM11_d N_XI26/XI9/NET35_XI26/XI9/MM11_g
+ N_VDD_XI26/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI10/MM2 N_XI26/XI10/NET34_XI26/XI10/MM2_d
+ N_XI26/XI10/NET33_XI26/XI10/MM2_g N_VSS_XI26/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI10/MM3 N_XI26/XI10/NET33_XI26/XI10/MM3_d N_WL<48>_XI26/XI10/MM3_g
+ N_BLN<5>_XI26/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI10/MM0 N_XI26/XI10/NET34_XI26/XI10/MM0_d N_WL<48>_XI26/XI10/MM0_g
+ N_BL<5>_XI26/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI10/MM1 N_XI26/XI10/NET33_XI26/XI10/MM1_d
+ N_XI26/XI10/NET34_XI26/XI10/MM1_g N_VSS_XI26/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI10/MM9 N_XI26/XI10/NET36_XI26/XI10/MM9_d N_WL<49>_XI26/XI10/MM9_g
+ N_BL<5>_XI26/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI10/MM6 N_XI26/XI10/NET35_XI26/XI10/MM6_d
+ N_XI26/XI10/NET36_XI26/XI10/MM6_g N_VSS_XI26/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI10/MM7 N_XI26/XI10/NET36_XI26/XI10/MM7_d
+ N_XI26/XI10/NET35_XI26/XI10/MM7_g N_VSS_XI26/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI10/MM8 N_XI26/XI10/NET35_XI26/XI10/MM8_d N_WL<49>_XI26/XI10/MM8_g
+ N_BLN<5>_XI26/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI10/MM5 N_XI26/XI10/NET34_XI26/XI10/MM5_d
+ N_XI26/XI10/NET33_XI26/XI10/MM5_g N_VDD_XI26/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI10/MM4 N_XI26/XI10/NET33_XI26/XI10/MM4_d
+ N_XI26/XI10/NET34_XI26/XI10/MM4_g N_VDD_XI26/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI10/MM10 N_XI26/XI10/NET35_XI26/XI10/MM10_d
+ N_XI26/XI10/NET36_XI26/XI10/MM10_g N_VDD_XI26/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI10/MM11 N_XI26/XI10/NET36_XI26/XI10/MM11_d
+ N_XI26/XI10/NET35_XI26/XI10/MM11_g N_VDD_XI26/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI11/MM2 N_XI26/XI11/NET34_XI26/XI11/MM2_d
+ N_XI26/XI11/NET33_XI26/XI11/MM2_g N_VSS_XI26/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI11/MM3 N_XI26/XI11/NET33_XI26/XI11/MM3_d N_WL<48>_XI26/XI11/MM3_g
+ N_BLN<4>_XI26/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI11/MM0 N_XI26/XI11/NET34_XI26/XI11/MM0_d N_WL<48>_XI26/XI11/MM0_g
+ N_BL<4>_XI26/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI11/MM1 N_XI26/XI11/NET33_XI26/XI11/MM1_d
+ N_XI26/XI11/NET34_XI26/XI11/MM1_g N_VSS_XI26/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI11/MM9 N_XI26/XI11/NET36_XI26/XI11/MM9_d N_WL<49>_XI26/XI11/MM9_g
+ N_BL<4>_XI26/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI11/MM6 N_XI26/XI11/NET35_XI26/XI11/MM6_d
+ N_XI26/XI11/NET36_XI26/XI11/MM6_g N_VSS_XI26/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI11/MM7 N_XI26/XI11/NET36_XI26/XI11/MM7_d
+ N_XI26/XI11/NET35_XI26/XI11/MM7_g N_VSS_XI26/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI11/MM8 N_XI26/XI11/NET35_XI26/XI11/MM8_d N_WL<49>_XI26/XI11/MM8_g
+ N_BLN<4>_XI26/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI11/MM5 N_XI26/XI11/NET34_XI26/XI11/MM5_d
+ N_XI26/XI11/NET33_XI26/XI11/MM5_g N_VDD_XI26/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI11/MM4 N_XI26/XI11/NET33_XI26/XI11/MM4_d
+ N_XI26/XI11/NET34_XI26/XI11/MM4_g N_VDD_XI26/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI11/MM10 N_XI26/XI11/NET35_XI26/XI11/MM10_d
+ N_XI26/XI11/NET36_XI26/XI11/MM10_g N_VDD_XI26/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI11/MM11 N_XI26/XI11/NET36_XI26/XI11/MM11_d
+ N_XI26/XI11/NET35_XI26/XI11/MM11_g N_VDD_XI26/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI12/MM2 N_XI26/XI12/NET34_XI26/XI12/MM2_d
+ N_XI26/XI12/NET33_XI26/XI12/MM2_g N_VSS_XI26/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI12/MM3 N_XI26/XI12/NET33_XI26/XI12/MM3_d N_WL<48>_XI26/XI12/MM3_g
+ N_BLN<3>_XI26/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI12/MM0 N_XI26/XI12/NET34_XI26/XI12/MM0_d N_WL<48>_XI26/XI12/MM0_g
+ N_BL<3>_XI26/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI12/MM1 N_XI26/XI12/NET33_XI26/XI12/MM1_d
+ N_XI26/XI12/NET34_XI26/XI12/MM1_g N_VSS_XI26/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI12/MM9 N_XI26/XI12/NET36_XI26/XI12/MM9_d N_WL<49>_XI26/XI12/MM9_g
+ N_BL<3>_XI26/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI12/MM6 N_XI26/XI12/NET35_XI26/XI12/MM6_d
+ N_XI26/XI12/NET36_XI26/XI12/MM6_g N_VSS_XI26/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI12/MM7 N_XI26/XI12/NET36_XI26/XI12/MM7_d
+ N_XI26/XI12/NET35_XI26/XI12/MM7_g N_VSS_XI26/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI12/MM8 N_XI26/XI12/NET35_XI26/XI12/MM8_d N_WL<49>_XI26/XI12/MM8_g
+ N_BLN<3>_XI26/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI12/MM5 N_XI26/XI12/NET34_XI26/XI12/MM5_d
+ N_XI26/XI12/NET33_XI26/XI12/MM5_g N_VDD_XI26/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI12/MM4 N_XI26/XI12/NET33_XI26/XI12/MM4_d
+ N_XI26/XI12/NET34_XI26/XI12/MM4_g N_VDD_XI26/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI12/MM10 N_XI26/XI12/NET35_XI26/XI12/MM10_d
+ N_XI26/XI12/NET36_XI26/XI12/MM10_g N_VDD_XI26/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI12/MM11 N_XI26/XI12/NET36_XI26/XI12/MM11_d
+ N_XI26/XI12/NET35_XI26/XI12/MM11_g N_VDD_XI26/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI13/MM2 N_XI26/XI13/NET34_XI26/XI13/MM2_d
+ N_XI26/XI13/NET33_XI26/XI13/MM2_g N_VSS_XI26/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI13/MM3 N_XI26/XI13/NET33_XI26/XI13/MM3_d N_WL<48>_XI26/XI13/MM3_g
+ N_BLN<2>_XI26/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI13/MM0 N_XI26/XI13/NET34_XI26/XI13/MM0_d N_WL<48>_XI26/XI13/MM0_g
+ N_BL<2>_XI26/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI13/MM1 N_XI26/XI13/NET33_XI26/XI13/MM1_d
+ N_XI26/XI13/NET34_XI26/XI13/MM1_g N_VSS_XI26/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI13/MM9 N_XI26/XI13/NET36_XI26/XI13/MM9_d N_WL<49>_XI26/XI13/MM9_g
+ N_BL<2>_XI26/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI13/MM6 N_XI26/XI13/NET35_XI26/XI13/MM6_d
+ N_XI26/XI13/NET36_XI26/XI13/MM6_g N_VSS_XI26/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI13/MM7 N_XI26/XI13/NET36_XI26/XI13/MM7_d
+ N_XI26/XI13/NET35_XI26/XI13/MM7_g N_VSS_XI26/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI13/MM8 N_XI26/XI13/NET35_XI26/XI13/MM8_d N_WL<49>_XI26/XI13/MM8_g
+ N_BLN<2>_XI26/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI13/MM5 N_XI26/XI13/NET34_XI26/XI13/MM5_d
+ N_XI26/XI13/NET33_XI26/XI13/MM5_g N_VDD_XI26/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI13/MM4 N_XI26/XI13/NET33_XI26/XI13/MM4_d
+ N_XI26/XI13/NET34_XI26/XI13/MM4_g N_VDD_XI26/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI13/MM10 N_XI26/XI13/NET35_XI26/XI13/MM10_d
+ N_XI26/XI13/NET36_XI26/XI13/MM10_g N_VDD_XI26/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI13/MM11 N_XI26/XI13/NET36_XI26/XI13/MM11_d
+ N_XI26/XI13/NET35_XI26/XI13/MM11_g N_VDD_XI26/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI14/MM2 N_XI26/XI14/NET34_XI26/XI14/MM2_d
+ N_XI26/XI14/NET33_XI26/XI14/MM2_g N_VSS_XI26/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI14/MM3 N_XI26/XI14/NET33_XI26/XI14/MM3_d N_WL<48>_XI26/XI14/MM3_g
+ N_BLN<1>_XI26/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI14/MM0 N_XI26/XI14/NET34_XI26/XI14/MM0_d N_WL<48>_XI26/XI14/MM0_g
+ N_BL<1>_XI26/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI14/MM1 N_XI26/XI14/NET33_XI26/XI14/MM1_d
+ N_XI26/XI14/NET34_XI26/XI14/MM1_g N_VSS_XI26/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI14/MM9 N_XI26/XI14/NET36_XI26/XI14/MM9_d N_WL<49>_XI26/XI14/MM9_g
+ N_BL<1>_XI26/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI14/MM6 N_XI26/XI14/NET35_XI26/XI14/MM6_d
+ N_XI26/XI14/NET36_XI26/XI14/MM6_g N_VSS_XI26/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI14/MM7 N_XI26/XI14/NET36_XI26/XI14/MM7_d
+ N_XI26/XI14/NET35_XI26/XI14/MM7_g N_VSS_XI26/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI14/MM8 N_XI26/XI14/NET35_XI26/XI14/MM8_d N_WL<49>_XI26/XI14/MM8_g
+ N_BLN<1>_XI26/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI14/MM5 N_XI26/XI14/NET34_XI26/XI14/MM5_d
+ N_XI26/XI14/NET33_XI26/XI14/MM5_g N_VDD_XI26/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI14/MM4 N_XI26/XI14/NET33_XI26/XI14/MM4_d
+ N_XI26/XI14/NET34_XI26/XI14/MM4_g N_VDD_XI26/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI14/MM10 N_XI26/XI14/NET35_XI26/XI14/MM10_d
+ N_XI26/XI14/NET36_XI26/XI14/MM10_g N_VDD_XI26/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI14/MM11 N_XI26/XI14/NET36_XI26/XI14/MM11_d
+ N_XI26/XI14/NET35_XI26/XI14/MM11_g N_VDD_XI26/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI15/MM2 N_XI26/XI15/NET34_XI26/XI15/MM2_d
+ N_XI26/XI15/NET33_XI26/XI15/MM2_g N_VSS_XI26/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI15/MM3 N_XI26/XI15/NET33_XI26/XI15/MM3_d N_WL<48>_XI26/XI15/MM3_g
+ N_BLN<0>_XI26/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI15/MM0 N_XI26/XI15/NET34_XI26/XI15/MM0_d N_WL<48>_XI26/XI15/MM0_g
+ N_BL<0>_XI26/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI15/MM1 N_XI26/XI15/NET33_XI26/XI15/MM1_d
+ N_XI26/XI15/NET34_XI26/XI15/MM1_g N_VSS_XI26/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI15/MM9 N_XI26/XI15/NET36_XI26/XI15/MM9_d N_WL<49>_XI26/XI15/MM9_g
+ N_BL<0>_XI26/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI15/MM6 N_XI26/XI15/NET35_XI26/XI15/MM6_d
+ N_XI26/XI15/NET36_XI26/XI15/MM6_g N_VSS_XI26/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI15/MM7 N_XI26/XI15/NET36_XI26/XI15/MM7_d
+ N_XI26/XI15/NET35_XI26/XI15/MM7_g N_VSS_XI26/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI26/XI15/MM8 N_XI26/XI15/NET35_XI26/XI15/MM8_d N_WL<49>_XI26/XI15/MM8_g
+ N_BLN<0>_XI26/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI26/XI15/MM5 N_XI26/XI15/NET34_XI26/XI15/MM5_d
+ N_XI26/XI15/NET33_XI26/XI15/MM5_g N_VDD_XI26/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI15/MM4 N_XI26/XI15/NET33_XI26/XI15/MM4_d
+ N_XI26/XI15/NET34_XI26/XI15/MM4_g N_VDD_XI26/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI15/MM10 N_XI26/XI15/NET35_XI26/XI15/MM10_d
+ N_XI26/XI15/NET36_XI26/XI15/MM10_g N_VDD_XI26/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI26/XI15/MM11 N_XI26/XI15/NET36_XI26/XI15/MM11_d
+ N_XI26/XI15/NET35_XI26/XI15/MM11_g N_VDD_XI26/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI0/MM2 N_XI27/XI0/NET34_XI27/XI0/MM2_d N_XI27/XI0/NET33_XI27/XI0/MM2_g
+ N_VSS_XI27/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI0/MM3 N_XI27/XI0/NET33_XI27/XI0/MM3_d N_WL<50>_XI27/XI0/MM3_g
+ N_BLN<15>_XI27/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI0/MM0 N_XI27/XI0/NET34_XI27/XI0/MM0_d N_WL<50>_XI27/XI0/MM0_g
+ N_BL<15>_XI27/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI0/MM1 N_XI27/XI0/NET33_XI27/XI0/MM1_d N_XI27/XI0/NET34_XI27/XI0/MM1_g
+ N_VSS_XI27/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI0/MM9 N_XI27/XI0/NET36_XI27/XI0/MM9_d N_WL<51>_XI27/XI0/MM9_g
+ N_BL<15>_XI27/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI0/MM6 N_XI27/XI0/NET35_XI27/XI0/MM6_d N_XI27/XI0/NET36_XI27/XI0/MM6_g
+ N_VSS_XI27/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI0/MM7 N_XI27/XI0/NET36_XI27/XI0/MM7_d N_XI27/XI0/NET35_XI27/XI0/MM7_g
+ N_VSS_XI27/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI0/MM8 N_XI27/XI0/NET35_XI27/XI0/MM8_d N_WL<51>_XI27/XI0/MM8_g
+ N_BLN<15>_XI27/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI0/MM5 N_XI27/XI0/NET34_XI27/XI0/MM5_d N_XI27/XI0/NET33_XI27/XI0/MM5_g
+ N_VDD_XI27/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI0/MM4 N_XI27/XI0/NET33_XI27/XI0/MM4_d N_XI27/XI0/NET34_XI27/XI0/MM4_g
+ N_VDD_XI27/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI0/MM10 N_XI27/XI0/NET35_XI27/XI0/MM10_d N_XI27/XI0/NET36_XI27/XI0/MM10_g
+ N_VDD_XI27/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI0/MM11 N_XI27/XI0/NET36_XI27/XI0/MM11_d N_XI27/XI0/NET35_XI27/XI0/MM11_g
+ N_VDD_XI27/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI1/MM2 N_XI27/XI1/NET34_XI27/XI1/MM2_d N_XI27/XI1/NET33_XI27/XI1/MM2_g
+ N_VSS_XI27/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI1/MM3 N_XI27/XI1/NET33_XI27/XI1/MM3_d N_WL<50>_XI27/XI1/MM3_g
+ N_BLN<14>_XI27/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI1/MM0 N_XI27/XI1/NET34_XI27/XI1/MM0_d N_WL<50>_XI27/XI1/MM0_g
+ N_BL<14>_XI27/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI1/MM1 N_XI27/XI1/NET33_XI27/XI1/MM1_d N_XI27/XI1/NET34_XI27/XI1/MM1_g
+ N_VSS_XI27/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI1/MM9 N_XI27/XI1/NET36_XI27/XI1/MM9_d N_WL<51>_XI27/XI1/MM9_g
+ N_BL<14>_XI27/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI1/MM6 N_XI27/XI1/NET35_XI27/XI1/MM6_d N_XI27/XI1/NET36_XI27/XI1/MM6_g
+ N_VSS_XI27/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI1/MM7 N_XI27/XI1/NET36_XI27/XI1/MM7_d N_XI27/XI1/NET35_XI27/XI1/MM7_g
+ N_VSS_XI27/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI1/MM8 N_XI27/XI1/NET35_XI27/XI1/MM8_d N_WL<51>_XI27/XI1/MM8_g
+ N_BLN<14>_XI27/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI1/MM5 N_XI27/XI1/NET34_XI27/XI1/MM5_d N_XI27/XI1/NET33_XI27/XI1/MM5_g
+ N_VDD_XI27/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI1/MM4 N_XI27/XI1/NET33_XI27/XI1/MM4_d N_XI27/XI1/NET34_XI27/XI1/MM4_g
+ N_VDD_XI27/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI1/MM10 N_XI27/XI1/NET35_XI27/XI1/MM10_d N_XI27/XI1/NET36_XI27/XI1/MM10_g
+ N_VDD_XI27/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI1/MM11 N_XI27/XI1/NET36_XI27/XI1/MM11_d N_XI27/XI1/NET35_XI27/XI1/MM11_g
+ N_VDD_XI27/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI2/MM2 N_XI27/XI2/NET34_XI27/XI2/MM2_d N_XI27/XI2/NET33_XI27/XI2/MM2_g
+ N_VSS_XI27/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI2/MM3 N_XI27/XI2/NET33_XI27/XI2/MM3_d N_WL<50>_XI27/XI2/MM3_g
+ N_BLN<13>_XI27/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI2/MM0 N_XI27/XI2/NET34_XI27/XI2/MM0_d N_WL<50>_XI27/XI2/MM0_g
+ N_BL<13>_XI27/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI2/MM1 N_XI27/XI2/NET33_XI27/XI2/MM1_d N_XI27/XI2/NET34_XI27/XI2/MM1_g
+ N_VSS_XI27/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI2/MM9 N_XI27/XI2/NET36_XI27/XI2/MM9_d N_WL<51>_XI27/XI2/MM9_g
+ N_BL<13>_XI27/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI2/MM6 N_XI27/XI2/NET35_XI27/XI2/MM6_d N_XI27/XI2/NET36_XI27/XI2/MM6_g
+ N_VSS_XI27/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI2/MM7 N_XI27/XI2/NET36_XI27/XI2/MM7_d N_XI27/XI2/NET35_XI27/XI2/MM7_g
+ N_VSS_XI27/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI2/MM8 N_XI27/XI2/NET35_XI27/XI2/MM8_d N_WL<51>_XI27/XI2/MM8_g
+ N_BLN<13>_XI27/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI2/MM5 N_XI27/XI2/NET34_XI27/XI2/MM5_d N_XI27/XI2/NET33_XI27/XI2/MM5_g
+ N_VDD_XI27/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI2/MM4 N_XI27/XI2/NET33_XI27/XI2/MM4_d N_XI27/XI2/NET34_XI27/XI2/MM4_g
+ N_VDD_XI27/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI2/MM10 N_XI27/XI2/NET35_XI27/XI2/MM10_d N_XI27/XI2/NET36_XI27/XI2/MM10_g
+ N_VDD_XI27/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI2/MM11 N_XI27/XI2/NET36_XI27/XI2/MM11_d N_XI27/XI2/NET35_XI27/XI2/MM11_g
+ N_VDD_XI27/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI3/MM2 N_XI27/XI3/NET34_XI27/XI3/MM2_d N_XI27/XI3/NET33_XI27/XI3/MM2_g
+ N_VSS_XI27/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI3/MM3 N_XI27/XI3/NET33_XI27/XI3/MM3_d N_WL<50>_XI27/XI3/MM3_g
+ N_BLN<12>_XI27/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI3/MM0 N_XI27/XI3/NET34_XI27/XI3/MM0_d N_WL<50>_XI27/XI3/MM0_g
+ N_BL<12>_XI27/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI3/MM1 N_XI27/XI3/NET33_XI27/XI3/MM1_d N_XI27/XI3/NET34_XI27/XI3/MM1_g
+ N_VSS_XI27/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI3/MM9 N_XI27/XI3/NET36_XI27/XI3/MM9_d N_WL<51>_XI27/XI3/MM9_g
+ N_BL<12>_XI27/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI3/MM6 N_XI27/XI3/NET35_XI27/XI3/MM6_d N_XI27/XI3/NET36_XI27/XI3/MM6_g
+ N_VSS_XI27/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI3/MM7 N_XI27/XI3/NET36_XI27/XI3/MM7_d N_XI27/XI3/NET35_XI27/XI3/MM7_g
+ N_VSS_XI27/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI3/MM8 N_XI27/XI3/NET35_XI27/XI3/MM8_d N_WL<51>_XI27/XI3/MM8_g
+ N_BLN<12>_XI27/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI3/MM5 N_XI27/XI3/NET34_XI27/XI3/MM5_d N_XI27/XI3/NET33_XI27/XI3/MM5_g
+ N_VDD_XI27/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI3/MM4 N_XI27/XI3/NET33_XI27/XI3/MM4_d N_XI27/XI3/NET34_XI27/XI3/MM4_g
+ N_VDD_XI27/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI3/MM10 N_XI27/XI3/NET35_XI27/XI3/MM10_d N_XI27/XI3/NET36_XI27/XI3/MM10_g
+ N_VDD_XI27/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI3/MM11 N_XI27/XI3/NET36_XI27/XI3/MM11_d N_XI27/XI3/NET35_XI27/XI3/MM11_g
+ N_VDD_XI27/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI4/MM2 N_XI27/XI4/NET34_XI27/XI4/MM2_d N_XI27/XI4/NET33_XI27/XI4/MM2_g
+ N_VSS_XI27/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI4/MM3 N_XI27/XI4/NET33_XI27/XI4/MM3_d N_WL<50>_XI27/XI4/MM3_g
+ N_BLN<11>_XI27/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI4/MM0 N_XI27/XI4/NET34_XI27/XI4/MM0_d N_WL<50>_XI27/XI4/MM0_g
+ N_BL<11>_XI27/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI4/MM1 N_XI27/XI4/NET33_XI27/XI4/MM1_d N_XI27/XI4/NET34_XI27/XI4/MM1_g
+ N_VSS_XI27/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI4/MM9 N_XI27/XI4/NET36_XI27/XI4/MM9_d N_WL<51>_XI27/XI4/MM9_g
+ N_BL<11>_XI27/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI4/MM6 N_XI27/XI4/NET35_XI27/XI4/MM6_d N_XI27/XI4/NET36_XI27/XI4/MM6_g
+ N_VSS_XI27/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI4/MM7 N_XI27/XI4/NET36_XI27/XI4/MM7_d N_XI27/XI4/NET35_XI27/XI4/MM7_g
+ N_VSS_XI27/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI4/MM8 N_XI27/XI4/NET35_XI27/XI4/MM8_d N_WL<51>_XI27/XI4/MM8_g
+ N_BLN<11>_XI27/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI4/MM5 N_XI27/XI4/NET34_XI27/XI4/MM5_d N_XI27/XI4/NET33_XI27/XI4/MM5_g
+ N_VDD_XI27/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI4/MM4 N_XI27/XI4/NET33_XI27/XI4/MM4_d N_XI27/XI4/NET34_XI27/XI4/MM4_g
+ N_VDD_XI27/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI4/MM10 N_XI27/XI4/NET35_XI27/XI4/MM10_d N_XI27/XI4/NET36_XI27/XI4/MM10_g
+ N_VDD_XI27/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI4/MM11 N_XI27/XI4/NET36_XI27/XI4/MM11_d N_XI27/XI4/NET35_XI27/XI4/MM11_g
+ N_VDD_XI27/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI5/MM2 N_XI27/XI5/NET34_XI27/XI5/MM2_d N_XI27/XI5/NET33_XI27/XI5/MM2_g
+ N_VSS_XI27/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI5/MM3 N_XI27/XI5/NET33_XI27/XI5/MM3_d N_WL<50>_XI27/XI5/MM3_g
+ N_BLN<10>_XI27/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI5/MM0 N_XI27/XI5/NET34_XI27/XI5/MM0_d N_WL<50>_XI27/XI5/MM0_g
+ N_BL<10>_XI27/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI5/MM1 N_XI27/XI5/NET33_XI27/XI5/MM1_d N_XI27/XI5/NET34_XI27/XI5/MM1_g
+ N_VSS_XI27/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI5/MM9 N_XI27/XI5/NET36_XI27/XI5/MM9_d N_WL<51>_XI27/XI5/MM9_g
+ N_BL<10>_XI27/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI5/MM6 N_XI27/XI5/NET35_XI27/XI5/MM6_d N_XI27/XI5/NET36_XI27/XI5/MM6_g
+ N_VSS_XI27/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI5/MM7 N_XI27/XI5/NET36_XI27/XI5/MM7_d N_XI27/XI5/NET35_XI27/XI5/MM7_g
+ N_VSS_XI27/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI5/MM8 N_XI27/XI5/NET35_XI27/XI5/MM8_d N_WL<51>_XI27/XI5/MM8_g
+ N_BLN<10>_XI27/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI5/MM5 N_XI27/XI5/NET34_XI27/XI5/MM5_d N_XI27/XI5/NET33_XI27/XI5/MM5_g
+ N_VDD_XI27/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI5/MM4 N_XI27/XI5/NET33_XI27/XI5/MM4_d N_XI27/XI5/NET34_XI27/XI5/MM4_g
+ N_VDD_XI27/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI5/MM10 N_XI27/XI5/NET35_XI27/XI5/MM10_d N_XI27/XI5/NET36_XI27/XI5/MM10_g
+ N_VDD_XI27/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI5/MM11 N_XI27/XI5/NET36_XI27/XI5/MM11_d N_XI27/XI5/NET35_XI27/XI5/MM11_g
+ N_VDD_XI27/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI6/MM2 N_XI27/XI6/NET34_XI27/XI6/MM2_d N_XI27/XI6/NET33_XI27/XI6/MM2_g
+ N_VSS_XI27/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM3 N_XI27/XI6/NET33_XI27/XI6/MM3_d N_WL<50>_XI27/XI6/MM3_g
+ N_BLN<9>_XI27/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM0 N_XI27/XI6/NET34_XI27/XI6/MM0_d N_WL<50>_XI27/XI6/MM0_g
+ N_BL<9>_XI27/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM1 N_XI27/XI6/NET33_XI27/XI6/MM1_d N_XI27/XI6/NET34_XI27/XI6/MM1_g
+ N_VSS_XI27/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM9 N_XI27/XI6/NET36_XI27/XI6/MM9_d N_WL<51>_XI27/XI6/MM9_g
+ N_BL<9>_XI27/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM6 N_XI27/XI6/NET35_XI27/XI6/MM6_d N_XI27/XI6/NET36_XI27/XI6/MM6_g
+ N_VSS_XI27/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM7 N_XI27/XI6/NET36_XI27/XI6/MM7_d N_XI27/XI6/NET35_XI27/XI6/MM7_g
+ N_VSS_XI27/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM8 N_XI27/XI6/NET35_XI27/XI6/MM8_d N_WL<51>_XI27/XI6/MM8_g
+ N_BLN<9>_XI27/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI6/MM5 N_XI27/XI6/NET34_XI27/XI6/MM5_d N_XI27/XI6/NET33_XI27/XI6/MM5_g
+ N_VDD_XI27/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI6/MM4 N_XI27/XI6/NET33_XI27/XI6/MM4_d N_XI27/XI6/NET34_XI27/XI6/MM4_g
+ N_VDD_XI27/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI6/MM10 N_XI27/XI6/NET35_XI27/XI6/MM10_d N_XI27/XI6/NET36_XI27/XI6/MM10_g
+ N_VDD_XI27/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI6/MM11 N_XI27/XI6/NET36_XI27/XI6/MM11_d N_XI27/XI6/NET35_XI27/XI6/MM11_g
+ N_VDD_XI27/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI7/MM2 N_XI27/XI7/NET34_XI27/XI7/MM2_d N_XI27/XI7/NET33_XI27/XI7/MM2_g
+ N_VSS_XI27/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM3 N_XI27/XI7/NET33_XI27/XI7/MM3_d N_WL<50>_XI27/XI7/MM3_g
+ N_BLN<8>_XI27/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM0 N_XI27/XI7/NET34_XI27/XI7/MM0_d N_WL<50>_XI27/XI7/MM0_g
+ N_BL<8>_XI27/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM1 N_XI27/XI7/NET33_XI27/XI7/MM1_d N_XI27/XI7/NET34_XI27/XI7/MM1_g
+ N_VSS_XI27/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM9 N_XI27/XI7/NET36_XI27/XI7/MM9_d N_WL<51>_XI27/XI7/MM9_g
+ N_BL<8>_XI27/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM6 N_XI27/XI7/NET35_XI27/XI7/MM6_d N_XI27/XI7/NET36_XI27/XI7/MM6_g
+ N_VSS_XI27/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM7 N_XI27/XI7/NET36_XI27/XI7/MM7_d N_XI27/XI7/NET35_XI27/XI7/MM7_g
+ N_VSS_XI27/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM8 N_XI27/XI7/NET35_XI27/XI7/MM8_d N_WL<51>_XI27/XI7/MM8_g
+ N_BLN<8>_XI27/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI7/MM5 N_XI27/XI7/NET34_XI27/XI7/MM5_d N_XI27/XI7/NET33_XI27/XI7/MM5_g
+ N_VDD_XI27/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI7/MM4 N_XI27/XI7/NET33_XI27/XI7/MM4_d N_XI27/XI7/NET34_XI27/XI7/MM4_g
+ N_VDD_XI27/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI7/MM10 N_XI27/XI7/NET35_XI27/XI7/MM10_d N_XI27/XI7/NET36_XI27/XI7/MM10_g
+ N_VDD_XI27/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI7/MM11 N_XI27/XI7/NET36_XI27/XI7/MM11_d N_XI27/XI7/NET35_XI27/XI7/MM11_g
+ N_VDD_XI27/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI8/MM2 N_XI27/XI8/NET34_XI27/XI8/MM2_d N_XI27/XI8/NET33_XI27/XI8/MM2_g
+ N_VSS_XI27/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM3 N_XI27/XI8/NET33_XI27/XI8/MM3_d N_WL<50>_XI27/XI8/MM3_g
+ N_BLN<7>_XI27/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM0 N_XI27/XI8/NET34_XI27/XI8/MM0_d N_WL<50>_XI27/XI8/MM0_g
+ N_BL<7>_XI27/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM1 N_XI27/XI8/NET33_XI27/XI8/MM1_d N_XI27/XI8/NET34_XI27/XI8/MM1_g
+ N_VSS_XI27/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM9 N_XI27/XI8/NET36_XI27/XI8/MM9_d N_WL<51>_XI27/XI8/MM9_g
+ N_BL<7>_XI27/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM6 N_XI27/XI8/NET35_XI27/XI8/MM6_d N_XI27/XI8/NET36_XI27/XI8/MM6_g
+ N_VSS_XI27/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM7 N_XI27/XI8/NET36_XI27/XI8/MM7_d N_XI27/XI8/NET35_XI27/XI8/MM7_g
+ N_VSS_XI27/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM8 N_XI27/XI8/NET35_XI27/XI8/MM8_d N_WL<51>_XI27/XI8/MM8_g
+ N_BLN<7>_XI27/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI8/MM5 N_XI27/XI8/NET34_XI27/XI8/MM5_d N_XI27/XI8/NET33_XI27/XI8/MM5_g
+ N_VDD_XI27/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI8/MM4 N_XI27/XI8/NET33_XI27/XI8/MM4_d N_XI27/XI8/NET34_XI27/XI8/MM4_g
+ N_VDD_XI27/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI8/MM10 N_XI27/XI8/NET35_XI27/XI8/MM10_d N_XI27/XI8/NET36_XI27/XI8/MM10_g
+ N_VDD_XI27/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI8/MM11 N_XI27/XI8/NET36_XI27/XI8/MM11_d N_XI27/XI8/NET35_XI27/XI8/MM11_g
+ N_VDD_XI27/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI9/MM2 N_XI27/XI9/NET34_XI27/XI9/MM2_d N_XI27/XI9/NET33_XI27/XI9/MM2_g
+ N_VSS_XI27/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM3 N_XI27/XI9/NET33_XI27/XI9/MM3_d N_WL<50>_XI27/XI9/MM3_g
+ N_BLN<6>_XI27/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM0 N_XI27/XI9/NET34_XI27/XI9/MM0_d N_WL<50>_XI27/XI9/MM0_g
+ N_BL<6>_XI27/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM1 N_XI27/XI9/NET33_XI27/XI9/MM1_d N_XI27/XI9/NET34_XI27/XI9/MM1_g
+ N_VSS_XI27/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM9 N_XI27/XI9/NET36_XI27/XI9/MM9_d N_WL<51>_XI27/XI9/MM9_g
+ N_BL<6>_XI27/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM6 N_XI27/XI9/NET35_XI27/XI9/MM6_d N_XI27/XI9/NET36_XI27/XI9/MM6_g
+ N_VSS_XI27/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM7 N_XI27/XI9/NET36_XI27/XI9/MM7_d N_XI27/XI9/NET35_XI27/XI9/MM7_g
+ N_VSS_XI27/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM8 N_XI27/XI9/NET35_XI27/XI9/MM8_d N_WL<51>_XI27/XI9/MM8_g
+ N_BLN<6>_XI27/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI9/MM5 N_XI27/XI9/NET34_XI27/XI9/MM5_d N_XI27/XI9/NET33_XI27/XI9/MM5_g
+ N_VDD_XI27/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI9/MM4 N_XI27/XI9/NET33_XI27/XI9/MM4_d N_XI27/XI9/NET34_XI27/XI9/MM4_g
+ N_VDD_XI27/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI9/MM10 N_XI27/XI9/NET35_XI27/XI9/MM10_d N_XI27/XI9/NET36_XI27/XI9/MM10_g
+ N_VDD_XI27/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI9/MM11 N_XI27/XI9/NET36_XI27/XI9/MM11_d N_XI27/XI9/NET35_XI27/XI9/MM11_g
+ N_VDD_XI27/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI10/MM2 N_XI27/XI10/NET34_XI27/XI10/MM2_d
+ N_XI27/XI10/NET33_XI27/XI10/MM2_g N_VSS_XI27/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI10/MM3 N_XI27/XI10/NET33_XI27/XI10/MM3_d N_WL<50>_XI27/XI10/MM3_g
+ N_BLN<5>_XI27/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI10/MM0 N_XI27/XI10/NET34_XI27/XI10/MM0_d N_WL<50>_XI27/XI10/MM0_g
+ N_BL<5>_XI27/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI10/MM1 N_XI27/XI10/NET33_XI27/XI10/MM1_d
+ N_XI27/XI10/NET34_XI27/XI10/MM1_g N_VSS_XI27/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI10/MM9 N_XI27/XI10/NET36_XI27/XI10/MM9_d N_WL<51>_XI27/XI10/MM9_g
+ N_BL<5>_XI27/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI10/MM6 N_XI27/XI10/NET35_XI27/XI10/MM6_d
+ N_XI27/XI10/NET36_XI27/XI10/MM6_g N_VSS_XI27/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI10/MM7 N_XI27/XI10/NET36_XI27/XI10/MM7_d
+ N_XI27/XI10/NET35_XI27/XI10/MM7_g N_VSS_XI27/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI10/MM8 N_XI27/XI10/NET35_XI27/XI10/MM8_d N_WL<51>_XI27/XI10/MM8_g
+ N_BLN<5>_XI27/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI10/MM5 N_XI27/XI10/NET34_XI27/XI10/MM5_d
+ N_XI27/XI10/NET33_XI27/XI10/MM5_g N_VDD_XI27/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI10/MM4 N_XI27/XI10/NET33_XI27/XI10/MM4_d
+ N_XI27/XI10/NET34_XI27/XI10/MM4_g N_VDD_XI27/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI10/MM10 N_XI27/XI10/NET35_XI27/XI10/MM10_d
+ N_XI27/XI10/NET36_XI27/XI10/MM10_g N_VDD_XI27/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI10/MM11 N_XI27/XI10/NET36_XI27/XI10/MM11_d
+ N_XI27/XI10/NET35_XI27/XI10/MM11_g N_VDD_XI27/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI11/MM2 N_XI27/XI11/NET34_XI27/XI11/MM2_d
+ N_XI27/XI11/NET33_XI27/XI11/MM2_g N_VSS_XI27/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI11/MM3 N_XI27/XI11/NET33_XI27/XI11/MM3_d N_WL<50>_XI27/XI11/MM3_g
+ N_BLN<4>_XI27/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI11/MM0 N_XI27/XI11/NET34_XI27/XI11/MM0_d N_WL<50>_XI27/XI11/MM0_g
+ N_BL<4>_XI27/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI11/MM1 N_XI27/XI11/NET33_XI27/XI11/MM1_d
+ N_XI27/XI11/NET34_XI27/XI11/MM1_g N_VSS_XI27/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI11/MM9 N_XI27/XI11/NET36_XI27/XI11/MM9_d N_WL<51>_XI27/XI11/MM9_g
+ N_BL<4>_XI27/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI11/MM6 N_XI27/XI11/NET35_XI27/XI11/MM6_d
+ N_XI27/XI11/NET36_XI27/XI11/MM6_g N_VSS_XI27/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI11/MM7 N_XI27/XI11/NET36_XI27/XI11/MM7_d
+ N_XI27/XI11/NET35_XI27/XI11/MM7_g N_VSS_XI27/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI11/MM8 N_XI27/XI11/NET35_XI27/XI11/MM8_d N_WL<51>_XI27/XI11/MM8_g
+ N_BLN<4>_XI27/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI11/MM5 N_XI27/XI11/NET34_XI27/XI11/MM5_d
+ N_XI27/XI11/NET33_XI27/XI11/MM5_g N_VDD_XI27/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI11/MM4 N_XI27/XI11/NET33_XI27/XI11/MM4_d
+ N_XI27/XI11/NET34_XI27/XI11/MM4_g N_VDD_XI27/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI11/MM10 N_XI27/XI11/NET35_XI27/XI11/MM10_d
+ N_XI27/XI11/NET36_XI27/XI11/MM10_g N_VDD_XI27/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI11/MM11 N_XI27/XI11/NET36_XI27/XI11/MM11_d
+ N_XI27/XI11/NET35_XI27/XI11/MM11_g N_VDD_XI27/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI12/MM2 N_XI27/XI12/NET34_XI27/XI12/MM2_d
+ N_XI27/XI12/NET33_XI27/XI12/MM2_g N_VSS_XI27/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI12/MM3 N_XI27/XI12/NET33_XI27/XI12/MM3_d N_WL<50>_XI27/XI12/MM3_g
+ N_BLN<3>_XI27/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI12/MM0 N_XI27/XI12/NET34_XI27/XI12/MM0_d N_WL<50>_XI27/XI12/MM0_g
+ N_BL<3>_XI27/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI12/MM1 N_XI27/XI12/NET33_XI27/XI12/MM1_d
+ N_XI27/XI12/NET34_XI27/XI12/MM1_g N_VSS_XI27/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI12/MM9 N_XI27/XI12/NET36_XI27/XI12/MM9_d N_WL<51>_XI27/XI12/MM9_g
+ N_BL<3>_XI27/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI12/MM6 N_XI27/XI12/NET35_XI27/XI12/MM6_d
+ N_XI27/XI12/NET36_XI27/XI12/MM6_g N_VSS_XI27/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI12/MM7 N_XI27/XI12/NET36_XI27/XI12/MM7_d
+ N_XI27/XI12/NET35_XI27/XI12/MM7_g N_VSS_XI27/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI12/MM8 N_XI27/XI12/NET35_XI27/XI12/MM8_d N_WL<51>_XI27/XI12/MM8_g
+ N_BLN<3>_XI27/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI12/MM5 N_XI27/XI12/NET34_XI27/XI12/MM5_d
+ N_XI27/XI12/NET33_XI27/XI12/MM5_g N_VDD_XI27/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI12/MM4 N_XI27/XI12/NET33_XI27/XI12/MM4_d
+ N_XI27/XI12/NET34_XI27/XI12/MM4_g N_VDD_XI27/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI12/MM10 N_XI27/XI12/NET35_XI27/XI12/MM10_d
+ N_XI27/XI12/NET36_XI27/XI12/MM10_g N_VDD_XI27/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI12/MM11 N_XI27/XI12/NET36_XI27/XI12/MM11_d
+ N_XI27/XI12/NET35_XI27/XI12/MM11_g N_VDD_XI27/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI13/MM2 N_XI27/XI13/NET34_XI27/XI13/MM2_d
+ N_XI27/XI13/NET33_XI27/XI13/MM2_g N_VSS_XI27/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI13/MM3 N_XI27/XI13/NET33_XI27/XI13/MM3_d N_WL<50>_XI27/XI13/MM3_g
+ N_BLN<2>_XI27/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI13/MM0 N_XI27/XI13/NET34_XI27/XI13/MM0_d N_WL<50>_XI27/XI13/MM0_g
+ N_BL<2>_XI27/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI13/MM1 N_XI27/XI13/NET33_XI27/XI13/MM1_d
+ N_XI27/XI13/NET34_XI27/XI13/MM1_g N_VSS_XI27/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI13/MM9 N_XI27/XI13/NET36_XI27/XI13/MM9_d N_WL<51>_XI27/XI13/MM9_g
+ N_BL<2>_XI27/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI13/MM6 N_XI27/XI13/NET35_XI27/XI13/MM6_d
+ N_XI27/XI13/NET36_XI27/XI13/MM6_g N_VSS_XI27/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI13/MM7 N_XI27/XI13/NET36_XI27/XI13/MM7_d
+ N_XI27/XI13/NET35_XI27/XI13/MM7_g N_VSS_XI27/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI13/MM8 N_XI27/XI13/NET35_XI27/XI13/MM8_d N_WL<51>_XI27/XI13/MM8_g
+ N_BLN<2>_XI27/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI13/MM5 N_XI27/XI13/NET34_XI27/XI13/MM5_d
+ N_XI27/XI13/NET33_XI27/XI13/MM5_g N_VDD_XI27/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI13/MM4 N_XI27/XI13/NET33_XI27/XI13/MM4_d
+ N_XI27/XI13/NET34_XI27/XI13/MM4_g N_VDD_XI27/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI13/MM10 N_XI27/XI13/NET35_XI27/XI13/MM10_d
+ N_XI27/XI13/NET36_XI27/XI13/MM10_g N_VDD_XI27/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI13/MM11 N_XI27/XI13/NET36_XI27/XI13/MM11_d
+ N_XI27/XI13/NET35_XI27/XI13/MM11_g N_VDD_XI27/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI14/MM2 N_XI27/XI14/NET34_XI27/XI14/MM2_d
+ N_XI27/XI14/NET33_XI27/XI14/MM2_g N_VSS_XI27/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI14/MM3 N_XI27/XI14/NET33_XI27/XI14/MM3_d N_WL<50>_XI27/XI14/MM3_g
+ N_BLN<1>_XI27/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI14/MM0 N_XI27/XI14/NET34_XI27/XI14/MM0_d N_WL<50>_XI27/XI14/MM0_g
+ N_BL<1>_XI27/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI14/MM1 N_XI27/XI14/NET33_XI27/XI14/MM1_d
+ N_XI27/XI14/NET34_XI27/XI14/MM1_g N_VSS_XI27/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI14/MM9 N_XI27/XI14/NET36_XI27/XI14/MM9_d N_WL<51>_XI27/XI14/MM9_g
+ N_BL<1>_XI27/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI14/MM6 N_XI27/XI14/NET35_XI27/XI14/MM6_d
+ N_XI27/XI14/NET36_XI27/XI14/MM6_g N_VSS_XI27/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI14/MM7 N_XI27/XI14/NET36_XI27/XI14/MM7_d
+ N_XI27/XI14/NET35_XI27/XI14/MM7_g N_VSS_XI27/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI14/MM8 N_XI27/XI14/NET35_XI27/XI14/MM8_d N_WL<51>_XI27/XI14/MM8_g
+ N_BLN<1>_XI27/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI14/MM5 N_XI27/XI14/NET34_XI27/XI14/MM5_d
+ N_XI27/XI14/NET33_XI27/XI14/MM5_g N_VDD_XI27/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI14/MM4 N_XI27/XI14/NET33_XI27/XI14/MM4_d
+ N_XI27/XI14/NET34_XI27/XI14/MM4_g N_VDD_XI27/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI14/MM10 N_XI27/XI14/NET35_XI27/XI14/MM10_d
+ N_XI27/XI14/NET36_XI27/XI14/MM10_g N_VDD_XI27/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI14/MM11 N_XI27/XI14/NET36_XI27/XI14/MM11_d
+ N_XI27/XI14/NET35_XI27/XI14/MM11_g N_VDD_XI27/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI15/MM2 N_XI27/XI15/NET34_XI27/XI15/MM2_d
+ N_XI27/XI15/NET33_XI27/XI15/MM2_g N_VSS_XI27/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI15/MM3 N_XI27/XI15/NET33_XI27/XI15/MM3_d N_WL<50>_XI27/XI15/MM3_g
+ N_BLN<0>_XI27/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI15/MM0 N_XI27/XI15/NET34_XI27/XI15/MM0_d N_WL<50>_XI27/XI15/MM0_g
+ N_BL<0>_XI27/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI15/MM1 N_XI27/XI15/NET33_XI27/XI15/MM1_d
+ N_XI27/XI15/NET34_XI27/XI15/MM1_g N_VSS_XI27/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI15/MM9 N_XI27/XI15/NET36_XI27/XI15/MM9_d N_WL<51>_XI27/XI15/MM9_g
+ N_BL<0>_XI27/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI15/MM6 N_XI27/XI15/NET35_XI27/XI15/MM6_d
+ N_XI27/XI15/NET36_XI27/XI15/MM6_g N_VSS_XI27/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI15/MM7 N_XI27/XI15/NET36_XI27/XI15/MM7_d
+ N_XI27/XI15/NET35_XI27/XI15/MM7_g N_VSS_XI27/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI27/XI15/MM8 N_XI27/XI15/NET35_XI27/XI15/MM8_d N_WL<51>_XI27/XI15/MM8_g
+ N_BLN<0>_XI27/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI27/XI15/MM5 N_XI27/XI15/NET34_XI27/XI15/MM5_d
+ N_XI27/XI15/NET33_XI27/XI15/MM5_g N_VDD_XI27/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI15/MM4 N_XI27/XI15/NET33_XI27/XI15/MM4_d
+ N_XI27/XI15/NET34_XI27/XI15/MM4_g N_VDD_XI27/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI15/MM10 N_XI27/XI15/NET35_XI27/XI15/MM10_d
+ N_XI27/XI15/NET36_XI27/XI15/MM10_g N_VDD_XI27/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI27/XI15/MM11 N_XI27/XI15/NET36_XI27/XI15/MM11_d
+ N_XI27/XI15/NET35_XI27/XI15/MM11_g N_VDD_XI27/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI0/MM2 N_XI28/XI0/NET34_XI28/XI0/MM2_d N_XI28/XI0/NET33_XI28/XI0/MM2_g
+ N_VSS_XI28/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI0/MM3 N_XI28/XI0/NET33_XI28/XI0/MM3_d N_WL<52>_XI28/XI0/MM3_g
+ N_BLN<15>_XI28/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI0/MM0 N_XI28/XI0/NET34_XI28/XI0/MM0_d N_WL<52>_XI28/XI0/MM0_g
+ N_BL<15>_XI28/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI0/MM1 N_XI28/XI0/NET33_XI28/XI0/MM1_d N_XI28/XI0/NET34_XI28/XI0/MM1_g
+ N_VSS_XI28/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI0/MM9 N_XI28/XI0/NET36_XI28/XI0/MM9_d N_WL<53>_XI28/XI0/MM9_g
+ N_BL<15>_XI28/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI0/MM6 N_XI28/XI0/NET35_XI28/XI0/MM6_d N_XI28/XI0/NET36_XI28/XI0/MM6_g
+ N_VSS_XI28/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI0/MM7 N_XI28/XI0/NET36_XI28/XI0/MM7_d N_XI28/XI0/NET35_XI28/XI0/MM7_g
+ N_VSS_XI28/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI0/MM8 N_XI28/XI0/NET35_XI28/XI0/MM8_d N_WL<53>_XI28/XI0/MM8_g
+ N_BLN<15>_XI28/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI0/MM5 N_XI28/XI0/NET34_XI28/XI0/MM5_d N_XI28/XI0/NET33_XI28/XI0/MM5_g
+ N_VDD_XI28/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI0/MM4 N_XI28/XI0/NET33_XI28/XI0/MM4_d N_XI28/XI0/NET34_XI28/XI0/MM4_g
+ N_VDD_XI28/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI0/MM10 N_XI28/XI0/NET35_XI28/XI0/MM10_d N_XI28/XI0/NET36_XI28/XI0/MM10_g
+ N_VDD_XI28/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI0/MM11 N_XI28/XI0/NET36_XI28/XI0/MM11_d N_XI28/XI0/NET35_XI28/XI0/MM11_g
+ N_VDD_XI28/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI1/MM2 N_XI28/XI1/NET34_XI28/XI1/MM2_d N_XI28/XI1/NET33_XI28/XI1/MM2_g
+ N_VSS_XI28/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI1/MM3 N_XI28/XI1/NET33_XI28/XI1/MM3_d N_WL<52>_XI28/XI1/MM3_g
+ N_BLN<14>_XI28/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI1/MM0 N_XI28/XI1/NET34_XI28/XI1/MM0_d N_WL<52>_XI28/XI1/MM0_g
+ N_BL<14>_XI28/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI1/MM1 N_XI28/XI1/NET33_XI28/XI1/MM1_d N_XI28/XI1/NET34_XI28/XI1/MM1_g
+ N_VSS_XI28/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI1/MM9 N_XI28/XI1/NET36_XI28/XI1/MM9_d N_WL<53>_XI28/XI1/MM9_g
+ N_BL<14>_XI28/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI1/MM6 N_XI28/XI1/NET35_XI28/XI1/MM6_d N_XI28/XI1/NET36_XI28/XI1/MM6_g
+ N_VSS_XI28/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI1/MM7 N_XI28/XI1/NET36_XI28/XI1/MM7_d N_XI28/XI1/NET35_XI28/XI1/MM7_g
+ N_VSS_XI28/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI1/MM8 N_XI28/XI1/NET35_XI28/XI1/MM8_d N_WL<53>_XI28/XI1/MM8_g
+ N_BLN<14>_XI28/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI1/MM5 N_XI28/XI1/NET34_XI28/XI1/MM5_d N_XI28/XI1/NET33_XI28/XI1/MM5_g
+ N_VDD_XI28/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI1/MM4 N_XI28/XI1/NET33_XI28/XI1/MM4_d N_XI28/XI1/NET34_XI28/XI1/MM4_g
+ N_VDD_XI28/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI1/MM10 N_XI28/XI1/NET35_XI28/XI1/MM10_d N_XI28/XI1/NET36_XI28/XI1/MM10_g
+ N_VDD_XI28/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI1/MM11 N_XI28/XI1/NET36_XI28/XI1/MM11_d N_XI28/XI1/NET35_XI28/XI1/MM11_g
+ N_VDD_XI28/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI2/MM2 N_XI28/XI2/NET34_XI28/XI2/MM2_d N_XI28/XI2/NET33_XI28/XI2/MM2_g
+ N_VSS_XI28/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI2/MM3 N_XI28/XI2/NET33_XI28/XI2/MM3_d N_WL<52>_XI28/XI2/MM3_g
+ N_BLN<13>_XI28/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI2/MM0 N_XI28/XI2/NET34_XI28/XI2/MM0_d N_WL<52>_XI28/XI2/MM0_g
+ N_BL<13>_XI28/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI2/MM1 N_XI28/XI2/NET33_XI28/XI2/MM1_d N_XI28/XI2/NET34_XI28/XI2/MM1_g
+ N_VSS_XI28/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI2/MM9 N_XI28/XI2/NET36_XI28/XI2/MM9_d N_WL<53>_XI28/XI2/MM9_g
+ N_BL<13>_XI28/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI2/MM6 N_XI28/XI2/NET35_XI28/XI2/MM6_d N_XI28/XI2/NET36_XI28/XI2/MM6_g
+ N_VSS_XI28/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI2/MM7 N_XI28/XI2/NET36_XI28/XI2/MM7_d N_XI28/XI2/NET35_XI28/XI2/MM7_g
+ N_VSS_XI28/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI2/MM8 N_XI28/XI2/NET35_XI28/XI2/MM8_d N_WL<53>_XI28/XI2/MM8_g
+ N_BLN<13>_XI28/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI2/MM5 N_XI28/XI2/NET34_XI28/XI2/MM5_d N_XI28/XI2/NET33_XI28/XI2/MM5_g
+ N_VDD_XI28/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI2/MM4 N_XI28/XI2/NET33_XI28/XI2/MM4_d N_XI28/XI2/NET34_XI28/XI2/MM4_g
+ N_VDD_XI28/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI2/MM10 N_XI28/XI2/NET35_XI28/XI2/MM10_d N_XI28/XI2/NET36_XI28/XI2/MM10_g
+ N_VDD_XI28/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI2/MM11 N_XI28/XI2/NET36_XI28/XI2/MM11_d N_XI28/XI2/NET35_XI28/XI2/MM11_g
+ N_VDD_XI28/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI3/MM2 N_XI28/XI3/NET34_XI28/XI3/MM2_d N_XI28/XI3/NET33_XI28/XI3/MM2_g
+ N_VSS_XI28/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI3/MM3 N_XI28/XI3/NET33_XI28/XI3/MM3_d N_WL<52>_XI28/XI3/MM3_g
+ N_BLN<12>_XI28/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI3/MM0 N_XI28/XI3/NET34_XI28/XI3/MM0_d N_WL<52>_XI28/XI3/MM0_g
+ N_BL<12>_XI28/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI3/MM1 N_XI28/XI3/NET33_XI28/XI3/MM1_d N_XI28/XI3/NET34_XI28/XI3/MM1_g
+ N_VSS_XI28/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI3/MM9 N_XI28/XI3/NET36_XI28/XI3/MM9_d N_WL<53>_XI28/XI3/MM9_g
+ N_BL<12>_XI28/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI3/MM6 N_XI28/XI3/NET35_XI28/XI3/MM6_d N_XI28/XI3/NET36_XI28/XI3/MM6_g
+ N_VSS_XI28/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI3/MM7 N_XI28/XI3/NET36_XI28/XI3/MM7_d N_XI28/XI3/NET35_XI28/XI3/MM7_g
+ N_VSS_XI28/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI3/MM8 N_XI28/XI3/NET35_XI28/XI3/MM8_d N_WL<53>_XI28/XI3/MM8_g
+ N_BLN<12>_XI28/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI3/MM5 N_XI28/XI3/NET34_XI28/XI3/MM5_d N_XI28/XI3/NET33_XI28/XI3/MM5_g
+ N_VDD_XI28/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI3/MM4 N_XI28/XI3/NET33_XI28/XI3/MM4_d N_XI28/XI3/NET34_XI28/XI3/MM4_g
+ N_VDD_XI28/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI3/MM10 N_XI28/XI3/NET35_XI28/XI3/MM10_d N_XI28/XI3/NET36_XI28/XI3/MM10_g
+ N_VDD_XI28/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI3/MM11 N_XI28/XI3/NET36_XI28/XI3/MM11_d N_XI28/XI3/NET35_XI28/XI3/MM11_g
+ N_VDD_XI28/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI4/MM2 N_XI28/XI4/NET34_XI28/XI4/MM2_d N_XI28/XI4/NET33_XI28/XI4/MM2_g
+ N_VSS_XI28/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI4/MM3 N_XI28/XI4/NET33_XI28/XI4/MM3_d N_WL<52>_XI28/XI4/MM3_g
+ N_BLN<11>_XI28/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI4/MM0 N_XI28/XI4/NET34_XI28/XI4/MM0_d N_WL<52>_XI28/XI4/MM0_g
+ N_BL<11>_XI28/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI4/MM1 N_XI28/XI4/NET33_XI28/XI4/MM1_d N_XI28/XI4/NET34_XI28/XI4/MM1_g
+ N_VSS_XI28/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI4/MM9 N_XI28/XI4/NET36_XI28/XI4/MM9_d N_WL<53>_XI28/XI4/MM9_g
+ N_BL<11>_XI28/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI4/MM6 N_XI28/XI4/NET35_XI28/XI4/MM6_d N_XI28/XI4/NET36_XI28/XI4/MM6_g
+ N_VSS_XI28/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI4/MM7 N_XI28/XI4/NET36_XI28/XI4/MM7_d N_XI28/XI4/NET35_XI28/XI4/MM7_g
+ N_VSS_XI28/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI4/MM8 N_XI28/XI4/NET35_XI28/XI4/MM8_d N_WL<53>_XI28/XI4/MM8_g
+ N_BLN<11>_XI28/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI4/MM5 N_XI28/XI4/NET34_XI28/XI4/MM5_d N_XI28/XI4/NET33_XI28/XI4/MM5_g
+ N_VDD_XI28/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI4/MM4 N_XI28/XI4/NET33_XI28/XI4/MM4_d N_XI28/XI4/NET34_XI28/XI4/MM4_g
+ N_VDD_XI28/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI4/MM10 N_XI28/XI4/NET35_XI28/XI4/MM10_d N_XI28/XI4/NET36_XI28/XI4/MM10_g
+ N_VDD_XI28/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI4/MM11 N_XI28/XI4/NET36_XI28/XI4/MM11_d N_XI28/XI4/NET35_XI28/XI4/MM11_g
+ N_VDD_XI28/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI5/MM2 N_XI28/XI5/NET34_XI28/XI5/MM2_d N_XI28/XI5/NET33_XI28/XI5/MM2_g
+ N_VSS_XI28/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI5/MM3 N_XI28/XI5/NET33_XI28/XI5/MM3_d N_WL<52>_XI28/XI5/MM3_g
+ N_BLN<10>_XI28/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI5/MM0 N_XI28/XI5/NET34_XI28/XI5/MM0_d N_WL<52>_XI28/XI5/MM0_g
+ N_BL<10>_XI28/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI5/MM1 N_XI28/XI5/NET33_XI28/XI5/MM1_d N_XI28/XI5/NET34_XI28/XI5/MM1_g
+ N_VSS_XI28/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI5/MM9 N_XI28/XI5/NET36_XI28/XI5/MM9_d N_WL<53>_XI28/XI5/MM9_g
+ N_BL<10>_XI28/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI5/MM6 N_XI28/XI5/NET35_XI28/XI5/MM6_d N_XI28/XI5/NET36_XI28/XI5/MM6_g
+ N_VSS_XI28/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI5/MM7 N_XI28/XI5/NET36_XI28/XI5/MM7_d N_XI28/XI5/NET35_XI28/XI5/MM7_g
+ N_VSS_XI28/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI5/MM8 N_XI28/XI5/NET35_XI28/XI5/MM8_d N_WL<53>_XI28/XI5/MM8_g
+ N_BLN<10>_XI28/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI5/MM5 N_XI28/XI5/NET34_XI28/XI5/MM5_d N_XI28/XI5/NET33_XI28/XI5/MM5_g
+ N_VDD_XI28/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI5/MM4 N_XI28/XI5/NET33_XI28/XI5/MM4_d N_XI28/XI5/NET34_XI28/XI5/MM4_g
+ N_VDD_XI28/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI5/MM10 N_XI28/XI5/NET35_XI28/XI5/MM10_d N_XI28/XI5/NET36_XI28/XI5/MM10_g
+ N_VDD_XI28/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI5/MM11 N_XI28/XI5/NET36_XI28/XI5/MM11_d N_XI28/XI5/NET35_XI28/XI5/MM11_g
+ N_VDD_XI28/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI6/MM2 N_XI28/XI6/NET34_XI28/XI6/MM2_d N_XI28/XI6/NET33_XI28/XI6/MM2_g
+ N_VSS_XI28/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM3 N_XI28/XI6/NET33_XI28/XI6/MM3_d N_WL<52>_XI28/XI6/MM3_g
+ N_BLN<9>_XI28/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM0 N_XI28/XI6/NET34_XI28/XI6/MM0_d N_WL<52>_XI28/XI6/MM0_g
+ N_BL<9>_XI28/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM1 N_XI28/XI6/NET33_XI28/XI6/MM1_d N_XI28/XI6/NET34_XI28/XI6/MM1_g
+ N_VSS_XI28/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM9 N_XI28/XI6/NET36_XI28/XI6/MM9_d N_WL<53>_XI28/XI6/MM9_g
+ N_BL<9>_XI28/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM6 N_XI28/XI6/NET35_XI28/XI6/MM6_d N_XI28/XI6/NET36_XI28/XI6/MM6_g
+ N_VSS_XI28/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM7 N_XI28/XI6/NET36_XI28/XI6/MM7_d N_XI28/XI6/NET35_XI28/XI6/MM7_g
+ N_VSS_XI28/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM8 N_XI28/XI6/NET35_XI28/XI6/MM8_d N_WL<53>_XI28/XI6/MM8_g
+ N_BLN<9>_XI28/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI6/MM5 N_XI28/XI6/NET34_XI28/XI6/MM5_d N_XI28/XI6/NET33_XI28/XI6/MM5_g
+ N_VDD_XI28/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI6/MM4 N_XI28/XI6/NET33_XI28/XI6/MM4_d N_XI28/XI6/NET34_XI28/XI6/MM4_g
+ N_VDD_XI28/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI6/MM10 N_XI28/XI6/NET35_XI28/XI6/MM10_d N_XI28/XI6/NET36_XI28/XI6/MM10_g
+ N_VDD_XI28/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI6/MM11 N_XI28/XI6/NET36_XI28/XI6/MM11_d N_XI28/XI6/NET35_XI28/XI6/MM11_g
+ N_VDD_XI28/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI7/MM2 N_XI28/XI7/NET34_XI28/XI7/MM2_d N_XI28/XI7/NET33_XI28/XI7/MM2_g
+ N_VSS_XI28/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM3 N_XI28/XI7/NET33_XI28/XI7/MM3_d N_WL<52>_XI28/XI7/MM3_g
+ N_BLN<8>_XI28/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM0 N_XI28/XI7/NET34_XI28/XI7/MM0_d N_WL<52>_XI28/XI7/MM0_g
+ N_BL<8>_XI28/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM1 N_XI28/XI7/NET33_XI28/XI7/MM1_d N_XI28/XI7/NET34_XI28/XI7/MM1_g
+ N_VSS_XI28/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM9 N_XI28/XI7/NET36_XI28/XI7/MM9_d N_WL<53>_XI28/XI7/MM9_g
+ N_BL<8>_XI28/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM6 N_XI28/XI7/NET35_XI28/XI7/MM6_d N_XI28/XI7/NET36_XI28/XI7/MM6_g
+ N_VSS_XI28/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM7 N_XI28/XI7/NET36_XI28/XI7/MM7_d N_XI28/XI7/NET35_XI28/XI7/MM7_g
+ N_VSS_XI28/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM8 N_XI28/XI7/NET35_XI28/XI7/MM8_d N_WL<53>_XI28/XI7/MM8_g
+ N_BLN<8>_XI28/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI7/MM5 N_XI28/XI7/NET34_XI28/XI7/MM5_d N_XI28/XI7/NET33_XI28/XI7/MM5_g
+ N_VDD_XI28/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI7/MM4 N_XI28/XI7/NET33_XI28/XI7/MM4_d N_XI28/XI7/NET34_XI28/XI7/MM4_g
+ N_VDD_XI28/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI7/MM10 N_XI28/XI7/NET35_XI28/XI7/MM10_d N_XI28/XI7/NET36_XI28/XI7/MM10_g
+ N_VDD_XI28/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI7/MM11 N_XI28/XI7/NET36_XI28/XI7/MM11_d N_XI28/XI7/NET35_XI28/XI7/MM11_g
+ N_VDD_XI28/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI8/MM2 N_XI28/XI8/NET34_XI28/XI8/MM2_d N_XI28/XI8/NET33_XI28/XI8/MM2_g
+ N_VSS_XI28/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM3 N_XI28/XI8/NET33_XI28/XI8/MM3_d N_WL<52>_XI28/XI8/MM3_g
+ N_BLN<7>_XI28/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM0 N_XI28/XI8/NET34_XI28/XI8/MM0_d N_WL<52>_XI28/XI8/MM0_g
+ N_BL<7>_XI28/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM1 N_XI28/XI8/NET33_XI28/XI8/MM1_d N_XI28/XI8/NET34_XI28/XI8/MM1_g
+ N_VSS_XI28/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM9 N_XI28/XI8/NET36_XI28/XI8/MM9_d N_WL<53>_XI28/XI8/MM9_g
+ N_BL<7>_XI28/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM6 N_XI28/XI8/NET35_XI28/XI8/MM6_d N_XI28/XI8/NET36_XI28/XI8/MM6_g
+ N_VSS_XI28/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM7 N_XI28/XI8/NET36_XI28/XI8/MM7_d N_XI28/XI8/NET35_XI28/XI8/MM7_g
+ N_VSS_XI28/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM8 N_XI28/XI8/NET35_XI28/XI8/MM8_d N_WL<53>_XI28/XI8/MM8_g
+ N_BLN<7>_XI28/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI8/MM5 N_XI28/XI8/NET34_XI28/XI8/MM5_d N_XI28/XI8/NET33_XI28/XI8/MM5_g
+ N_VDD_XI28/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI8/MM4 N_XI28/XI8/NET33_XI28/XI8/MM4_d N_XI28/XI8/NET34_XI28/XI8/MM4_g
+ N_VDD_XI28/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI8/MM10 N_XI28/XI8/NET35_XI28/XI8/MM10_d N_XI28/XI8/NET36_XI28/XI8/MM10_g
+ N_VDD_XI28/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI8/MM11 N_XI28/XI8/NET36_XI28/XI8/MM11_d N_XI28/XI8/NET35_XI28/XI8/MM11_g
+ N_VDD_XI28/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI9/MM2 N_XI28/XI9/NET34_XI28/XI9/MM2_d N_XI28/XI9/NET33_XI28/XI9/MM2_g
+ N_VSS_XI28/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM3 N_XI28/XI9/NET33_XI28/XI9/MM3_d N_WL<52>_XI28/XI9/MM3_g
+ N_BLN<6>_XI28/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM0 N_XI28/XI9/NET34_XI28/XI9/MM0_d N_WL<52>_XI28/XI9/MM0_g
+ N_BL<6>_XI28/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM1 N_XI28/XI9/NET33_XI28/XI9/MM1_d N_XI28/XI9/NET34_XI28/XI9/MM1_g
+ N_VSS_XI28/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM9 N_XI28/XI9/NET36_XI28/XI9/MM9_d N_WL<53>_XI28/XI9/MM9_g
+ N_BL<6>_XI28/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM6 N_XI28/XI9/NET35_XI28/XI9/MM6_d N_XI28/XI9/NET36_XI28/XI9/MM6_g
+ N_VSS_XI28/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM7 N_XI28/XI9/NET36_XI28/XI9/MM7_d N_XI28/XI9/NET35_XI28/XI9/MM7_g
+ N_VSS_XI28/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM8 N_XI28/XI9/NET35_XI28/XI9/MM8_d N_WL<53>_XI28/XI9/MM8_g
+ N_BLN<6>_XI28/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI9/MM5 N_XI28/XI9/NET34_XI28/XI9/MM5_d N_XI28/XI9/NET33_XI28/XI9/MM5_g
+ N_VDD_XI28/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI9/MM4 N_XI28/XI9/NET33_XI28/XI9/MM4_d N_XI28/XI9/NET34_XI28/XI9/MM4_g
+ N_VDD_XI28/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI9/MM10 N_XI28/XI9/NET35_XI28/XI9/MM10_d N_XI28/XI9/NET36_XI28/XI9/MM10_g
+ N_VDD_XI28/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI9/MM11 N_XI28/XI9/NET36_XI28/XI9/MM11_d N_XI28/XI9/NET35_XI28/XI9/MM11_g
+ N_VDD_XI28/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI10/MM2 N_XI28/XI10/NET34_XI28/XI10/MM2_d
+ N_XI28/XI10/NET33_XI28/XI10/MM2_g N_VSS_XI28/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI10/MM3 N_XI28/XI10/NET33_XI28/XI10/MM3_d N_WL<52>_XI28/XI10/MM3_g
+ N_BLN<5>_XI28/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI10/MM0 N_XI28/XI10/NET34_XI28/XI10/MM0_d N_WL<52>_XI28/XI10/MM0_g
+ N_BL<5>_XI28/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI10/MM1 N_XI28/XI10/NET33_XI28/XI10/MM1_d
+ N_XI28/XI10/NET34_XI28/XI10/MM1_g N_VSS_XI28/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI10/MM9 N_XI28/XI10/NET36_XI28/XI10/MM9_d N_WL<53>_XI28/XI10/MM9_g
+ N_BL<5>_XI28/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI10/MM6 N_XI28/XI10/NET35_XI28/XI10/MM6_d
+ N_XI28/XI10/NET36_XI28/XI10/MM6_g N_VSS_XI28/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI10/MM7 N_XI28/XI10/NET36_XI28/XI10/MM7_d
+ N_XI28/XI10/NET35_XI28/XI10/MM7_g N_VSS_XI28/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI10/MM8 N_XI28/XI10/NET35_XI28/XI10/MM8_d N_WL<53>_XI28/XI10/MM8_g
+ N_BLN<5>_XI28/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI10/MM5 N_XI28/XI10/NET34_XI28/XI10/MM5_d
+ N_XI28/XI10/NET33_XI28/XI10/MM5_g N_VDD_XI28/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI10/MM4 N_XI28/XI10/NET33_XI28/XI10/MM4_d
+ N_XI28/XI10/NET34_XI28/XI10/MM4_g N_VDD_XI28/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI10/MM10 N_XI28/XI10/NET35_XI28/XI10/MM10_d
+ N_XI28/XI10/NET36_XI28/XI10/MM10_g N_VDD_XI28/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI10/MM11 N_XI28/XI10/NET36_XI28/XI10/MM11_d
+ N_XI28/XI10/NET35_XI28/XI10/MM11_g N_VDD_XI28/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI11/MM2 N_XI28/XI11/NET34_XI28/XI11/MM2_d
+ N_XI28/XI11/NET33_XI28/XI11/MM2_g N_VSS_XI28/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI11/MM3 N_XI28/XI11/NET33_XI28/XI11/MM3_d N_WL<52>_XI28/XI11/MM3_g
+ N_BLN<4>_XI28/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI11/MM0 N_XI28/XI11/NET34_XI28/XI11/MM0_d N_WL<52>_XI28/XI11/MM0_g
+ N_BL<4>_XI28/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI11/MM1 N_XI28/XI11/NET33_XI28/XI11/MM1_d
+ N_XI28/XI11/NET34_XI28/XI11/MM1_g N_VSS_XI28/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI11/MM9 N_XI28/XI11/NET36_XI28/XI11/MM9_d N_WL<53>_XI28/XI11/MM9_g
+ N_BL<4>_XI28/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI11/MM6 N_XI28/XI11/NET35_XI28/XI11/MM6_d
+ N_XI28/XI11/NET36_XI28/XI11/MM6_g N_VSS_XI28/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI11/MM7 N_XI28/XI11/NET36_XI28/XI11/MM7_d
+ N_XI28/XI11/NET35_XI28/XI11/MM7_g N_VSS_XI28/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI11/MM8 N_XI28/XI11/NET35_XI28/XI11/MM8_d N_WL<53>_XI28/XI11/MM8_g
+ N_BLN<4>_XI28/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI11/MM5 N_XI28/XI11/NET34_XI28/XI11/MM5_d
+ N_XI28/XI11/NET33_XI28/XI11/MM5_g N_VDD_XI28/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI11/MM4 N_XI28/XI11/NET33_XI28/XI11/MM4_d
+ N_XI28/XI11/NET34_XI28/XI11/MM4_g N_VDD_XI28/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI11/MM10 N_XI28/XI11/NET35_XI28/XI11/MM10_d
+ N_XI28/XI11/NET36_XI28/XI11/MM10_g N_VDD_XI28/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI11/MM11 N_XI28/XI11/NET36_XI28/XI11/MM11_d
+ N_XI28/XI11/NET35_XI28/XI11/MM11_g N_VDD_XI28/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI12/MM2 N_XI28/XI12/NET34_XI28/XI12/MM2_d
+ N_XI28/XI12/NET33_XI28/XI12/MM2_g N_VSS_XI28/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI12/MM3 N_XI28/XI12/NET33_XI28/XI12/MM3_d N_WL<52>_XI28/XI12/MM3_g
+ N_BLN<3>_XI28/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI12/MM0 N_XI28/XI12/NET34_XI28/XI12/MM0_d N_WL<52>_XI28/XI12/MM0_g
+ N_BL<3>_XI28/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI12/MM1 N_XI28/XI12/NET33_XI28/XI12/MM1_d
+ N_XI28/XI12/NET34_XI28/XI12/MM1_g N_VSS_XI28/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI12/MM9 N_XI28/XI12/NET36_XI28/XI12/MM9_d N_WL<53>_XI28/XI12/MM9_g
+ N_BL<3>_XI28/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI12/MM6 N_XI28/XI12/NET35_XI28/XI12/MM6_d
+ N_XI28/XI12/NET36_XI28/XI12/MM6_g N_VSS_XI28/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI12/MM7 N_XI28/XI12/NET36_XI28/XI12/MM7_d
+ N_XI28/XI12/NET35_XI28/XI12/MM7_g N_VSS_XI28/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI12/MM8 N_XI28/XI12/NET35_XI28/XI12/MM8_d N_WL<53>_XI28/XI12/MM8_g
+ N_BLN<3>_XI28/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI12/MM5 N_XI28/XI12/NET34_XI28/XI12/MM5_d
+ N_XI28/XI12/NET33_XI28/XI12/MM5_g N_VDD_XI28/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI12/MM4 N_XI28/XI12/NET33_XI28/XI12/MM4_d
+ N_XI28/XI12/NET34_XI28/XI12/MM4_g N_VDD_XI28/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI12/MM10 N_XI28/XI12/NET35_XI28/XI12/MM10_d
+ N_XI28/XI12/NET36_XI28/XI12/MM10_g N_VDD_XI28/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI12/MM11 N_XI28/XI12/NET36_XI28/XI12/MM11_d
+ N_XI28/XI12/NET35_XI28/XI12/MM11_g N_VDD_XI28/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI13/MM2 N_XI28/XI13/NET34_XI28/XI13/MM2_d
+ N_XI28/XI13/NET33_XI28/XI13/MM2_g N_VSS_XI28/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI13/MM3 N_XI28/XI13/NET33_XI28/XI13/MM3_d N_WL<52>_XI28/XI13/MM3_g
+ N_BLN<2>_XI28/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI13/MM0 N_XI28/XI13/NET34_XI28/XI13/MM0_d N_WL<52>_XI28/XI13/MM0_g
+ N_BL<2>_XI28/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI13/MM1 N_XI28/XI13/NET33_XI28/XI13/MM1_d
+ N_XI28/XI13/NET34_XI28/XI13/MM1_g N_VSS_XI28/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI13/MM9 N_XI28/XI13/NET36_XI28/XI13/MM9_d N_WL<53>_XI28/XI13/MM9_g
+ N_BL<2>_XI28/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI13/MM6 N_XI28/XI13/NET35_XI28/XI13/MM6_d
+ N_XI28/XI13/NET36_XI28/XI13/MM6_g N_VSS_XI28/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI13/MM7 N_XI28/XI13/NET36_XI28/XI13/MM7_d
+ N_XI28/XI13/NET35_XI28/XI13/MM7_g N_VSS_XI28/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI13/MM8 N_XI28/XI13/NET35_XI28/XI13/MM8_d N_WL<53>_XI28/XI13/MM8_g
+ N_BLN<2>_XI28/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI13/MM5 N_XI28/XI13/NET34_XI28/XI13/MM5_d
+ N_XI28/XI13/NET33_XI28/XI13/MM5_g N_VDD_XI28/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI13/MM4 N_XI28/XI13/NET33_XI28/XI13/MM4_d
+ N_XI28/XI13/NET34_XI28/XI13/MM4_g N_VDD_XI28/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI13/MM10 N_XI28/XI13/NET35_XI28/XI13/MM10_d
+ N_XI28/XI13/NET36_XI28/XI13/MM10_g N_VDD_XI28/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI13/MM11 N_XI28/XI13/NET36_XI28/XI13/MM11_d
+ N_XI28/XI13/NET35_XI28/XI13/MM11_g N_VDD_XI28/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI14/MM2 N_XI28/XI14/NET34_XI28/XI14/MM2_d
+ N_XI28/XI14/NET33_XI28/XI14/MM2_g N_VSS_XI28/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI14/MM3 N_XI28/XI14/NET33_XI28/XI14/MM3_d N_WL<52>_XI28/XI14/MM3_g
+ N_BLN<1>_XI28/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI14/MM0 N_XI28/XI14/NET34_XI28/XI14/MM0_d N_WL<52>_XI28/XI14/MM0_g
+ N_BL<1>_XI28/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI14/MM1 N_XI28/XI14/NET33_XI28/XI14/MM1_d
+ N_XI28/XI14/NET34_XI28/XI14/MM1_g N_VSS_XI28/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI14/MM9 N_XI28/XI14/NET36_XI28/XI14/MM9_d N_WL<53>_XI28/XI14/MM9_g
+ N_BL<1>_XI28/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI14/MM6 N_XI28/XI14/NET35_XI28/XI14/MM6_d
+ N_XI28/XI14/NET36_XI28/XI14/MM6_g N_VSS_XI28/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI14/MM7 N_XI28/XI14/NET36_XI28/XI14/MM7_d
+ N_XI28/XI14/NET35_XI28/XI14/MM7_g N_VSS_XI28/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI14/MM8 N_XI28/XI14/NET35_XI28/XI14/MM8_d N_WL<53>_XI28/XI14/MM8_g
+ N_BLN<1>_XI28/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI14/MM5 N_XI28/XI14/NET34_XI28/XI14/MM5_d
+ N_XI28/XI14/NET33_XI28/XI14/MM5_g N_VDD_XI28/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI14/MM4 N_XI28/XI14/NET33_XI28/XI14/MM4_d
+ N_XI28/XI14/NET34_XI28/XI14/MM4_g N_VDD_XI28/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI14/MM10 N_XI28/XI14/NET35_XI28/XI14/MM10_d
+ N_XI28/XI14/NET36_XI28/XI14/MM10_g N_VDD_XI28/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI14/MM11 N_XI28/XI14/NET36_XI28/XI14/MM11_d
+ N_XI28/XI14/NET35_XI28/XI14/MM11_g N_VDD_XI28/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI15/MM2 N_XI28/XI15/NET34_XI28/XI15/MM2_d
+ N_XI28/XI15/NET33_XI28/XI15/MM2_g N_VSS_XI28/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI15/MM3 N_XI28/XI15/NET33_XI28/XI15/MM3_d N_WL<52>_XI28/XI15/MM3_g
+ N_BLN<0>_XI28/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI15/MM0 N_XI28/XI15/NET34_XI28/XI15/MM0_d N_WL<52>_XI28/XI15/MM0_g
+ N_BL<0>_XI28/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI15/MM1 N_XI28/XI15/NET33_XI28/XI15/MM1_d
+ N_XI28/XI15/NET34_XI28/XI15/MM1_g N_VSS_XI28/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI15/MM9 N_XI28/XI15/NET36_XI28/XI15/MM9_d N_WL<53>_XI28/XI15/MM9_g
+ N_BL<0>_XI28/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI15/MM6 N_XI28/XI15/NET35_XI28/XI15/MM6_d
+ N_XI28/XI15/NET36_XI28/XI15/MM6_g N_VSS_XI28/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI15/MM7 N_XI28/XI15/NET36_XI28/XI15/MM7_d
+ N_XI28/XI15/NET35_XI28/XI15/MM7_g N_VSS_XI28/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI28/XI15/MM8 N_XI28/XI15/NET35_XI28/XI15/MM8_d N_WL<53>_XI28/XI15/MM8_g
+ N_BLN<0>_XI28/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI28/XI15/MM5 N_XI28/XI15/NET34_XI28/XI15/MM5_d
+ N_XI28/XI15/NET33_XI28/XI15/MM5_g N_VDD_XI28/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI15/MM4 N_XI28/XI15/NET33_XI28/XI15/MM4_d
+ N_XI28/XI15/NET34_XI28/XI15/MM4_g N_VDD_XI28/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI15/MM10 N_XI28/XI15/NET35_XI28/XI15/MM10_d
+ N_XI28/XI15/NET36_XI28/XI15/MM10_g N_VDD_XI28/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI28/XI15/MM11 N_XI28/XI15/NET36_XI28/XI15/MM11_d
+ N_XI28/XI15/NET35_XI28/XI15/MM11_g N_VDD_XI28/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI0/MM2 N_XI29/XI0/NET34_XI29/XI0/MM2_d N_XI29/XI0/NET33_XI29/XI0/MM2_g
+ N_VSS_XI29/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI0/MM3 N_XI29/XI0/NET33_XI29/XI0/MM3_d N_WL<54>_XI29/XI0/MM3_g
+ N_BLN<15>_XI29/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI0/MM0 N_XI29/XI0/NET34_XI29/XI0/MM0_d N_WL<54>_XI29/XI0/MM0_g
+ N_BL<15>_XI29/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI0/MM1 N_XI29/XI0/NET33_XI29/XI0/MM1_d N_XI29/XI0/NET34_XI29/XI0/MM1_g
+ N_VSS_XI29/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI0/MM9 N_XI29/XI0/NET36_XI29/XI0/MM9_d N_WL<55>_XI29/XI0/MM9_g
+ N_BL<15>_XI29/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI0/MM6 N_XI29/XI0/NET35_XI29/XI0/MM6_d N_XI29/XI0/NET36_XI29/XI0/MM6_g
+ N_VSS_XI29/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI0/MM7 N_XI29/XI0/NET36_XI29/XI0/MM7_d N_XI29/XI0/NET35_XI29/XI0/MM7_g
+ N_VSS_XI29/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI0/MM8 N_XI29/XI0/NET35_XI29/XI0/MM8_d N_WL<55>_XI29/XI0/MM8_g
+ N_BLN<15>_XI29/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI0/MM5 N_XI29/XI0/NET34_XI29/XI0/MM5_d N_XI29/XI0/NET33_XI29/XI0/MM5_g
+ N_VDD_XI29/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI0/MM4 N_XI29/XI0/NET33_XI29/XI0/MM4_d N_XI29/XI0/NET34_XI29/XI0/MM4_g
+ N_VDD_XI29/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI0/MM10 N_XI29/XI0/NET35_XI29/XI0/MM10_d N_XI29/XI0/NET36_XI29/XI0/MM10_g
+ N_VDD_XI29/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI0/MM11 N_XI29/XI0/NET36_XI29/XI0/MM11_d N_XI29/XI0/NET35_XI29/XI0/MM11_g
+ N_VDD_XI29/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI1/MM2 N_XI29/XI1/NET34_XI29/XI1/MM2_d N_XI29/XI1/NET33_XI29/XI1/MM2_g
+ N_VSS_XI29/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI1/MM3 N_XI29/XI1/NET33_XI29/XI1/MM3_d N_WL<54>_XI29/XI1/MM3_g
+ N_BLN<14>_XI29/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI1/MM0 N_XI29/XI1/NET34_XI29/XI1/MM0_d N_WL<54>_XI29/XI1/MM0_g
+ N_BL<14>_XI29/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI1/MM1 N_XI29/XI1/NET33_XI29/XI1/MM1_d N_XI29/XI1/NET34_XI29/XI1/MM1_g
+ N_VSS_XI29/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI1/MM9 N_XI29/XI1/NET36_XI29/XI1/MM9_d N_WL<55>_XI29/XI1/MM9_g
+ N_BL<14>_XI29/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI1/MM6 N_XI29/XI1/NET35_XI29/XI1/MM6_d N_XI29/XI1/NET36_XI29/XI1/MM6_g
+ N_VSS_XI29/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI1/MM7 N_XI29/XI1/NET36_XI29/XI1/MM7_d N_XI29/XI1/NET35_XI29/XI1/MM7_g
+ N_VSS_XI29/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI1/MM8 N_XI29/XI1/NET35_XI29/XI1/MM8_d N_WL<55>_XI29/XI1/MM8_g
+ N_BLN<14>_XI29/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI1/MM5 N_XI29/XI1/NET34_XI29/XI1/MM5_d N_XI29/XI1/NET33_XI29/XI1/MM5_g
+ N_VDD_XI29/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI1/MM4 N_XI29/XI1/NET33_XI29/XI1/MM4_d N_XI29/XI1/NET34_XI29/XI1/MM4_g
+ N_VDD_XI29/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI1/MM10 N_XI29/XI1/NET35_XI29/XI1/MM10_d N_XI29/XI1/NET36_XI29/XI1/MM10_g
+ N_VDD_XI29/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI1/MM11 N_XI29/XI1/NET36_XI29/XI1/MM11_d N_XI29/XI1/NET35_XI29/XI1/MM11_g
+ N_VDD_XI29/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI2/MM2 N_XI29/XI2/NET34_XI29/XI2/MM2_d N_XI29/XI2/NET33_XI29/XI2/MM2_g
+ N_VSS_XI29/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI2/MM3 N_XI29/XI2/NET33_XI29/XI2/MM3_d N_WL<54>_XI29/XI2/MM3_g
+ N_BLN<13>_XI29/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI2/MM0 N_XI29/XI2/NET34_XI29/XI2/MM0_d N_WL<54>_XI29/XI2/MM0_g
+ N_BL<13>_XI29/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI2/MM1 N_XI29/XI2/NET33_XI29/XI2/MM1_d N_XI29/XI2/NET34_XI29/XI2/MM1_g
+ N_VSS_XI29/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI2/MM9 N_XI29/XI2/NET36_XI29/XI2/MM9_d N_WL<55>_XI29/XI2/MM9_g
+ N_BL<13>_XI29/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI2/MM6 N_XI29/XI2/NET35_XI29/XI2/MM6_d N_XI29/XI2/NET36_XI29/XI2/MM6_g
+ N_VSS_XI29/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI2/MM7 N_XI29/XI2/NET36_XI29/XI2/MM7_d N_XI29/XI2/NET35_XI29/XI2/MM7_g
+ N_VSS_XI29/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI2/MM8 N_XI29/XI2/NET35_XI29/XI2/MM8_d N_WL<55>_XI29/XI2/MM8_g
+ N_BLN<13>_XI29/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI2/MM5 N_XI29/XI2/NET34_XI29/XI2/MM5_d N_XI29/XI2/NET33_XI29/XI2/MM5_g
+ N_VDD_XI29/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI2/MM4 N_XI29/XI2/NET33_XI29/XI2/MM4_d N_XI29/XI2/NET34_XI29/XI2/MM4_g
+ N_VDD_XI29/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI2/MM10 N_XI29/XI2/NET35_XI29/XI2/MM10_d N_XI29/XI2/NET36_XI29/XI2/MM10_g
+ N_VDD_XI29/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI2/MM11 N_XI29/XI2/NET36_XI29/XI2/MM11_d N_XI29/XI2/NET35_XI29/XI2/MM11_g
+ N_VDD_XI29/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI3/MM2 N_XI29/XI3/NET34_XI29/XI3/MM2_d N_XI29/XI3/NET33_XI29/XI3/MM2_g
+ N_VSS_XI29/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI3/MM3 N_XI29/XI3/NET33_XI29/XI3/MM3_d N_WL<54>_XI29/XI3/MM3_g
+ N_BLN<12>_XI29/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI3/MM0 N_XI29/XI3/NET34_XI29/XI3/MM0_d N_WL<54>_XI29/XI3/MM0_g
+ N_BL<12>_XI29/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI3/MM1 N_XI29/XI3/NET33_XI29/XI3/MM1_d N_XI29/XI3/NET34_XI29/XI3/MM1_g
+ N_VSS_XI29/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI3/MM9 N_XI29/XI3/NET36_XI29/XI3/MM9_d N_WL<55>_XI29/XI3/MM9_g
+ N_BL<12>_XI29/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI3/MM6 N_XI29/XI3/NET35_XI29/XI3/MM6_d N_XI29/XI3/NET36_XI29/XI3/MM6_g
+ N_VSS_XI29/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI3/MM7 N_XI29/XI3/NET36_XI29/XI3/MM7_d N_XI29/XI3/NET35_XI29/XI3/MM7_g
+ N_VSS_XI29/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI3/MM8 N_XI29/XI3/NET35_XI29/XI3/MM8_d N_WL<55>_XI29/XI3/MM8_g
+ N_BLN<12>_XI29/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI3/MM5 N_XI29/XI3/NET34_XI29/XI3/MM5_d N_XI29/XI3/NET33_XI29/XI3/MM5_g
+ N_VDD_XI29/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI3/MM4 N_XI29/XI3/NET33_XI29/XI3/MM4_d N_XI29/XI3/NET34_XI29/XI3/MM4_g
+ N_VDD_XI29/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI3/MM10 N_XI29/XI3/NET35_XI29/XI3/MM10_d N_XI29/XI3/NET36_XI29/XI3/MM10_g
+ N_VDD_XI29/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI3/MM11 N_XI29/XI3/NET36_XI29/XI3/MM11_d N_XI29/XI3/NET35_XI29/XI3/MM11_g
+ N_VDD_XI29/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI4/MM2 N_XI29/XI4/NET34_XI29/XI4/MM2_d N_XI29/XI4/NET33_XI29/XI4/MM2_g
+ N_VSS_XI29/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI4/MM3 N_XI29/XI4/NET33_XI29/XI4/MM3_d N_WL<54>_XI29/XI4/MM3_g
+ N_BLN<11>_XI29/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI4/MM0 N_XI29/XI4/NET34_XI29/XI4/MM0_d N_WL<54>_XI29/XI4/MM0_g
+ N_BL<11>_XI29/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI4/MM1 N_XI29/XI4/NET33_XI29/XI4/MM1_d N_XI29/XI4/NET34_XI29/XI4/MM1_g
+ N_VSS_XI29/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI4/MM9 N_XI29/XI4/NET36_XI29/XI4/MM9_d N_WL<55>_XI29/XI4/MM9_g
+ N_BL<11>_XI29/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI4/MM6 N_XI29/XI4/NET35_XI29/XI4/MM6_d N_XI29/XI4/NET36_XI29/XI4/MM6_g
+ N_VSS_XI29/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI4/MM7 N_XI29/XI4/NET36_XI29/XI4/MM7_d N_XI29/XI4/NET35_XI29/XI4/MM7_g
+ N_VSS_XI29/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI4/MM8 N_XI29/XI4/NET35_XI29/XI4/MM8_d N_WL<55>_XI29/XI4/MM8_g
+ N_BLN<11>_XI29/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI4/MM5 N_XI29/XI4/NET34_XI29/XI4/MM5_d N_XI29/XI4/NET33_XI29/XI4/MM5_g
+ N_VDD_XI29/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI4/MM4 N_XI29/XI4/NET33_XI29/XI4/MM4_d N_XI29/XI4/NET34_XI29/XI4/MM4_g
+ N_VDD_XI29/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI4/MM10 N_XI29/XI4/NET35_XI29/XI4/MM10_d N_XI29/XI4/NET36_XI29/XI4/MM10_g
+ N_VDD_XI29/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI4/MM11 N_XI29/XI4/NET36_XI29/XI4/MM11_d N_XI29/XI4/NET35_XI29/XI4/MM11_g
+ N_VDD_XI29/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI5/MM2 N_XI29/XI5/NET34_XI29/XI5/MM2_d N_XI29/XI5/NET33_XI29/XI5/MM2_g
+ N_VSS_XI29/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI5/MM3 N_XI29/XI5/NET33_XI29/XI5/MM3_d N_WL<54>_XI29/XI5/MM3_g
+ N_BLN<10>_XI29/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI5/MM0 N_XI29/XI5/NET34_XI29/XI5/MM0_d N_WL<54>_XI29/XI5/MM0_g
+ N_BL<10>_XI29/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI5/MM1 N_XI29/XI5/NET33_XI29/XI5/MM1_d N_XI29/XI5/NET34_XI29/XI5/MM1_g
+ N_VSS_XI29/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI5/MM9 N_XI29/XI5/NET36_XI29/XI5/MM9_d N_WL<55>_XI29/XI5/MM9_g
+ N_BL<10>_XI29/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI5/MM6 N_XI29/XI5/NET35_XI29/XI5/MM6_d N_XI29/XI5/NET36_XI29/XI5/MM6_g
+ N_VSS_XI29/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI5/MM7 N_XI29/XI5/NET36_XI29/XI5/MM7_d N_XI29/XI5/NET35_XI29/XI5/MM7_g
+ N_VSS_XI29/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI5/MM8 N_XI29/XI5/NET35_XI29/XI5/MM8_d N_WL<55>_XI29/XI5/MM8_g
+ N_BLN<10>_XI29/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI5/MM5 N_XI29/XI5/NET34_XI29/XI5/MM5_d N_XI29/XI5/NET33_XI29/XI5/MM5_g
+ N_VDD_XI29/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI5/MM4 N_XI29/XI5/NET33_XI29/XI5/MM4_d N_XI29/XI5/NET34_XI29/XI5/MM4_g
+ N_VDD_XI29/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI5/MM10 N_XI29/XI5/NET35_XI29/XI5/MM10_d N_XI29/XI5/NET36_XI29/XI5/MM10_g
+ N_VDD_XI29/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI5/MM11 N_XI29/XI5/NET36_XI29/XI5/MM11_d N_XI29/XI5/NET35_XI29/XI5/MM11_g
+ N_VDD_XI29/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI6/MM2 N_XI29/XI6/NET34_XI29/XI6/MM2_d N_XI29/XI6/NET33_XI29/XI6/MM2_g
+ N_VSS_XI29/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM3 N_XI29/XI6/NET33_XI29/XI6/MM3_d N_WL<54>_XI29/XI6/MM3_g
+ N_BLN<9>_XI29/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM0 N_XI29/XI6/NET34_XI29/XI6/MM0_d N_WL<54>_XI29/XI6/MM0_g
+ N_BL<9>_XI29/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM1 N_XI29/XI6/NET33_XI29/XI6/MM1_d N_XI29/XI6/NET34_XI29/XI6/MM1_g
+ N_VSS_XI29/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM9 N_XI29/XI6/NET36_XI29/XI6/MM9_d N_WL<55>_XI29/XI6/MM9_g
+ N_BL<9>_XI29/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM6 N_XI29/XI6/NET35_XI29/XI6/MM6_d N_XI29/XI6/NET36_XI29/XI6/MM6_g
+ N_VSS_XI29/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM7 N_XI29/XI6/NET36_XI29/XI6/MM7_d N_XI29/XI6/NET35_XI29/XI6/MM7_g
+ N_VSS_XI29/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM8 N_XI29/XI6/NET35_XI29/XI6/MM8_d N_WL<55>_XI29/XI6/MM8_g
+ N_BLN<9>_XI29/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI6/MM5 N_XI29/XI6/NET34_XI29/XI6/MM5_d N_XI29/XI6/NET33_XI29/XI6/MM5_g
+ N_VDD_XI29/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI6/MM4 N_XI29/XI6/NET33_XI29/XI6/MM4_d N_XI29/XI6/NET34_XI29/XI6/MM4_g
+ N_VDD_XI29/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI6/MM10 N_XI29/XI6/NET35_XI29/XI6/MM10_d N_XI29/XI6/NET36_XI29/XI6/MM10_g
+ N_VDD_XI29/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI6/MM11 N_XI29/XI6/NET36_XI29/XI6/MM11_d N_XI29/XI6/NET35_XI29/XI6/MM11_g
+ N_VDD_XI29/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI7/MM2 N_XI29/XI7/NET34_XI29/XI7/MM2_d N_XI29/XI7/NET33_XI29/XI7/MM2_g
+ N_VSS_XI29/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM3 N_XI29/XI7/NET33_XI29/XI7/MM3_d N_WL<54>_XI29/XI7/MM3_g
+ N_BLN<8>_XI29/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM0 N_XI29/XI7/NET34_XI29/XI7/MM0_d N_WL<54>_XI29/XI7/MM0_g
+ N_BL<8>_XI29/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM1 N_XI29/XI7/NET33_XI29/XI7/MM1_d N_XI29/XI7/NET34_XI29/XI7/MM1_g
+ N_VSS_XI29/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM9 N_XI29/XI7/NET36_XI29/XI7/MM9_d N_WL<55>_XI29/XI7/MM9_g
+ N_BL<8>_XI29/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM6 N_XI29/XI7/NET35_XI29/XI7/MM6_d N_XI29/XI7/NET36_XI29/XI7/MM6_g
+ N_VSS_XI29/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM7 N_XI29/XI7/NET36_XI29/XI7/MM7_d N_XI29/XI7/NET35_XI29/XI7/MM7_g
+ N_VSS_XI29/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM8 N_XI29/XI7/NET35_XI29/XI7/MM8_d N_WL<55>_XI29/XI7/MM8_g
+ N_BLN<8>_XI29/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI7/MM5 N_XI29/XI7/NET34_XI29/XI7/MM5_d N_XI29/XI7/NET33_XI29/XI7/MM5_g
+ N_VDD_XI29/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI7/MM4 N_XI29/XI7/NET33_XI29/XI7/MM4_d N_XI29/XI7/NET34_XI29/XI7/MM4_g
+ N_VDD_XI29/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI7/MM10 N_XI29/XI7/NET35_XI29/XI7/MM10_d N_XI29/XI7/NET36_XI29/XI7/MM10_g
+ N_VDD_XI29/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI7/MM11 N_XI29/XI7/NET36_XI29/XI7/MM11_d N_XI29/XI7/NET35_XI29/XI7/MM11_g
+ N_VDD_XI29/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI8/MM2 N_XI29/XI8/NET34_XI29/XI8/MM2_d N_XI29/XI8/NET33_XI29/XI8/MM2_g
+ N_VSS_XI29/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM3 N_XI29/XI8/NET33_XI29/XI8/MM3_d N_WL<54>_XI29/XI8/MM3_g
+ N_BLN<7>_XI29/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM0 N_XI29/XI8/NET34_XI29/XI8/MM0_d N_WL<54>_XI29/XI8/MM0_g
+ N_BL<7>_XI29/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM1 N_XI29/XI8/NET33_XI29/XI8/MM1_d N_XI29/XI8/NET34_XI29/XI8/MM1_g
+ N_VSS_XI29/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM9 N_XI29/XI8/NET36_XI29/XI8/MM9_d N_WL<55>_XI29/XI8/MM9_g
+ N_BL<7>_XI29/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM6 N_XI29/XI8/NET35_XI29/XI8/MM6_d N_XI29/XI8/NET36_XI29/XI8/MM6_g
+ N_VSS_XI29/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM7 N_XI29/XI8/NET36_XI29/XI8/MM7_d N_XI29/XI8/NET35_XI29/XI8/MM7_g
+ N_VSS_XI29/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM8 N_XI29/XI8/NET35_XI29/XI8/MM8_d N_WL<55>_XI29/XI8/MM8_g
+ N_BLN<7>_XI29/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI8/MM5 N_XI29/XI8/NET34_XI29/XI8/MM5_d N_XI29/XI8/NET33_XI29/XI8/MM5_g
+ N_VDD_XI29/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI8/MM4 N_XI29/XI8/NET33_XI29/XI8/MM4_d N_XI29/XI8/NET34_XI29/XI8/MM4_g
+ N_VDD_XI29/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI8/MM10 N_XI29/XI8/NET35_XI29/XI8/MM10_d N_XI29/XI8/NET36_XI29/XI8/MM10_g
+ N_VDD_XI29/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI8/MM11 N_XI29/XI8/NET36_XI29/XI8/MM11_d N_XI29/XI8/NET35_XI29/XI8/MM11_g
+ N_VDD_XI29/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI9/MM2 N_XI29/XI9/NET34_XI29/XI9/MM2_d N_XI29/XI9/NET33_XI29/XI9/MM2_g
+ N_VSS_XI29/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM3 N_XI29/XI9/NET33_XI29/XI9/MM3_d N_WL<54>_XI29/XI9/MM3_g
+ N_BLN<6>_XI29/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM0 N_XI29/XI9/NET34_XI29/XI9/MM0_d N_WL<54>_XI29/XI9/MM0_g
+ N_BL<6>_XI29/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM1 N_XI29/XI9/NET33_XI29/XI9/MM1_d N_XI29/XI9/NET34_XI29/XI9/MM1_g
+ N_VSS_XI29/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM9 N_XI29/XI9/NET36_XI29/XI9/MM9_d N_WL<55>_XI29/XI9/MM9_g
+ N_BL<6>_XI29/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM6 N_XI29/XI9/NET35_XI29/XI9/MM6_d N_XI29/XI9/NET36_XI29/XI9/MM6_g
+ N_VSS_XI29/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM7 N_XI29/XI9/NET36_XI29/XI9/MM7_d N_XI29/XI9/NET35_XI29/XI9/MM7_g
+ N_VSS_XI29/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM8 N_XI29/XI9/NET35_XI29/XI9/MM8_d N_WL<55>_XI29/XI9/MM8_g
+ N_BLN<6>_XI29/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI9/MM5 N_XI29/XI9/NET34_XI29/XI9/MM5_d N_XI29/XI9/NET33_XI29/XI9/MM5_g
+ N_VDD_XI29/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI9/MM4 N_XI29/XI9/NET33_XI29/XI9/MM4_d N_XI29/XI9/NET34_XI29/XI9/MM4_g
+ N_VDD_XI29/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI9/MM10 N_XI29/XI9/NET35_XI29/XI9/MM10_d N_XI29/XI9/NET36_XI29/XI9/MM10_g
+ N_VDD_XI29/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI9/MM11 N_XI29/XI9/NET36_XI29/XI9/MM11_d N_XI29/XI9/NET35_XI29/XI9/MM11_g
+ N_VDD_XI29/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI10/MM2 N_XI29/XI10/NET34_XI29/XI10/MM2_d
+ N_XI29/XI10/NET33_XI29/XI10/MM2_g N_VSS_XI29/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI10/MM3 N_XI29/XI10/NET33_XI29/XI10/MM3_d N_WL<54>_XI29/XI10/MM3_g
+ N_BLN<5>_XI29/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI10/MM0 N_XI29/XI10/NET34_XI29/XI10/MM0_d N_WL<54>_XI29/XI10/MM0_g
+ N_BL<5>_XI29/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI10/MM1 N_XI29/XI10/NET33_XI29/XI10/MM1_d
+ N_XI29/XI10/NET34_XI29/XI10/MM1_g N_VSS_XI29/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI10/MM9 N_XI29/XI10/NET36_XI29/XI10/MM9_d N_WL<55>_XI29/XI10/MM9_g
+ N_BL<5>_XI29/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI10/MM6 N_XI29/XI10/NET35_XI29/XI10/MM6_d
+ N_XI29/XI10/NET36_XI29/XI10/MM6_g N_VSS_XI29/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI10/MM7 N_XI29/XI10/NET36_XI29/XI10/MM7_d
+ N_XI29/XI10/NET35_XI29/XI10/MM7_g N_VSS_XI29/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI10/MM8 N_XI29/XI10/NET35_XI29/XI10/MM8_d N_WL<55>_XI29/XI10/MM8_g
+ N_BLN<5>_XI29/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI10/MM5 N_XI29/XI10/NET34_XI29/XI10/MM5_d
+ N_XI29/XI10/NET33_XI29/XI10/MM5_g N_VDD_XI29/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI10/MM4 N_XI29/XI10/NET33_XI29/XI10/MM4_d
+ N_XI29/XI10/NET34_XI29/XI10/MM4_g N_VDD_XI29/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI10/MM10 N_XI29/XI10/NET35_XI29/XI10/MM10_d
+ N_XI29/XI10/NET36_XI29/XI10/MM10_g N_VDD_XI29/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI10/MM11 N_XI29/XI10/NET36_XI29/XI10/MM11_d
+ N_XI29/XI10/NET35_XI29/XI10/MM11_g N_VDD_XI29/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI11/MM2 N_XI29/XI11/NET34_XI29/XI11/MM2_d
+ N_XI29/XI11/NET33_XI29/XI11/MM2_g N_VSS_XI29/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI11/MM3 N_XI29/XI11/NET33_XI29/XI11/MM3_d N_WL<54>_XI29/XI11/MM3_g
+ N_BLN<4>_XI29/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI11/MM0 N_XI29/XI11/NET34_XI29/XI11/MM0_d N_WL<54>_XI29/XI11/MM0_g
+ N_BL<4>_XI29/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI11/MM1 N_XI29/XI11/NET33_XI29/XI11/MM1_d
+ N_XI29/XI11/NET34_XI29/XI11/MM1_g N_VSS_XI29/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI11/MM9 N_XI29/XI11/NET36_XI29/XI11/MM9_d N_WL<55>_XI29/XI11/MM9_g
+ N_BL<4>_XI29/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI11/MM6 N_XI29/XI11/NET35_XI29/XI11/MM6_d
+ N_XI29/XI11/NET36_XI29/XI11/MM6_g N_VSS_XI29/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI11/MM7 N_XI29/XI11/NET36_XI29/XI11/MM7_d
+ N_XI29/XI11/NET35_XI29/XI11/MM7_g N_VSS_XI29/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI11/MM8 N_XI29/XI11/NET35_XI29/XI11/MM8_d N_WL<55>_XI29/XI11/MM8_g
+ N_BLN<4>_XI29/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI11/MM5 N_XI29/XI11/NET34_XI29/XI11/MM5_d
+ N_XI29/XI11/NET33_XI29/XI11/MM5_g N_VDD_XI29/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI11/MM4 N_XI29/XI11/NET33_XI29/XI11/MM4_d
+ N_XI29/XI11/NET34_XI29/XI11/MM4_g N_VDD_XI29/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI11/MM10 N_XI29/XI11/NET35_XI29/XI11/MM10_d
+ N_XI29/XI11/NET36_XI29/XI11/MM10_g N_VDD_XI29/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI11/MM11 N_XI29/XI11/NET36_XI29/XI11/MM11_d
+ N_XI29/XI11/NET35_XI29/XI11/MM11_g N_VDD_XI29/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI12/MM2 N_XI29/XI12/NET34_XI29/XI12/MM2_d
+ N_XI29/XI12/NET33_XI29/XI12/MM2_g N_VSS_XI29/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI12/MM3 N_XI29/XI12/NET33_XI29/XI12/MM3_d N_WL<54>_XI29/XI12/MM3_g
+ N_BLN<3>_XI29/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI12/MM0 N_XI29/XI12/NET34_XI29/XI12/MM0_d N_WL<54>_XI29/XI12/MM0_g
+ N_BL<3>_XI29/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI12/MM1 N_XI29/XI12/NET33_XI29/XI12/MM1_d
+ N_XI29/XI12/NET34_XI29/XI12/MM1_g N_VSS_XI29/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI12/MM9 N_XI29/XI12/NET36_XI29/XI12/MM9_d N_WL<55>_XI29/XI12/MM9_g
+ N_BL<3>_XI29/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI12/MM6 N_XI29/XI12/NET35_XI29/XI12/MM6_d
+ N_XI29/XI12/NET36_XI29/XI12/MM6_g N_VSS_XI29/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI12/MM7 N_XI29/XI12/NET36_XI29/XI12/MM7_d
+ N_XI29/XI12/NET35_XI29/XI12/MM7_g N_VSS_XI29/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI12/MM8 N_XI29/XI12/NET35_XI29/XI12/MM8_d N_WL<55>_XI29/XI12/MM8_g
+ N_BLN<3>_XI29/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI12/MM5 N_XI29/XI12/NET34_XI29/XI12/MM5_d
+ N_XI29/XI12/NET33_XI29/XI12/MM5_g N_VDD_XI29/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI12/MM4 N_XI29/XI12/NET33_XI29/XI12/MM4_d
+ N_XI29/XI12/NET34_XI29/XI12/MM4_g N_VDD_XI29/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI12/MM10 N_XI29/XI12/NET35_XI29/XI12/MM10_d
+ N_XI29/XI12/NET36_XI29/XI12/MM10_g N_VDD_XI29/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI12/MM11 N_XI29/XI12/NET36_XI29/XI12/MM11_d
+ N_XI29/XI12/NET35_XI29/XI12/MM11_g N_VDD_XI29/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI13/MM2 N_XI29/XI13/NET34_XI29/XI13/MM2_d
+ N_XI29/XI13/NET33_XI29/XI13/MM2_g N_VSS_XI29/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI13/MM3 N_XI29/XI13/NET33_XI29/XI13/MM3_d N_WL<54>_XI29/XI13/MM3_g
+ N_BLN<2>_XI29/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI13/MM0 N_XI29/XI13/NET34_XI29/XI13/MM0_d N_WL<54>_XI29/XI13/MM0_g
+ N_BL<2>_XI29/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI13/MM1 N_XI29/XI13/NET33_XI29/XI13/MM1_d
+ N_XI29/XI13/NET34_XI29/XI13/MM1_g N_VSS_XI29/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI13/MM9 N_XI29/XI13/NET36_XI29/XI13/MM9_d N_WL<55>_XI29/XI13/MM9_g
+ N_BL<2>_XI29/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI13/MM6 N_XI29/XI13/NET35_XI29/XI13/MM6_d
+ N_XI29/XI13/NET36_XI29/XI13/MM6_g N_VSS_XI29/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI13/MM7 N_XI29/XI13/NET36_XI29/XI13/MM7_d
+ N_XI29/XI13/NET35_XI29/XI13/MM7_g N_VSS_XI29/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI13/MM8 N_XI29/XI13/NET35_XI29/XI13/MM8_d N_WL<55>_XI29/XI13/MM8_g
+ N_BLN<2>_XI29/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI13/MM5 N_XI29/XI13/NET34_XI29/XI13/MM5_d
+ N_XI29/XI13/NET33_XI29/XI13/MM5_g N_VDD_XI29/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI13/MM4 N_XI29/XI13/NET33_XI29/XI13/MM4_d
+ N_XI29/XI13/NET34_XI29/XI13/MM4_g N_VDD_XI29/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI13/MM10 N_XI29/XI13/NET35_XI29/XI13/MM10_d
+ N_XI29/XI13/NET36_XI29/XI13/MM10_g N_VDD_XI29/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI13/MM11 N_XI29/XI13/NET36_XI29/XI13/MM11_d
+ N_XI29/XI13/NET35_XI29/XI13/MM11_g N_VDD_XI29/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI14/MM2 N_XI29/XI14/NET34_XI29/XI14/MM2_d
+ N_XI29/XI14/NET33_XI29/XI14/MM2_g N_VSS_XI29/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI14/MM3 N_XI29/XI14/NET33_XI29/XI14/MM3_d N_WL<54>_XI29/XI14/MM3_g
+ N_BLN<1>_XI29/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI14/MM0 N_XI29/XI14/NET34_XI29/XI14/MM0_d N_WL<54>_XI29/XI14/MM0_g
+ N_BL<1>_XI29/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI14/MM1 N_XI29/XI14/NET33_XI29/XI14/MM1_d
+ N_XI29/XI14/NET34_XI29/XI14/MM1_g N_VSS_XI29/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI14/MM9 N_XI29/XI14/NET36_XI29/XI14/MM9_d N_WL<55>_XI29/XI14/MM9_g
+ N_BL<1>_XI29/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI14/MM6 N_XI29/XI14/NET35_XI29/XI14/MM6_d
+ N_XI29/XI14/NET36_XI29/XI14/MM6_g N_VSS_XI29/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI14/MM7 N_XI29/XI14/NET36_XI29/XI14/MM7_d
+ N_XI29/XI14/NET35_XI29/XI14/MM7_g N_VSS_XI29/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI14/MM8 N_XI29/XI14/NET35_XI29/XI14/MM8_d N_WL<55>_XI29/XI14/MM8_g
+ N_BLN<1>_XI29/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI14/MM5 N_XI29/XI14/NET34_XI29/XI14/MM5_d
+ N_XI29/XI14/NET33_XI29/XI14/MM5_g N_VDD_XI29/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI14/MM4 N_XI29/XI14/NET33_XI29/XI14/MM4_d
+ N_XI29/XI14/NET34_XI29/XI14/MM4_g N_VDD_XI29/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI14/MM10 N_XI29/XI14/NET35_XI29/XI14/MM10_d
+ N_XI29/XI14/NET36_XI29/XI14/MM10_g N_VDD_XI29/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI14/MM11 N_XI29/XI14/NET36_XI29/XI14/MM11_d
+ N_XI29/XI14/NET35_XI29/XI14/MM11_g N_VDD_XI29/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI15/MM2 N_XI29/XI15/NET34_XI29/XI15/MM2_d
+ N_XI29/XI15/NET33_XI29/XI15/MM2_g N_VSS_XI29/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI15/MM3 N_XI29/XI15/NET33_XI29/XI15/MM3_d N_WL<54>_XI29/XI15/MM3_g
+ N_BLN<0>_XI29/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI15/MM0 N_XI29/XI15/NET34_XI29/XI15/MM0_d N_WL<54>_XI29/XI15/MM0_g
+ N_BL<0>_XI29/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI15/MM1 N_XI29/XI15/NET33_XI29/XI15/MM1_d
+ N_XI29/XI15/NET34_XI29/XI15/MM1_g N_VSS_XI29/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI15/MM9 N_XI29/XI15/NET36_XI29/XI15/MM9_d N_WL<55>_XI29/XI15/MM9_g
+ N_BL<0>_XI29/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI15/MM6 N_XI29/XI15/NET35_XI29/XI15/MM6_d
+ N_XI29/XI15/NET36_XI29/XI15/MM6_g N_VSS_XI29/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI15/MM7 N_XI29/XI15/NET36_XI29/XI15/MM7_d
+ N_XI29/XI15/NET35_XI29/XI15/MM7_g N_VSS_XI29/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI29/XI15/MM8 N_XI29/XI15/NET35_XI29/XI15/MM8_d N_WL<55>_XI29/XI15/MM8_g
+ N_BLN<0>_XI29/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI29/XI15/MM5 N_XI29/XI15/NET34_XI29/XI15/MM5_d
+ N_XI29/XI15/NET33_XI29/XI15/MM5_g N_VDD_XI29/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI15/MM4 N_XI29/XI15/NET33_XI29/XI15/MM4_d
+ N_XI29/XI15/NET34_XI29/XI15/MM4_g N_VDD_XI29/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI15/MM10 N_XI29/XI15/NET35_XI29/XI15/MM10_d
+ N_XI29/XI15/NET36_XI29/XI15/MM10_g N_VDD_XI29/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI29/XI15/MM11 N_XI29/XI15/NET36_XI29/XI15/MM11_d
+ N_XI29/XI15/NET35_XI29/XI15/MM11_g N_VDD_XI29/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI0/MM2 N_XI30/XI0/NET34_XI30/XI0/MM2_d N_XI30/XI0/NET33_XI30/XI0/MM2_g
+ N_VSS_XI30/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI0/MM3 N_XI30/XI0/NET33_XI30/XI0/MM3_d N_WL<56>_XI30/XI0/MM3_g
+ N_BLN<15>_XI30/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI0/MM0 N_XI30/XI0/NET34_XI30/XI0/MM0_d N_WL<56>_XI30/XI0/MM0_g
+ N_BL<15>_XI30/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI0/MM1 N_XI30/XI0/NET33_XI30/XI0/MM1_d N_XI30/XI0/NET34_XI30/XI0/MM1_g
+ N_VSS_XI30/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI0/MM9 N_XI30/XI0/NET36_XI30/XI0/MM9_d N_WL<57>_XI30/XI0/MM9_g
+ N_BL<15>_XI30/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI0/MM6 N_XI30/XI0/NET35_XI30/XI0/MM6_d N_XI30/XI0/NET36_XI30/XI0/MM6_g
+ N_VSS_XI30/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI0/MM7 N_XI30/XI0/NET36_XI30/XI0/MM7_d N_XI30/XI0/NET35_XI30/XI0/MM7_g
+ N_VSS_XI30/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI0/MM8 N_XI30/XI0/NET35_XI30/XI0/MM8_d N_WL<57>_XI30/XI0/MM8_g
+ N_BLN<15>_XI30/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI0/MM5 N_XI30/XI0/NET34_XI30/XI0/MM5_d N_XI30/XI0/NET33_XI30/XI0/MM5_g
+ N_VDD_XI30/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI0/MM4 N_XI30/XI0/NET33_XI30/XI0/MM4_d N_XI30/XI0/NET34_XI30/XI0/MM4_g
+ N_VDD_XI30/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI0/MM10 N_XI30/XI0/NET35_XI30/XI0/MM10_d N_XI30/XI0/NET36_XI30/XI0/MM10_g
+ N_VDD_XI30/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI0/MM11 N_XI30/XI0/NET36_XI30/XI0/MM11_d N_XI30/XI0/NET35_XI30/XI0/MM11_g
+ N_VDD_XI30/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI1/MM2 N_XI30/XI1/NET34_XI30/XI1/MM2_d N_XI30/XI1/NET33_XI30/XI1/MM2_g
+ N_VSS_XI30/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI1/MM3 N_XI30/XI1/NET33_XI30/XI1/MM3_d N_WL<56>_XI30/XI1/MM3_g
+ N_BLN<14>_XI30/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI1/MM0 N_XI30/XI1/NET34_XI30/XI1/MM0_d N_WL<56>_XI30/XI1/MM0_g
+ N_BL<14>_XI30/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI1/MM1 N_XI30/XI1/NET33_XI30/XI1/MM1_d N_XI30/XI1/NET34_XI30/XI1/MM1_g
+ N_VSS_XI30/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI1/MM9 N_XI30/XI1/NET36_XI30/XI1/MM9_d N_WL<57>_XI30/XI1/MM9_g
+ N_BL<14>_XI30/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI1/MM6 N_XI30/XI1/NET35_XI30/XI1/MM6_d N_XI30/XI1/NET36_XI30/XI1/MM6_g
+ N_VSS_XI30/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI1/MM7 N_XI30/XI1/NET36_XI30/XI1/MM7_d N_XI30/XI1/NET35_XI30/XI1/MM7_g
+ N_VSS_XI30/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI1/MM8 N_XI30/XI1/NET35_XI30/XI1/MM8_d N_WL<57>_XI30/XI1/MM8_g
+ N_BLN<14>_XI30/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI1/MM5 N_XI30/XI1/NET34_XI30/XI1/MM5_d N_XI30/XI1/NET33_XI30/XI1/MM5_g
+ N_VDD_XI30/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI1/MM4 N_XI30/XI1/NET33_XI30/XI1/MM4_d N_XI30/XI1/NET34_XI30/XI1/MM4_g
+ N_VDD_XI30/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI1/MM10 N_XI30/XI1/NET35_XI30/XI1/MM10_d N_XI30/XI1/NET36_XI30/XI1/MM10_g
+ N_VDD_XI30/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI1/MM11 N_XI30/XI1/NET36_XI30/XI1/MM11_d N_XI30/XI1/NET35_XI30/XI1/MM11_g
+ N_VDD_XI30/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI2/MM2 N_XI30/XI2/NET34_XI30/XI2/MM2_d N_XI30/XI2/NET33_XI30/XI2/MM2_g
+ N_VSS_XI30/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI2/MM3 N_XI30/XI2/NET33_XI30/XI2/MM3_d N_WL<56>_XI30/XI2/MM3_g
+ N_BLN<13>_XI30/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI2/MM0 N_XI30/XI2/NET34_XI30/XI2/MM0_d N_WL<56>_XI30/XI2/MM0_g
+ N_BL<13>_XI30/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI2/MM1 N_XI30/XI2/NET33_XI30/XI2/MM1_d N_XI30/XI2/NET34_XI30/XI2/MM1_g
+ N_VSS_XI30/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI2/MM9 N_XI30/XI2/NET36_XI30/XI2/MM9_d N_WL<57>_XI30/XI2/MM9_g
+ N_BL<13>_XI30/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI2/MM6 N_XI30/XI2/NET35_XI30/XI2/MM6_d N_XI30/XI2/NET36_XI30/XI2/MM6_g
+ N_VSS_XI30/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI2/MM7 N_XI30/XI2/NET36_XI30/XI2/MM7_d N_XI30/XI2/NET35_XI30/XI2/MM7_g
+ N_VSS_XI30/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI2/MM8 N_XI30/XI2/NET35_XI30/XI2/MM8_d N_WL<57>_XI30/XI2/MM8_g
+ N_BLN<13>_XI30/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI2/MM5 N_XI30/XI2/NET34_XI30/XI2/MM5_d N_XI30/XI2/NET33_XI30/XI2/MM5_g
+ N_VDD_XI30/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI2/MM4 N_XI30/XI2/NET33_XI30/XI2/MM4_d N_XI30/XI2/NET34_XI30/XI2/MM4_g
+ N_VDD_XI30/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI2/MM10 N_XI30/XI2/NET35_XI30/XI2/MM10_d N_XI30/XI2/NET36_XI30/XI2/MM10_g
+ N_VDD_XI30/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI2/MM11 N_XI30/XI2/NET36_XI30/XI2/MM11_d N_XI30/XI2/NET35_XI30/XI2/MM11_g
+ N_VDD_XI30/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI3/MM2 N_XI30/XI3/NET34_XI30/XI3/MM2_d N_XI30/XI3/NET33_XI30/XI3/MM2_g
+ N_VSS_XI30/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI3/MM3 N_XI30/XI3/NET33_XI30/XI3/MM3_d N_WL<56>_XI30/XI3/MM3_g
+ N_BLN<12>_XI30/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI3/MM0 N_XI30/XI3/NET34_XI30/XI3/MM0_d N_WL<56>_XI30/XI3/MM0_g
+ N_BL<12>_XI30/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI3/MM1 N_XI30/XI3/NET33_XI30/XI3/MM1_d N_XI30/XI3/NET34_XI30/XI3/MM1_g
+ N_VSS_XI30/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI3/MM9 N_XI30/XI3/NET36_XI30/XI3/MM9_d N_WL<57>_XI30/XI3/MM9_g
+ N_BL<12>_XI30/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI3/MM6 N_XI30/XI3/NET35_XI30/XI3/MM6_d N_XI30/XI3/NET36_XI30/XI3/MM6_g
+ N_VSS_XI30/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI3/MM7 N_XI30/XI3/NET36_XI30/XI3/MM7_d N_XI30/XI3/NET35_XI30/XI3/MM7_g
+ N_VSS_XI30/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI3/MM8 N_XI30/XI3/NET35_XI30/XI3/MM8_d N_WL<57>_XI30/XI3/MM8_g
+ N_BLN<12>_XI30/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI3/MM5 N_XI30/XI3/NET34_XI30/XI3/MM5_d N_XI30/XI3/NET33_XI30/XI3/MM5_g
+ N_VDD_XI30/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI3/MM4 N_XI30/XI3/NET33_XI30/XI3/MM4_d N_XI30/XI3/NET34_XI30/XI3/MM4_g
+ N_VDD_XI30/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI3/MM10 N_XI30/XI3/NET35_XI30/XI3/MM10_d N_XI30/XI3/NET36_XI30/XI3/MM10_g
+ N_VDD_XI30/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI3/MM11 N_XI30/XI3/NET36_XI30/XI3/MM11_d N_XI30/XI3/NET35_XI30/XI3/MM11_g
+ N_VDD_XI30/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI4/MM2 N_XI30/XI4/NET34_XI30/XI4/MM2_d N_XI30/XI4/NET33_XI30/XI4/MM2_g
+ N_VSS_XI30/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI4/MM3 N_XI30/XI4/NET33_XI30/XI4/MM3_d N_WL<56>_XI30/XI4/MM3_g
+ N_BLN<11>_XI30/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI4/MM0 N_XI30/XI4/NET34_XI30/XI4/MM0_d N_WL<56>_XI30/XI4/MM0_g
+ N_BL<11>_XI30/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI4/MM1 N_XI30/XI4/NET33_XI30/XI4/MM1_d N_XI30/XI4/NET34_XI30/XI4/MM1_g
+ N_VSS_XI30/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI4/MM9 N_XI30/XI4/NET36_XI30/XI4/MM9_d N_WL<57>_XI30/XI4/MM9_g
+ N_BL<11>_XI30/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI4/MM6 N_XI30/XI4/NET35_XI30/XI4/MM6_d N_XI30/XI4/NET36_XI30/XI4/MM6_g
+ N_VSS_XI30/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI4/MM7 N_XI30/XI4/NET36_XI30/XI4/MM7_d N_XI30/XI4/NET35_XI30/XI4/MM7_g
+ N_VSS_XI30/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI4/MM8 N_XI30/XI4/NET35_XI30/XI4/MM8_d N_WL<57>_XI30/XI4/MM8_g
+ N_BLN<11>_XI30/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI4/MM5 N_XI30/XI4/NET34_XI30/XI4/MM5_d N_XI30/XI4/NET33_XI30/XI4/MM5_g
+ N_VDD_XI30/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI4/MM4 N_XI30/XI4/NET33_XI30/XI4/MM4_d N_XI30/XI4/NET34_XI30/XI4/MM4_g
+ N_VDD_XI30/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI4/MM10 N_XI30/XI4/NET35_XI30/XI4/MM10_d N_XI30/XI4/NET36_XI30/XI4/MM10_g
+ N_VDD_XI30/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI4/MM11 N_XI30/XI4/NET36_XI30/XI4/MM11_d N_XI30/XI4/NET35_XI30/XI4/MM11_g
+ N_VDD_XI30/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI5/MM2 N_XI30/XI5/NET34_XI30/XI5/MM2_d N_XI30/XI5/NET33_XI30/XI5/MM2_g
+ N_VSS_XI30/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI5/MM3 N_XI30/XI5/NET33_XI30/XI5/MM3_d N_WL<56>_XI30/XI5/MM3_g
+ N_BLN<10>_XI30/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI5/MM0 N_XI30/XI5/NET34_XI30/XI5/MM0_d N_WL<56>_XI30/XI5/MM0_g
+ N_BL<10>_XI30/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI5/MM1 N_XI30/XI5/NET33_XI30/XI5/MM1_d N_XI30/XI5/NET34_XI30/XI5/MM1_g
+ N_VSS_XI30/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI5/MM9 N_XI30/XI5/NET36_XI30/XI5/MM9_d N_WL<57>_XI30/XI5/MM9_g
+ N_BL<10>_XI30/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI5/MM6 N_XI30/XI5/NET35_XI30/XI5/MM6_d N_XI30/XI5/NET36_XI30/XI5/MM6_g
+ N_VSS_XI30/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI5/MM7 N_XI30/XI5/NET36_XI30/XI5/MM7_d N_XI30/XI5/NET35_XI30/XI5/MM7_g
+ N_VSS_XI30/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI5/MM8 N_XI30/XI5/NET35_XI30/XI5/MM8_d N_WL<57>_XI30/XI5/MM8_g
+ N_BLN<10>_XI30/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI5/MM5 N_XI30/XI5/NET34_XI30/XI5/MM5_d N_XI30/XI5/NET33_XI30/XI5/MM5_g
+ N_VDD_XI30/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI5/MM4 N_XI30/XI5/NET33_XI30/XI5/MM4_d N_XI30/XI5/NET34_XI30/XI5/MM4_g
+ N_VDD_XI30/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI5/MM10 N_XI30/XI5/NET35_XI30/XI5/MM10_d N_XI30/XI5/NET36_XI30/XI5/MM10_g
+ N_VDD_XI30/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI5/MM11 N_XI30/XI5/NET36_XI30/XI5/MM11_d N_XI30/XI5/NET35_XI30/XI5/MM11_g
+ N_VDD_XI30/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI6/MM2 N_XI30/XI6/NET34_XI30/XI6/MM2_d N_XI30/XI6/NET33_XI30/XI6/MM2_g
+ N_VSS_XI30/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM3 N_XI30/XI6/NET33_XI30/XI6/MM3_d N_WL<56>_XI30/XI6/MM3_g
+ N_BLN<9>_XI30/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM0 N_XI30/XI6/NET34_XI30/XI6/MM0_d N_WL<56>_XI30/XI6/MM0_g
+ N_BL<9>_XI30/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM1 N_XI30/XI6/NET33_XI30/XI6/MM1_d N_XI30/XI6/NET34_XI30/XI6/MM1_g
+ N_VSS_XI30/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM9 N_XI30/XI6/NET36_XI30/XI6/MM9_d N_WL<57>_XI30/XI6/MM9_g
+ N_BL<9>_XI30/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM6 N_XI30/XI6/NET35_XI30/XI6/MM6_d N_XI30/XI6/NET36_XI30/XI6/MM6_g
+ N_VSS_XI30/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM7 N_XI30/XI6/NET36_XI30/XI6/MM7_d N_XI30/XI6/NET35_XI30/XI6/MM7_g
+ N_VSS_XI30/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM8 N_XI30/XI6/NET35_XI30/XI6/MM8_d N_WL<57>_XI30/XI6/MM8_g
+ N_BLN<9>_XI30/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI6/MM5 N_XI30/XI6/NET34_XI30/XI6/MM5_d N_XI30/XI6/NET33_XI30/XI6/MM5_g
+ N_VDD_XI30/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI6/MM4 N_XI30/XI6/NET33_XI30/XI6/MM4_d N_XI30/XI6/NET34_XI30/XI6/MM4_g
+ N_VDD_XI30/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI6/MM10 N_XI30/XI6/NET35_XI30/XI6/MM10_d N_XI30/XI6/NET36_XI30/XI6/MM10_g
+ N_VDD_XI30/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI6/MM11 N_XI30/XI6/NET36_XI30/XI6/MM11_d N_XI30/XI6/NET35_XI30/XI6/MM11_g
+ N_VDD_XI30/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI7/MM2 N_XI30/XI7/NET34_XI30/XI7/MM2_d N_XI30/XI7/NET33_XI30/XI7/MM2_g
+ N_VSS_XI30/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM3 N_XI30/XI7/NET33_XI30/XI7/MM3_d N_WL<56>_XI30/XI7/MM3_g
+ N_BLN<8>_XI30/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM0 N_XI30/XI7/NET34_XI30/XI7/MM0_d N_WL<56>_XI30/XI7/MM0_g
+ N_BL<8>_XI30/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM1 N_XI30/XI7/NET33_XI30/XI7/MM1_d N_XI30/XI7/NET34_XI30/XI7/MM1_g
+ N_VSS_XI30/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM9 N_XI30/XI7/NET36_XI30/XI7/MM9_d N_WL<57>_XI30/XI7/MM9_g
+ N_BL<8>_XI30/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM6 N_XI30/XI7/NET35_XI30/XI7/MM6_d N_XI30/XI7/NET36_XI30/XI7/MM6_g
+ N_VSS_XI30/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM7 N_XI30/XI7/NET36_XI30/XI7/MM7_d N_XI30/XI7/NET35_XI30/XI7/MM7_g
+ N_VSS_XI30/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM8 N_XI30/XI7/NET35_XI30/XI7/MM8_d N_WL<57>_XI30/XI7/MM8_g
+ N_BLN<8>_XI30/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI7/MM5 N_XI30/XI7/NET34_XI30/XI7/MM5_d N_XI30/XI7/NET33_XI30/XI7/MM5_g
+ N_VDD_XI30/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI7/MM4 N_XI30/XI7/NET33_XI30/XI7/MM4_d N_XI30/XI7/NET34_XI30/XI7/MM4_g
+ N_VDD_XI30/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI7/MM10 N_XI30/XI7/NET35_XI30/XI7/MM10_d N_XI30/XI7/NET36_XI30/XI7/MM10_g
+ N_VDD_XI30/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI7/MM11 N_XI30/XI7/NET36_XI30/XI7/MM11_d N_XI30/XI7/NET35_XI30/XI7/MM11_g
+ N_VDD_XI30/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI8/MM2 N_XI30/XI8/NET34_XI30/XI8/MM2_d N_XI30/XI8/NET33_XI30/XI8/MM2_g
+ N_VSS_XI30/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM3 N_XI30/XI8/NET33_XI30/XI8/MM3_d N_WL<56>_XI30/XI8/MM3_g
+ N_BLN<7>_XI30/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM0 N_XI30/XI8/NET34_XI30/XI8/MM0_d N_WL<56>_XI30/XI8/MM0_g
+ N_BL<7>_XI30/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM1 N_XI30/XI8/NET33_XI30/XI8/MM1_d N_XI30/XI8/NET34_XI30/XI8/MM1_g
+ N_VSS_XI30/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM9 N_XI30/XI8/NET36_XI30/XI8/MM9_d N_WL<57>_XI30/XI8/MM9_g
+ N_BL<7>_XI30/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM6 N_XI30/XI8/NET35_XI30/XI8/MM6_d N_XI30/XI8/NET36_XI30/XI8/MM6_g
+ N_VSS_XI30/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM7 N_XI30/XI8/NET36_XI30/XI8/MM7_d N_XI30/XI8/NET35_XI30/XI8/MM7_g
+ N_VSS_XI30/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM8 N_XI30/XI8/NET35_XI30/XI8/MM8_d N_WL<57>_XI30/XI8/MM8_g
+ N_BLN<7>_XI30/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI8/MM5 N_XI30/XI8/NET34_XI30/XI8/MM5_d N_XI30/XI8/NET33_XI30/XI8/MM5_g
+ N_VDD_XI30/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI8/MM4 N_XI30/XI8/NET33_XI30/XI8/MM4_d N_XI30/XI8/NET34_XI30/XI8/MM4_g
+ N_VDD_XI30/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI8/MM10 N_XI30/XI8/NET35_XI30/XI8/MM10_d N_XI30/XI8/NET36_XI30/XI8/MM10_g
+ N_VDD_XI30/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI8/MM11 N_XI30/XI8/NET36_XI30/XI8/MM11_d N_XI30/XI8/NET35_XI30/XI8/MM11_g
+ N_VDD_XI30/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI9/MM2 N_XI30/XI9/NET34_XI30/XI9/MM2_d N_XI30/XI9/NET33_XI30/XI9/MM2_g
+ N_VSS_XI30/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM3 N_XI30/XI9/NET33_XI30/XI9/MM3_d N_WL<56>_XI30/XI9/MM3_g
+ N_BLN<6>_XI30/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM0 N_XI30/XI9/NET34_XI30/XI9/MM0_d N_WL<56>_XI30/XI9/MM0_g
+ N_BL<6>_XI30/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM1 N_XI30/XI9/NET33_XI30/XI9/MM1_d N_XI30/XI9/NET34_XI30/XI9/MM1_g
+ N_VSS_XI30/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM9 N_XI30/XI9/NET36_XI30/XI9/MM9_d N_WL<57>_XI30/XI9/MM9_g
+ N_BL<6>_XI30/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM6 N_XI30/XI9/NET35_XI30/XI9/MM6_d N_XI30/XI9/NET36_XI30/XI9/MM6_g
+ N_VSS_XI30/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM7 N_XI30/XI9/NET36_XI30/XI9/MM7_d N_XI30/XI9/NET35_XI30/XI9/MM7_g
+ N_VSS_XI30/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM8 N_XI30/XI9/NET35_XI30/XI9/MM8_d N_WL<57>_XI30/XI9/MM8_g
+ N_BLN<6>_XI30/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI9/MM5 N_XI30/XI9/NET34_XI30/XI9/MM5_d N_XI30/XI9/NET33_XI30/XI9/MM5_g
+ N_VDD_XI30/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI9/MM4 N_XI30/XI9/NET33_XI30/XI9/MM4_d N_XI30/XI9/NET34_XI30/XI9/MM4_g
+ N_VDD_XI30/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI9/MM10 N_XI30/XI9/NET35_XI30/XI9/MM10_d N_XI30/XI9/NET36_XI30/XI9/MM10_g
+ N_VDD_XI30/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI9/MM11 N_XI30/XI9/NET36_XI30/XI9/MM11_d N_XI30/XI9/NET35_XI30/XI9/MM11_g
+ N_VDD_XI30/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI10/MM2 N_XI30/XI10/NET34_XI30/XI10/MM2_d
+ N_XI30/XI10/NET33_XI30/XI10/MM2_g N_VSS_XI30/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI10/MM3 N_XI30/XI10/NET33_XI30/XI10/MM3_d N_WL<56>_XI30/XI10/MM3_g
+ N_BLN<5>_XI30/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI10/MM0 N_XI30/XI10/NET34_XI30/XI10/MM0_d N_WL<56>_XI30/XI10/MM0_g
+ N_BL<5>_XI30/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI10/MM1 N_XI30/XI10/NET33_XI30/XI10/MM1_d
+ N_XI30/XI10/NET34_XI30/XI10/MM1_g N_VSS_XI30/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI10/MM9 N_XI30/XI10/NET36_XI30/XI10/MM9_d N_WL<57>_XI30/XI10/MM9_g
+ N_BL<5>_XI30/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI10/MM6 N_XI30/XI10/NET35_XI30/XI10/MM6_d
+ N_XI30/XI10/NET36_XI30/XI10/MM6_g N_VSS_XI30/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI10/MM7 N_XI30/XI10/NET36_XI30/XI10/MM7_d
+ N_XI30/XI10/NET35_XI30/XI10/MM7_g N_VSS_XI30/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI10/MM8 N_XI30/XI10/NET35_XI30/XI10/MM8_d N_WL<57>_XI30/XI10/MM8_g
+ N_BLN<5>_XI30/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI10/MM5 N_XI30/XI10/NET34_XI30/XI10/MM5_d
+ N_XI30/XI10/NET33_XI30/XI10/MM5_g N_VDD_XI30/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI10/MM4 N_XI30/XI10/NET33_XI30/XI10/MM4_d
+ N_XI30/XI10/NET34_XI30/XI10/MM4_g N_VDD_XI30/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI10/MM10 N_XI30/XI10/NET35_XI30/XI10/MM10_d
+ N_XI30/XI10/NET36_XI30/XI10/MM10_g N_VDD_XI30/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI10/MM11 N_XI30/XI10/NET36_XI30/XI10/MM11_d
+ N_XI30/XI10/NET35_XI30/XI10/MM11_g N_VDD_XI30/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI11/MM2 N_XI30/XI11/NET34_XI30/XI11/MM2_d
+ N_XI30/XI11/NET33_XI30/XI11/MM2_g N_VSS_XI30/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI11/MM3 N_XI30/XI11/NET33_XI30/XI11/MM3_d N_WL<56>_XI30/XI11/MM3_g
+ N_BLN<4>_XI30/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI11/MM0 N_XI30/XI11/NET34_XI30/XI11/MM0_d N_WL<56>_XI30/XI11/MM0_g
+ N_BL<4>_XI30/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI11/MM1 N_XI30/XI11/NET33_XI30/XI11/MM1_d
+ N_XI30/XI11/NET34_XI30/XI11/MM1_g N_VSS_XI30/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI11/MM9 N_XI30/XI11/NET36_XI30/XI11/MM9_d N_WL<57>_XI30/XI11/MM9_g
+ N_BL<4>_XI30/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI11/MM6 N_XI30/XI11/NET35_XI30/XI11/MM6_d
+ N_XI30/XI11/NET36_XI30/XI11/MM6_g N_VSS_XI30/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI11/MM7 N_XI30/XI11/NET36_XI30/XI11/MM7_d
+ N_XI30/XI11/NET35_XI30/XI11/MM7_g N_VSS_XI30/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI11/MM8 N_XI30/XI11/NET35_XI30/XI11/MM8_d N_WL<57>_XI30/XI11/MM8_g
+ N_BLN<4>_XI30/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI11/MM5 N_XI30/XI11/NET34_XI30/XI11/MM5_d
+ N_XI30/XI11/NET33_XI30/XI11/MM5_g N_VDD_XI30/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI11/MM4 N_XI30/XI11/NET33_XI30/XI11/MM4_d
+ N_XI30/XI11/NET34_XI30/XI11/MM4_g N_VDD_XI30/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI11/MM10 N_XI30/XI11/NET35_XI30/XI11/MM10_d
+ N_XI30/XI11/NET36_XI30/XI11/MM10_g N_VDD_XI30/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI11/MM11 N_XI30/XI11/NET36_XI30/XI11/MM11_d
+ N_XI30/XI11/NET35_XI30/XI11/MM11_g N_VDD_XI30/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI12/MM2 N_XI30/XI12/NET34_XI30/XI12/MM2_d
+ N_XI30/XI12/NET33_XI30/XI12/MM2_g N_VSS_XI30/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI12/MM3 N_XI30/XI12/NET33_XI30/XI12/MM3_d N_WL<56>_XI30/XI12/MM3_g
+ N_BLN<3>_XI30/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI12/MM0 N_XI30/XI12/NET34_XI30/XI12/MM0_d N_WL<56>_XI30/XI12/MM0_g
+ N_BL<3>_XI30/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI12/MM1 N_XI30/XI12/NET33_XI30/XI12/MM1_d
+ N_XI30/XI12/NET34_XI30/XI12/MM1_g N_VSS_XI30/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI12/MM9 N_XI30/XI12/NET36_XI30/XI12/MM9_d N_WL<57>_XI30/XI12/MM9_g
+ N_BL<3>_XI30/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI12/MM6 N_XI30/XI12/NET35_XI30/XI12/MM6_d
+ N_XI30/XI12/NET36_XI30/XI12/MM6_g N_VSS_XI30/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI12/MM7 N_XI30/XI12/NET36_XI30/XI12/MM7_d
+ N_XI30/XI12/NET35_XI30/XI12/MM7_g N_VSS_XI30/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI12/MM8 N_XI30/XI12/NET35_XI30/XI12/MM8_d N_WL<57>_XI30/XI12/MM8_g
+ N_BLN<3>_XI30/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI12/MM5 N_XI30/XI12/NET34_XI30/XI12/MM5_d
+ N_XI30/XI12/NET33_XI30/XI12/MM5_g N_VDD_XI30/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI12/MM4 N_XI30/XI12/NET33_XI30/XI12/MM4_d
+ N_XI30/XI12/NET34_XI30/XI12/MM4_g N_VDD_XI30/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI12/MM10 N_XI30/XI12/NET35_XI30/XI12/MM10_d
+ N_XI30/XI12/NET36_XI30/XI12/MM10_g N_VDD_XI30/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI12/MM11 N_XI30/XI12/NET36_XI30/XI12/MM11_d
+ N_XI30/XI12/NET35_XI30/XI12/MM11_g N_VDD_XI30/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI13/MM2 N_XI30/XI13/NET34_XI30/XI13/MM2_d
+ N_XI30/XI13/NET33_XI30/XI13/MM2_g N_VSS_XI30/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI13/MM3 N_XI30/XI13/NET33_XI30/XI13/MM3_d N_WL<56>_XI30/XI13/MM3_g
+ N_BLN<2>_XI30/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI13/MM0 N_XI30/XI13/NET34_XI30/XI13/MM0_d N_WL<56>_XI30/XI13/MM0_g
+ N_BL<2>_XI30/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI13/MM1 N_XI30/XI13/NET33_XI30/XI13/MM1_d
+ N_XI30/XI13/NET34_XI30/XI13/MM1_g N_VSS_XI30/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI13/MM9 N_XI30/XI13/NET36_XI30/XI13/MM9_d N_WL<57>_XI30/XI13/MM9_g
+ N_BL<2>_XI30/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI13/MM6 N_XI30/XI13/NET35_XI30/XI13/MM6_d
+ N_XI30/XI13/NET36_XI30/XI13/MM6_g N_VSS_XI30/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI13/MM7 N_XI30/XI13/NET36_XI30/XI13/MM7_d
+ N_XI30/XI13/NET35_XI30/XI13/MM7_g N_VSS_XI30/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI13/MM8 N_XI30/XI13/NET35_XI30/XI13/MM8_d N_WL<57>_XI30/XI13/MM8_g
+ N_BLN<2>_XI30/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI13/MM5 N_XI30/XI13/NET34_XI30/XI13/MM5_d
+ N_XI30/XI13/NET33_XI30/XI13/MM5_g N_VDD_XI30/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI13/MM4 N_XI30/XI13/NET33_XI30/XI13/MM4_d
+ N_XI30/XI13/NET34_XI30/XI13/MM4_g N_VDD_XI30/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI13/MM10 N_XI30/XI13/NET35_XI30/XI13/MM10_d
+ N_XI30/XI13/NET36_XI30/XI13/MM10_g N_VDD_XI30/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI13/MM11 N_XI30/XI13/NET36_XI30/XI13/MM11_d
+ N_XI30/XI13/NET35_XI30/XI13/MM11_g N_VDD_XI30/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI14/MM2 N_XI30/XI14/NET34_XI30/XI14/MM2_d
+ N_XI30/XI14/NET33_XI30/XI14/MM2_g N_VSS_XI30/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI14/MM3 N_XI30/XI14/NET33_XI30/XI14/MM3_d N_WL<56>_XI30/XI14/MM3_g
+ N_BLN<1>_XI30/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI14/MM0 N_XI30/XI14/NET34_XI30/XI14/MM0_d N_WL<56>_XI30/XI14/MM0_g
+ N_BL<1>_XI30/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI14/MM1 N_XI30/XI14/NET33_XI30/XI14/MM1_d
+ N_XI30/XI14/NET34_XI30/XI14/MM1_g N_VSS_XI30/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI14/MM9 N_XI30/XI14/NET36_XI30/XI14/MM9_d N_WL<57>_XI30/XI14/MM9_g
+ N_BL<1>_XI30/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI14/MM6 N_XI30/XI14/NET35_XI30/XI14/MM6_d
+ N_XI30/XI14/NET36_XI30/XI14/MM6_g N_VSS_XI30/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI14/MM7 N_XI30/XI14/NET36_XI30/XI14/MM7_d
+ N_XI30/XI14/NET35_XI30/XI14/MM7_g N_VSS_XI30/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI14/MM8 N_XI30/XI14/NET35_XI30/XI14/MM8_d N_WL<57>_XI30/XI14/MM8_g
+ N_BLN<1>_XI30/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI14/MM5 N_XI30/XI14/NET34_XI30/XI14/MM5_d
+ N_XI30/XI14/NET33_XI30/XI14/MM5_g N_VDD_XI30/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI14/MM4 N_XI30/XI14/NET33_XI30/XI14/MM4_d
+ N_XI30/XI14/NET34_XI30/XI14/MM4_g N_VDD_XI30/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI14/MM10 N_XI30/XI14/NET35_XI30/XI14/MM10_d
+ N_XI30/XI14/NET36_XI30/XI14/MM10_g N_VDD_XI30/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI14/MM11 N_XI30/XI14/NET36_XI30/XI14/MM11_d
+ N_XI30/XI14/NET35_XI30/XI14/MM11_g N_VDD_XI30/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI15/MM2 N_XI30/XI15/NET34_XI30/XI15/MM2_d
+ N_XI30/XI15/NET33_XI30/XI15/MM2_g N_VSS_XI30/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI15/MM3 N_XI30/XI15/NET33_XI30/XI15/MM3_d N_WL<56>_XI30/XI15/MM3_g
+ N_BLN<0>_XI30/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI15/MM0 N_XI30/XI15/NET34_XI30/XI15/MM0_d N_WL<56>_XI30/XI15/MM0_g
+ N_BL<0>_XI30/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI15/MM1 N_XI30/XI15/NET33_XI30/XI15/MM1_d
+ N_XI30/XI15/NET34_XI30/XI15/MM1_g N_VSS_XI30/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI15/MM9 N_XI30/XI15/NET36_XI30/XI15/MM9_d N_WL<57>_XI30/XI15/MM9_g
+ N_BL<0>_XI30/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI15/MM6 N_XI30/XI15/NET35_XI30/XI15/MM6_d
+ N_XI30/XI15/NET36_XI30/XI15/MM6_g N_VSS_XI30/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI15/MM7 N_XI30/XI15/NET36_XI30/XI15/MM7_d
+ N_XI30/XI15/NET35_XI30/XI15/MM7_g N_VSS_XI30/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI30/XI15/MM8 N_XI30/XI15/NET35_XI30/XI15/MM8_d N_WL<57>_XI30/XI15/MM8_g
+ N_BLN<0>_XI30/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI30/XI15/MM5 N_XI30/XI15/NET34_XI30/XI15/MM5_d
+ N_XI30/XI15/NET33_XI30/XI15/MM5_g N_VDD_XI30/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI15/MM4 N_XI30/XI15/NET33_XI30/XI15/MM4_d
+ N_XI30/XI15/NET34_XI30/XI15/MM4_g N_VDD_XI30/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI15/MM10 N_XI30/XI15/NET35_XI30/XI15/MM10_d
+ N_XI30/XI15/NET36_XI30/XI15/MM10_g N_VDD_XI30/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI30/XI15/MM11 N_XI30/XI15/NET36_XI30/XI15/MM11_d
+ N_XI30/XI15/NET35_XI30/XI15/MM11_g N_VDD_XI30/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI0/MM2 N_XI31/XI0/NET34_XI31/XI0/MM2_d N_XI31/XI0/NET33_XI31/XI0/MM2_g
+ N_VSS_XI31/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI0/MM3 N_XI31/XI0/NET33_XI31/XI0/MM3_d N_WL<58>_XI31/XI0/MM3_g
+ N_BLN<15>_XI31/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI0/MM0 N_XI31/XI0/NET34_XI31/XI0/MM0_d N_WL<58>_XI31/XI0/MM0_g
+ N_BL<15>_XI31/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI0/MM1 N_XI31/XI0/NET33_XI31/XI0/MM1_d N_XI31/XI0/NET34_XI31/XI0/MM1_g
+ N_VSS_XI31/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI0/MM9 N_XI31/XI0/NET36_XI31/XI0/MM9_d N_WL<59>_XI31/XI0/MM9_g
+ N_BL<15>_XI31/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI0/MM6 N_XI31/XI0/NET35_XI31/XI0/MM6_d N_XI31/XI0/NET36_XI31/XI0/MM6_g
+ N_VSS_XI31/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI0/MM7 N_XI31/XI0/NET36_XI31/XI0/MM7_d N_XI31/XI0/NET35_XI31/XI0/MM7_g
+ N_VSS_XI31/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI0/MM8 N_XI31/XI0/NET35_XI31/XI0/MM8_d N_WL<59>_XI31/XI0/MM8_g
+ N_BLN<15>_XI31/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI0/MM5 N_XI31/XI0/NET34_XI31/XI0/MM5_d N_XI31/XI0/NET33_XI31/XI0/MM5_g
+ N_VDD_XI31/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI0/MM4 N_XI31/XI0/NET33_XI31/XI0/MM4_d N_XI31/XI0/NET34_XI31/XI0/MM4_g
+ N_VDD_XI31/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI0/MM10 N_XI31/XI0/NET35_XI31/XI0/MM10_d N_XI31/XI0/NET36_XI31/XI0/MM10_g
+ N_VDD_XI31/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI0/MM11 N_XI31/XI0/NET36_XI31/XI0/MM11_d N_XI31/XI0/NET35_XI31/XI0/MM11_g
+ N_VDD_XI31/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI1/MM2 N_XI31/XI1/NET34_XI31/XI1/MM2_d N_XI31/XI1/NET33_XI31/XI1/MM2_g
+ N_VSS_XI31/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI1/MM3 N_XI31/XI1/NET33_XI31/XI1/MM3_d N_WL<58>_XI31/XI1/MM3_g
+ N_BLN<14>_XI31/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI1/MM0 N_XI31/XI1/NET34_XI31/XI1/MM0_d N_WL<58>_XI31/XI1/MM0_g
+ N_BL<14>_XI31/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI1/MM1 N_XI31/XI1/NET33_XI31/XI1/MM1_d N_XI31/XI1/NET34_XI31/XI1/MM1_g
+ N_VSS_XI31/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI1/MM9 N_XI31/XI1/NET36_XI31/XI1/MM9_d N_WL<59>_XI31/XI1/MM9_g
+ N_BL<14>_XI31/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI1/MM6 N_XI31/XI1/NET35_XI31/XI1/MM6_d N_XI31/XI1/NET36_XI31/XI1/MM6_g
+ N_VSS_XI31/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI1/MM7 N_XI31/XI1/NET36_XI31/XI1/MM7_d N_XI31/XI1/NET35_XI31/XI1/MM7_g
+ N_VSS_XI31/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI1/MM8 N_XI31/XI1/NET35_XI31/XI1/MM8_d N_WL<59>_XI31/XI1/MM8_g
+ N_BLN<14>_XI31/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI1/MM5 N_XI31/XI1/NET34_XI31/XI1/MM5_d N_XI31/XI1/NET33_XI31/XI1/MM5_g
+ N_VDD_XI31/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI1/MM4 N_XI31/XI1/NET33_XI31/XI1/MM4_d N_XI31/XI1/NET34_XI31/XI1/MM4_g
+ N_VDD_XI31/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI1/MM10 N_XI31/XI1/NET35_XI31/XI1/MM10_d N_XI31/XI1/NET36_XI31/XI1/MM10_g
+ N_VDD_XI31/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI1/MM11 N_XI31/XI1/NET36_XI31/XI1/MM11_d N_XI31/XI1/NET35_XI31/XI1/MM11_g
+ N_VDD_XI31/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI2/MM2 N_XI31/XI2/NET34_XI31/XI2/MM2_d N_XI31/XI2/NET33_XI31/XI2/MM2_g
+ N_VSS_XI31/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI2/MM3 N_XI31/XI2/NET33_XI31/XI2/MM3_d N_WL<58>_XI31/XI2/MM3_g
+ N_BLN<13>_XI31/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI2/MM0 N_XI31/XI2/NET34_XI31/XI2/MM0_d N_WL<58>_XI31/XI2/MM0_g
+ N_BL<13>_XI31/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI2/MM1 N_XI31/XI2/NET33_XI31/XI2/MM1_d N_XI31/XI2/NET34_XI31/XI2/MM1_g
+ N_VSS_XI31/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI2/MM9 N_XI31/XI2/NET36_XI31/XI2/MM9_d N_WL<59>_XI31/XI2/MM9_g
+ N_BL<13>_XI31/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI2/MM6 N_XI31/XI2/NET35_XI31/XI2/MM6_d N_XI31/XI2/NET36_XI31/XI2/MM6_g
+ N_VSS_XI31/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI2/MM7 N_XI31/XI2/NET36_XI31/XI2/MM7_d N_XI31/XI2/NET35_XI31/XI2/MM7_g
+ N_VSS_XI31/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI2/MM8 N_XI31/XI2/NET35_XI31/XI2/MM8_d N_WL<59>_XI31/XI2/MM8_g
+ N_BLN<13>_XI31/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI2/MM5 N_XI31/XI2/NET34_XI31/XI2/MM5_d N_XI31/XI2/NET33_XI31/XI2/MM5_g
+ N_VDD_XI31/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI2/MM4 N_XI31/XI2/NET33_XI31/XI2/MM4_d N_XI31/XI2/NET34_XI31/XI2/MM4_g
+ N_VDD_XI31/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI2/MM10 N_XI31/XI2/NET35_XI31/XI2/MM10_d N_XI31/XI2/NET36_XI31/XI2/MM10_g
+ N_VDD_XI31/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI2/MM11 N_XI31/XI2/NET36_XI31/XI2/MM11_d N_XI31/XI2/NET35_XI31/XI2/MM11_g
+ N_VDD_XI31/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI3/MM2 N_XI31/XI3/NET34_XI31/XI3/MM2_d N_XI31/XI3/NET33_XI31/XI3/MM2_g
+ N_VSS_XI31/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI3/MM3 N_XI31/XI3/NET33_XI31/XI3/MM3_d N_WL<58>_XI31/XI3/MM3_g
+ N_BLN<12>_XI31/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI3/MM0 N_XI31/XI3/NET34_XI31/XI3/MM0_d N_WL<58>_XI31/XI3/MM0_g
+ N_BL<12>_XI31/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI3/MM1 N_XI31/XI3/NET33_XI31/XI3/MM1_d N_XI31/XI3/NET34_XI31/XI3/MM1_g
+ N_VSS_XI31/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI3/MM9 N_XI31/XI3/NET36_XI31/XI3/MM9_d N_WL<59>_XI31/XI3/MM9_g
+ N_BL<12>_XI31/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI3/MM6 N_XI31/XI3/NET35_XI31/XI3/MM6_d N_XI31/XI3/NET36_XI31/XI3/MM6_g
+ N_VSS_XI31/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI3/MM7 N_XI31/XI3/NET36_XI31/XI3/MM7_d N_XI31/XI3/NET35_XI31/XI3/MM7_g
+ N_VSS_XI31/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI3/MM8 N_XI31/XI3/NET35_XI31/XI3/MM8_d N_WL<59>_XI31/XI3/MM8_g
+ N_BLN<12>_XI31/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI3/MM5 N_XI31/XI3/NET34_XI31/XI3/MM5_d N_XI31/XI3/NET33_XI31/XI3/MM5_g
+ N_VDD_XI31/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI3/MM4 N_XI31/XI3/NET33_XI31/XI3/MM4_d N_XI31/XI3/NET34_XI31/XI3/MM4_g
+ N_VDD_XI31/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI3/MM10 N_XI31/XI3/NET35_XI31/XI3/MM10_d N_XI31/XI3/NET36_XI31/XI3/MM10_g
+ N_VDD_XI31/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI3/MM11 N_XI31/XI3/NET36_XI31/XI3/MM11_d N_XI31/XI3/NET35_XI31/XI3/MM11_g
+ N_VDD_XI31/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI4/MM2 N_XI31/XI4/NET34_XI31/XI4/MM2_d N_XI31/XI4/NET33_XI31/XI4/MM2_g
+ N_VSS_XI31/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI4/MM3 N_XI31/XI4/NET33_XI31/XI4/MM3_d N_WL<58>_XI31/XI4/MM3_g
+ N_BLN<11>_XI31/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI4/MM0 N_XI31/XI4/NET34_XI31/XI4/MM0_d N_WL<58>_XI31/XI4/MM0_g
+ N_BL<11>_XI31/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI4/MM1 N_XI31/XI4/NET33_XI31/XI4/MM1_d N_XI31/XI4/NET34_XI31/XI4/MM1_g
+ N_VSS_XI31/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI4/MM9 N_XI31/XI4/NET36_XI31/XI4/MM9_d N_WL<59>_XI31/XI4/MM9_g
+ N_BL<11>_XI31/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI4/MM6 N_XI31/XI4/NET35_XI31/XI4/MM6_d N_XI31/XI4/NET36_XI31/XI4/MM6_g
+ N_VSS_XI31/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI4/MM7 N_XI31/XI4/NET36_XI31/XI4/MM7_d N_XI31/XI4/NET35_XI31/XI4/MM7_g
+ N_VSS_XI31/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI4/MM8 N_XI31/XI4/NET35_XI31/XI4/MM8_d N_WL<59>_XI31/XI4/MM8_g
+ N_BLN<11>_XI31/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI4/MM5 N_XI31/XI4/NET34_XI31/XI4/MM5_d N_XI31/XI4/NET33_XI31/XI4/MM5_g
+ N_VDD_XI31/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI4/MM4 N_XI31/XI4/NET33_XI31/XI4/MM4_d N_XI31/XI4/NET34_XI31/XI4/MM4_g
+ N_VDD_XI31/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI4/MM10 N_XI31/XI4/NET35_XI31/XI4/MM10_d N_XI31/XI4/NET36_XI31/XI4/MM10_g
+ N_VDD_XI31/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI4/MM11 N_XI31/XI4/NET36_XI31/XI4/MM11_d N_XI31/XI4/NET35_XI31/XI4/MM11_g
+ N_VDD_XI31/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI5/MM2 N_XI31/XI5/NET34_XI31/XI5/MM2_d N_XI31/XI5/NET33_XI31/XI5/MM2_g
+ N_VSS_XI31/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI5/MM3 N_XI31/XI5/NET33_XI31/XI5/MM3_d N_WL<58>_XI31/XI5/MM3_g
+ N_BLN<10>_XI31/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI5/MM0 N_XI31/XI5/NET34_XI31/XI5/MM0_d N_WL<58>_XI31/XI5/MM0_g
+ N_BL<10>_XI31/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI5/MM1 N_XI31/XI5/NET33_XI31/XI5/MM1_d N_XI31/XI5/NET34_XI31/XI5/MM1_g
+ N_VSS_XI31/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI5/MM9 N_XI31/XI5/NET36_XI31/XI5/MM9_d N_WL<59>_XI31/XI5/MM9_g
+ N_BL<10>_XI31/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI5/MM6 N_XI31/XI5/NET35_XI31/XI5/MM6_d N_XI31/XI5/NET36_XI31/XI5/MM6_g
+ N_VSS_XI31/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI5/MM7 N_XI31/XI5/NET36_XI31/XI5/MM7_d N_XI31/XI5/NET35_XI31/XI5/MM7_g
+ N_VSS_XI31/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI5/MM8 N_XI31/XI5/NET35_XI31/XI5/MM8_d N_WL<59>_XI31/XI5/MM8_g
+ N_BLN<10>_XI31/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI5/MM5 N_XI31/XI5/NET34_XI31/XI5/MM5_d N_XI31/XI5/NET33_XI31/XI5/MM5_g
+ N_VDD_XI31/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI5/MM4 N_XI31/XI5/NET33_XI31/XI5/MM4_d N_XI31/XI5/NET34_XI31/XI5/MM4_g
+ N_VDD_XI31/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI5/MM10 N_XI31/XI5/NET35_XI31/XI5/MM10_d N_XI31/XI5/NET36_XI31/XI5/MM10_g
+ N_VDD_XI31/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI5/MM11 N_XI31/XI5/NET36_XI31/XI5/MM11_d N_XI31/XI5/NET35_XI31/XI5/MM11_g
+ N_VDD_XI31/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI6/MM2 N_XI31/XI6/NET34_XI31/XI6/MM2_d N_XI31/XI6/NET33_XI31/XI6/MM2_g
+ N_VSS_XI31/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM3 N_XI31/XI6/NET33_XI31/XI6/MM3_d N_WL<58>_XI31/XI6/MM3_g
+ N_BLN<9>_XI31/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM0 N_XI31/XI6/NET34_XI31/XI6/MM0_d N_WL<58>_XI31/XI6/MM0_g
+ N_BL<9>_XI31/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM1 N_XI31/XI6/NET33_XI31/XI6/MM1_d N_XI31/XI6/NET34_XI31/XI6/MM1_g
+ N_VSS_XI31/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM9 N_XI31/XI6/NET36_XI31/XI6/MM9_d N_WL<59>_XI31/XI6/MM9_g
+ N_BL<9>_XI31/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM6 N_XI31/XI6/NET35_XI31/XI6/MM6_d N_XI31/XI6/NET36_XI31/XI6/MM6_g
+ N_VSS_XI31/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM7 N_XI31/XI6/NET36_XI31/XI6/MM7_d N_XI31/XI6/NET35_XI31/XI6/MM7_g
+ N_VSS_XI31/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM8 N_XI31/XI6/NET35_XI31/XI6/MM8_d N_WL<59>_XI31/XI6/MM8_g
+ N_BLN<9>_XI31/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI6/MM5 N_XI31/XI6/NET34_XI31/XI6/MM5_d N_XI31/XI6/NET33_XI31/XI6/MM5_g
+ N_VDD_XI31/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI6/MM4 N_XI31/XI6/NET33_XI31/XI6/MM4_d N_XI31/XI6/NET34_XI31/XI6/MM4_g
+ N_VDD_XI31/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI6/MM10 N_XI31/XI6/NET35_XI31/XI6/MM10_d N_XI31/XI6/NET36_XI31/XI6/MM10_g
+ N_VDD_XI31/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI6/MM11 N_XI31/XI6/NET36_XI31/XI6/MM11_d N_XI31/XI6/NET35_XI31/XI6/MM11_g
+ N_VDD_XI31/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI7/MM2 N_XI31/XI7/NET34_XI31/XI7/MM2_d N_XI31/XI7/NET33_XI31/XI7/MM2_g
+ N_VSS_XI31/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM3 N_XI31/XI7/NET33_XI31/XI7/MM3_d N_WL<58>_XI31/XI7/MM3_g
+ N_BLN<8>_XI31/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM0 N_XI31/XI7/NET34_XI31/XI7/MM0_d N_WL<58>_XI31/XI7/MM0_g
+ N_BL<8>_XI31/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM1 N_XI31/XI7/NET33_XI31/XI7/MM1_d N_XI31/XI7/NET34_XI31/XI7/MM1_g
+ N_VSS_XI31/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM9 N_XI31/XI7/NET36_XI31/XI7/MM9_d N_WL<59>_XI31/XI7/MM9_g
+ N_BL<8>_XI31/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM6 N_XI31/XI7/NET35_XI31/XI7/MM6_d N_XI31/XI7/NET36_XI31/XI7/MM6_g
+ N_VSS_XI31/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM7 N_XI31/XI7/NET36_XI31/XI7/MM7_d N_XI31/XI7/NET35_XI31/XI7/MM7_g
+ N_VSS_XI31/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM8 N_XI31/XI7/NET35_XI31/XI7/MM8_d N_WL<59>_XI31/XI7/MM8_g
+ N_BLN<8>_XI31/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI7/MM5 N_XI31/XI7/NET34_XI31/XI7/MM5_d N_XI31/XI7/NET33_XI31/XI7/MM5_g
+ N_VDD_XI31/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI7/MM4 N_XI31/XI7/NET33_XI31/XI7/MM4_d N_XI31/XI7/NET34_XI31/XI7/MM4_g
+ N_VDD_XI31/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI7/MM10 N_XI31/XI7/NET35_XI31/XI7/MM10_d N_XI31/XI7/NET36_XI31/XI7/MM10_g
+ N_VDD_XI31/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI7/MM11 N_XI31/XI7/NET36_XI31/XI7/MM11_d N_XI31/XI7/NET35_XI31/XI7/MM11_g
+ N_VDD_XI31/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI8/MM2 N_XI31/XI8/NET34_XI31/XI8/MM2_d N_XI31/XI8/NET33_XI31/XI8/MM2_g
+ N_VSS_XI31/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM3 N_XI31/XI8/NET33_XI31/XI8/MM3_d N_WL<58>_XI31/XI8/MM3_g
+ N_BLN<7>_XI31/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM0 N_XI31/XI8/NET34_XI31/XI8/MM0_d N_WL<58>_XI31/XI8/MM0_g
+ N_BL<7>_XI31/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM1 N_XI31/XI8/NET33_XI31/XI8/MM1_d N_XI31/XI8/NET34_XI31/XI8/MM1_g
+ N_VSS_XI31/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM9 N_XI31/XI8/NET36_XI31/XI8/MM9_d N_WL<59>_XI31/XI8/MM9_g
+ N_BL<7>_XI31/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM6 N_XI31/XI8/NET35_XI31/XI8/MM6_d N_XI31/XI8/NET36_XI31/XI8/MM6_g
+ N_VSS_XI31/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM7 N_XI31/XI8/NET36_XI31/XI8/MM7_d N_XI31/XI8/NET35_XI31/XI8/MM7_g
+ N_VSS_XI31/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM8 N_XI31/XI8/NET35_XI31/XI8/MM8_d N_WL<59>_XI31/XI8/MM8_g
+ N_BLN<7>_XI31/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI8/MM5 N_XI31/XI8/NET34_XI31/XI8/MM5_d N_XI31/XI8/NET33_XI31/XI8/MM5_g
+ N_VDD_XI31/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI8/MM4 N_XI31/XI8/NET33_XI31/XI8/MM4_d N_XI31/XI8/NET34_XI31/XI8/MM4_g
+ N_VDD_XI31/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI8/MM10 N_XI31/XI8/NET35_XI31/XI8/MM10_d N_XI31/XI8/NET36_XI31/XI8/MM10_g
+ N_VDD_XI31/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI8/MM11 N_XI31/XI8/NET36_XI31/XI8/MM11_d N_XI31/XI8/NET35_XI31/XI8/MM11_g
+ N_VDD_XI31/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI9/MM2 N_XI31/XI9/NET34_XI31/XI9/MM2_d N_XI31/XI9/NET33_XI31/XI9/MM2_g
+ N_VSS_XI31/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM3 N_XI31/XI9/NET33_XI31/XI9/MM3_d N_WL<58>_XI31/XI9/MM3_g
+ N_BLN<6>_XI31/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM0 N_XI31/XI9/NET34_XI31/XI9/MM0_d N_WL<58>_XI31/XI9/MM0_g
+ N_BL<6>_XI31/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM1 N_XI31/XI9/NET33_XI31/XI9/MM1_d N_XI31/XI9/NET34_XI31/XI9/MM1_g
+ N_VSS_XI31/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM9 N_XI31/XI9/NET36_XI31/XI9/MM9_d N_WL<59>_XI31/XI9/MM9_g
+ N_BL<6>_XI31/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM6 N_XI31/XI9/NET35_XI31/XI9/MM6_d N_XI31/XI9/NET36_XI31/XI9/MM6_g
+ N_VSS_XI31/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM7 N_XI31/XI9/NET36_XI31/XI9/MM7_d N_XI31/XI9/NET35_XI31/XI9/MM7_g
+ N_VSS_XI31/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM8 N_XI31/XI9/NET35_XI31/XI9/MM8_d N_WL<59>_XI31/XI9/MM8_g
+ N_BLN<6>_XI31/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI9/MM5 N_XI31/XI9/NET34_XI31/XI9/MM5_d N_XI31/XI9/NET33_XI31/XI9/MM5_g
+ N_VDD_XI31/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI9/MM4 N_XI31/XI9/NET33_XI31/XI9/MM4_d N_XI31/XI9/NET34_XI31/XI9/MM4_g
+ N_VDD_XI31/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI9/MM10 N_XI31/XI9/NET35_XI31/XI9/MM10_d N_XI31/XI9/NET36_XI31/XI9/MM10_g
+ N_VDD_XI31/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI9/MM11 N_XI31/XI9/NET36_XI31/XI9/MM11_d N_XI31/XI9/NET35_XI31/XI9/MM11_g
+ N_VDD_XI31/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI10/MM2 N_XI31/XI10/NET34_XI31/XI10/MM2_d
+ N_XI31/XI10/NET33_XI31/XI10/MM2_g N_VSS_XI31/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI10/MM3 N_XI31/XI10/NET33_XI31/XI10/MM3_d N_WL<58>_XI31/XI10/MM3_g
+ N_BLN<5>_XI31/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI10/MM0 N_XI31/XI10/NET34_XI31/XI10/MM0_d N_WL<58>_XI31/XI10/MM0_g
+ N_BL<5>_XI31/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI10/MM1 N_XI31/XI10/NET33_XI31/XI10/MM1_d
+ N_XI31/XI10/NET34_XI31/XI10/MM1_g N_VSS_XI31/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI10/MM9 N_XI31/XI10/NET36_XI31/XI10/MM9_d N_WL<59>_XI31/XI10/MM9_g
+ N_BL<5>_XI31/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI10/MM6 N_XI31/XI10/NET35_XI31/XI10/MM6_d
+ N_XI31/XI10/NET36_XI31/XI10/MM6_g N_VSS_XI31/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI10/MM7 N_XI31/XI10/NET36_XI31/XI10/MM7_d
+ N_XI31/XI10/NET35_XI31/XI10/MM7_g N_VSS_XI31/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI10/MM8 N_XI31/XI10/NET35_XI31/XI10/MM8_d N_WL<59>_XI31/XI10/MM8_g
+ N_BLN<5>_XI31/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI10/MM5 N_XI31/XI10/NET34_XI31/XI10/MM5_d
+ N_XI31/XI10/NET33_XI31/XI10/MM5_g N_VDD_XI31/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI10/MM4 N_XI31/XI10/NET33_XI31/XI10/MM4_d
+ N_XI31/XI10/NET34_XI31/XI10/MM4_g N_VDD_XI31/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI10/MM10 N_XI31/XI10/NET35_XI31/XI10/MM10_d
+ N_XI31/XI10/NET36_XI31/XI10/MM10_g N_VDD_XI31/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI10/MM11 N_XI31/XI10/NET36_XI31/XI10/MM11_d
+ N_XI31/XI10/NET35_XI31/XI10/MM11_g N_VDD_XI31/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI11/MM2 N_XI31/XI11/NET34_XI31/XI11/MM2_d
+ N_XI31/XI11/NET33_XI31/XI11/MM2_g N_VSS_XI31/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI11/MM3 N_XI31/XI11/NET33_XI31/XI11/MM3_d N_WL<58>_XI31/XI11/MM3_g
+ N_BLN<4>_XI31/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI11/MM0 N_XI31/XI11/NET34_XI31/XI11/MM0_d N_WL<58>_XI31/XI11/MM0_g
+ N_BL<4>_XI31/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI11/MM1 N_XI31/XI11/NET33_XI31/XI11/MM1_d
+ N_XI31/XI11/NET34_XI31/XI11/MM1_g N_VSS_XI31/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI11/MM9 N_XI31/XI11/NET36_XI31/XI11/MM9_d N_WL<59>_XI31/XI11/MM9_g
+ N_BL<4>_XI31/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI11/MM6 N_XI31/XI11/NET35_XI31/XI11/MM6_d
+ N_XI31/XI11/NET36_XI31/XI11/MM6_g N_VSS_XI31/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI11/MM7 N_XI31/XI11/NET36_XI31/XI11/MM7_d
+ N_XI31/XI11/NET35_XI31/XI11/MM7_g N_VSS_XI31/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI11/MM8 N_XI31/XI11/NET35_XI31/XI11/MM8_d N_WL<59>_XI31/XI11/MM8_g
+ N_BLN<4>_XI31/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI11/MM5 N_XI31/XI11/NET34_XI31/XI11/MM5_d
+ N_XI31/XI11/NET33_XI31/XI11/MM5_g N_VDD_XI31/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI11/MM4 N_XI31/XI11/NET33_XI31/XI11/MM4_d
+ N_XI31/XI11/NET34_XI31/XI11/MM4_g N_VDD_XI31/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI11/MM10 N_XI31/XI11/NET35_XI31/XI11/MM10_d
+ N_XI31/XI11/NET36_XI31/XI11/MM10_g N_VDD_XI31/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI11/MM11 N_XI31/XI11/NET36_XI31/XI11/MM11_d
+ N_XI31/XI11/NET35_XI31/XI11/MM11_g N_VDD_XI31/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI12/MM2 N_XI31/XI12/NET34_XI31/XI12/MM2_d
+ N_XI31/XI12/NET33_XI31/XI12/MM2_g N_VSS_XI31/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI12/MM3 N_XI31/XI12/NET33_XI31/XI12/MM3_d N_WL<58>_XI31/XI12/MM3_g
+ N_BLN<3>_XI31/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI12/MM0 N_XI31/XI12/NET34_XI31/XI12/MM0_d N_WL<58>_XI31/XI12/MM0_g
+ N_BL<3>_XI31/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI12/MM1 N_XI31/XI12/NET33_XI31/XI12/MM1_d
+ N_XI31/XI12/NET34_XI31/XI12/MM1_g N_VSS_XI31/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI12/MM9 N_XI31/XI12/NET36_XI31/XI12/MM9_d N_WL<59>_XI31/XI12/MM9_g
+ N_BL<3>_XI31/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI12/MM6 N_XI31/XI12/NET35_XI31/XI12/MM6_d
+ N_XI31/XI12/NET36_XI31/XI12/MM6_g N_VSS_XI31/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI12/MM7 N_XI31/XI12/NET36_XI31/XI12/MM7_d
+ N_XI31/XI12/NET35_XI31/XI12/MM7_g N_VSS_XI31/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI12/MM8 N_XI31/XI12/NET35_XI31/XI12/MM8_d N_WL<59>_XI31/XI12/MM8_g
+ N_BLN<3>_XI31/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI12/MM5 N_XI31/XI12/NET34_XI31/XI12/MM5_d
+ N_XI31/XI12/NET33_XI31/XI12/MM5_g N_VDD_XI31/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI12/MM4 N_XI31/XI12/NET33_XI31/XI12/MM4_d
+ N_XI31/XI12/NET34_XI31/XI12/MM4_g N_VDD_XI31/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI12/MM10 N_XI31/XI12/NET35_XI31/XI12/MM10_d
+ N_XI31/XI12/NET36_XI31/XI12/MM10_g N_VDD_XI31/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI12/MM11 N_XI31/XI12/NET36_XI31/XI12/MM11_d
+ N_XI31/XI12/NET35_XI31/XI12/MM11_g N_VDD_XI31/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI13/MM2 N_XI31/XI13/NET34_XI31/XI13/MM2_d
+ N_XI31/XI13/NET33_XI31/XI13/MM2_g N_VSS_XI31/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI13/MM3 N_XI31/XI13/NET33_XI31/XI13/MM3_d N_WL<58>_XI31/XI13/MM3_g
+ N_BLN<2>_XI31/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI13/MM0 N_XI31/XI13/NET34_XI31/XI13/MM0_d N_WL<58>_XI31/XI13/MM0_g
+ N_BL<2>_XI31/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI13/MM1 N_XI31/XI13/NET33_XI31/XI13/MM1_d
+ N_XI31/XI13/NET34_XI31/XI13/MM1_g N_VSS_XI31/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI13/MM9 N_XI31/XI13/NET36_XI31/XI13/MM9_d N_WL<59>_XI31/XI13/MM9_g
+ N_BL<2>_XI31/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI13/MM6 N_XI31/XI13/NET35_XI31/XI13/MM6_d
+ N_XI31/XI13/NET36_XI31/XI13/MM6_g N_VSS_XI31/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI13/MM7 N_XI31/XI13/NET36_XI31/XI13/MM7_d
+ N_XI31/XI13/NET35_XI31/XI13/MM7_g N_VSS_XI31/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI13/MM8 N_XI31/XI13/NET35_XI31/XI13/MM8_d N_WL<59>_XI31/XI13/MM8_g
+ N_BLN<2>_XI31/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI13/MM5 N_XI31/XI13/NET34_XI31/XI13/MM5_d
+ N_XI31/XI13/NET33_XI31/XI13/MM5_g N_VDD_XI31/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI13/MM4 N_XI31/XI13/NET33_XI31/XI13/MM4_d
+ N_XI31/XI13/NET34_XI31/XI13/MM4_g N_VDD_XI31/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI13/MM10 N_XI31/XI13/NET35_XI31/XI13/MM10_d
+ N_XI31/XI13/NET36_XI31/XI13/MM10_g N_VDD_XI31/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI13/MM11 N_XI31/XI13/NET36_XI31/XI13/MM11_d
+ N_XI31/XI13/NET35_XI31/XI13/MM11_g N_VDD_XI31/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI14/MM2 N_XI31/XI14/NET34_XI31/XI14/MM2_d
+ N_XI31/XI14/NET33_XI31/XI14/MM2_g N_VSS_XI31/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI14/MM3 N_XI31/XI14/NET33_XI31/XI14/MM3_d N_WL<58>_XI31/XI14/MM3_g
+ N_BLN<1>_XI31/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI14/MM0 N_XI31/XI14/NET34_XI31/XI14/MM0_d N_WL<58>_XI31/XI14/MM0_g
+ N_BL<1>_XI31/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI14/MM1 N_XI31/XI14/NET33_XI31/XI14/MM1_d
+ N_XI31/XI14/NET34_XI31/XI14/MM1_g N_VSS_XI31/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI14/MM9 N_XI31/XI14/NET36_XI31/XI14/MM9_d N_WL<59>_XI31/XI14/MM9_g
+ N_BL<1>_XI31/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI14/MM6 N_XI31/XI14/NET35_XI31/XI14/MM6_d
+ N_XI31/XI14/NET36_XI31/XI14/MM6_g N_VSS_XI31/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI14/MM7 N_XI31/XI14/NET36_XI31/XI14/MM7_d
+ N_XI31/XI14/NET35_XI31/XI14/MM7_g N_VSS_XI31/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI14/MM8 N_XI31/XI14/NET35_XI31/XI14/MM8_d N_WL<59>_XI31/XI14/MM8_g
+ N_BLN<1>_XI31/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI14/MM5 N_XI31/XI14/NET34_XI31/XI14/MM5_d
+ N_XI31/XI14/NET33_XI31/XI14/MM5_g N_VDD_XI31/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI14/MM4 N_XI31/XI14/NET33_XI31/XI14/MM4_d
+ N_XI31/XI14/NET34_XI31/XI14/MM4_g N_VDD_XI31/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI14/MM10 N_XI31/XI14/NET35_XI31/XI14/MM10_d
+ N_XI31/XI14/NET36_XI31/XI14/MM10_g N_VDD_XI31/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI14/MM11 N_XI31/XI14/NET36_XI31/XI14/MM11_d
+ N_XI31/XI14/NET35_XI31/XI14/MM11_g N_VDD_XI31/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI15/MM2 N_XI31/XI15/NET34_XI31/XI15/MM2_d
+ N_XI31/XI15/NET33_XI31/XI15/MM2_g N_VSS_XI31/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI15/MM3 N_XI31/XI15/NET33_XI31/XI15/MM3_d N_WL<58>_XI31/XI15/MM3_g
+ N_BLN<0>_XI31/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI15/MM0 N_XI31/XI15/NET34_XI31/XI15/MM0_d N_WL<58>_XI31/XI15/MM0_g
+ N_BL<0>_XI31/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI15/MM1 N_XI31/XI15/NET33_XI31/XI15/MM1_d
+ N_XI31/XI15/NET34_XI31/XI15/MM1_g N_VSS_XI31/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI15/MM9 N_XI31/XI15/NET36_XI31/XI15/MM9_d N_WL<59>_XI31/XI15/MM9_g
+ N_BL<0>_XI31/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI15/MM6 N_XI31/XI15/NET35_XI31/XI15/MM6_d
+ N_XI31/XI15/NET36_XI31/XI15/MM6_g N_VSS_XI31/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI15/MM7 N_XI31/XI15/NET36_XI31/XI15/MM7_d
+ N_XI31/XI15/NET35_XI31/XI15/MM7_g N_VSS_XI31/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI31/XI15/MM8 N_XI31/XI15/NET35_XI31/XI15/MM8_d N_WL<59>_XI31/XI15/MM8_g
+ N_BLN<0>_XI31/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI31/XI15/MM5 N_XI31/XI15/NET34_XI31/XI15/MM5_d
+ N_XI31/XI15/NET33_XI31/XI15/MM5_g N_VDD_XI31/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI15/MM4 N_XI31/XI15/NET33_XI31/XI15/MM4_d
+ N_XI31/XI15/NET34_XI31/XI15/MM4_g N_VDD_XI31/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI15/MM10 N_XI31/XI15/NET35_XI31/XI15/MM10_d
+ N_XI31/XI15/NET36_XI31/XI15/MM10_g N_VDD_XI31/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI31/XI15/MM11 N_XI31/XI15/NET36_XI31/XI15/MM11_d
+ N_XI31/XI15/NET35_XI31/XI15/MM11_g N_VDD_XI31/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI0/MM2 N_XI32/XI0/NET34_XI32/XI0/MM2_d N_XI32/XI0/NET33_XI32/XI0/MM2_g
+ N_VSS_XI32/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI0/MM3 N_XI32/XI0/NET33_XI32/XI0/MM3_d N_WL<60>_XI32/XI0/MM3_g
+ N_BLN<15>_XI32/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI0/MM0 N_XI32/XI0/NET34_XI32/XI0/MM0_d N_WL<60>_XI32/XI0/MM0_g
+ N_BL<15>_XI32/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI0/MM1 N_XI32/XI0/NET33_XI32/XI0/MM1_d N_XI32/XI0/NET34_XI32/XI0/MM1_g
+ N_VSS_XI32/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI0/MM9 N_XI32/XI0/NET36_XI32/XI0/MM9_d N_WL<61>_XI32/XI0/MM9_g
+ N_BL<15>_XI32/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI0/MM6 N_XI32/XI0/NET35_XI32/XI0/MM6_d N_XI32/XI0/NET36_XI32/XI0/MM6_g
+ N_VSS_XI32/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI0/MM7 N_XI32/XI0/NET36_XI32/XI0/MM7_d N_XI32/XI0/NET35_XI32/XI0/MM7_g
+ N_VSS_XI32/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI0/MM8 N_XI32/XI0/NET35_XI32/XI0/MM8_d N_WL<61>_XI32/XI0/MM8_g
+ N_BLN<15>_XI32/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI0/MM5 N_XI32/XI0/NET34_XI32/XI0/MM5_d N_XI32/XI0/NET33_XI32/XI0/MM5_g
+ N_VDD_XI32/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI0/MM4 N_XI32/XI0/NET33_XI32/XI0/MM4_d N_XI32/XI0/NET34_XI32/XI0/MM4_g
+ N_VDD_XI32/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI0/MM10 N_XI32/XI0/NET35_XI32/XI0/MM10_d N_XI32/XI0/NET36_XI32/XI0/MM10_g
+ N_VDD_XI32/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI0/MM11 N_XI32/XI0/NET36_XI32/XI0/MM11_d N_XI32/XI0/NET35_XI32/XI0/MM11_g
+ N_VDD_XI32/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI1/MM2 N_XI32/XI1/NET34_XI32/XI1/MM2_d N_XI32/XI1/NET33_XI32/XI1/MM2_g
+ N_VSS_XI32/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI1/MM3 N_XI32/XI1/NET33_XI32/XI1/MM3_d N_WL<60>_XI32/XI1/MM3_g
+ N_BLN<14>_XI32/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI1/MM0 N_XI32/XI1/NET34_XI32/XI1/MM0_d N_WL<60>_XI32/XI1/MM0_g
+ N_BL<14>_XI32/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI1/MM1 N_XI32/XI1/NET33_XI32/XI1/MM1_d N_XI32/XI1/NET34_XI32/XI1/MM1_g
+ N_VSS_XI32/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI1/MM9 N_XI32/XI1/NET36_XI32/XI1/MM9_d N_WL<61>_XI32/XI1/MM9_g
+ N_BL<14>_XI32/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI1/MM6 N_XI32/XI1/NET35_XI32/XI1/MM6_d N_XI32/XI1/NET36_XI32/XI1/MM6_g
+ N_VSS_XI32/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI1/MM7 N_XI32/XI1/NET36_XI32/XI1/MM7_d N_XI32/XI1/NET35_XI32/XI1/MM7_g
+ N_VSS_XI32/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI1/MM8 N_XI32/XI1/NET35_XI32/XI1/MM8_d N_WL<61>_XI32/XI1/MM8_g
+ N_BLN<14>_XI32/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI1/MM5 N_XI32/XI1/NET34_XI32/XI1/MM5_d N_XI32/XI1/NET33_XI32/XI1/MM5_g
+ N_VDD_XI32/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI1/MM4 N_XI32/XI1/NET33_XI32/XI1/MM4_d N_XI32/XI1/NET34_XI32/XI1/MM4_g
+ N_VDD_XI32/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI1/MM10 N_XI32/XI1/NET35_XI32/XI1/MM10_d N_XI32/XI1/NET36_XI32/XI1/MM10_g
+ N_VDD_XI32/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI1/MM11 N_XI32/XI1/NET36_XI32/XI1/MM11_d N_XI32/XI1/NET35_XI32/XI1/MM11_g
+ N_VDD_XI32/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI2/MM2 N_XI32/XI2/NET34_XI32/XI2/MM2_d N_XI32/XI2/NET33_XI32/XI2/MM2_g
+ N_VSS_XI32/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI2/MM3 N_XI32/XI2/NET33_XI32/XI2/MM3_d N_WL<60>_XI32/XI2/MM3_g
+ N_BLN<13>_XI32/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI2/MM0 N_XI32/XI2/NET34_XI32/XI2/MM0_d N_WL<60>_XI32/XI2/MM0_g
+ N_BL<13>_XI32/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI2/MM1 N_XI32/XI2/NET33_XI32/XI2/MM1_d N_XI32/XI2/NET34_XI32/XI2/MM1_g
+ N_VSS_XI32/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI2/MM9 N_XI32/XI2/NET36_XI32/XI2/MM9_d N_WL<61>_XI32/XI2/MM9_g
+ N_BL<13>_XI32/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI2/MM6 N_XI32/XI2/NET35_XI32/XI2/MM6_d N_XI32/XI2/NET36_XI32/XI2/MM6_g
+ N_VSS_XI32/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI2/MM7 N_XI32/XI2/NET36_XI32/XI2/MM7_d N_XI32/XI2/NET35_XI32/XI2/MM7_g
+ N_VSS_XI32/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI2/MM8 N_XI32/XI2/NET35_XI32/XI2/MM8_d N_WL<61>_XI32/XI2/MM8_g
+ N_BLN<13>_XI32/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI2/MM5 N_XI32/XI2/NET34_XI32/XI2/MM5_d N_XI32/XI2/NET33_XI32/XI2/MM5_g
+ N_VDD_XI32/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI2/MM4 N_XI32/XI2/NET33_XI32/XI2/MM4_d N_XI32/XI2/NET34_XI32/XI2/MM4_g
+ N_VDD_XI32/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI2/MM10 N_XI32/XI2/NET35_XI32/XI2/MM10_d N_XI32/XI2/NET36_XI32/XI2/MM10_g
+ N_VDD_XI32/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI2/MM11 N_XI32/XI2/NET36_XI32/XI2/MM11_d N_XI32/XI2/NET35_XI32/XI2/MM11_g
+ N_VDD_XI32/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI3/MM2 N_XI32/XI3/NET34_XI32/XI3/MM2_d N_XI32/XI3/NET33_XI32/XI3/MM2_g
+ N_VSS_XI32/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI3/MM3 N_XI32/XI3/NET33_XI32/XI3/MM3_d N_WL<60>_XI32/XI3/MM3_g
+ N_BLN<12>_XI32/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI3/MM0 N_XI32/XI3/NET34_XI32/XI3/MM0_d N_WL<60>_XI32/XI3/MM0_g
+ N_BL<12>_XI32/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI3/MM1 N_XI32/XI3/NET33_XI32/XI3/MM1_d N_XI32/XI3/NET34_XI32/XI3/MM1_g
+ N_VSS_XI32/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI3/MM9 N_XI32/XI3/NET36_XI32/XI3/MM9_d N_WL<61>_XI32/XI3/MM9_g
+ N_BL<12>_XI32/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI3/MM6 N_XI32/XI3/NET35_XI32/XI3/MM6_d N_XI32/XI3/NET36_XI32/XI3/MM6_g
+ N_VSS_XI32/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI3/MM7 N_XI32/XI3/NET36_XI32/XI3/MM7_d N_XI32/XI3/NET35_XI32/XI3/MM7_g
+ N_VSS_XI32/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI3/MM8 N_XI32/XI3/NET35_XI32/XI3/MM8_d N_WL<61>_XI32/XI3/MM8_g
+ N_BLN<12>_XI32/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI3/MM5 N_XI32/XI3/NET34_XI32/XI3/MM5_d N_XI32/XI3/NET33_XI32/XI3/MM5_g
+ N_VDD_XI32/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI3/MM4 N_XI32/XI3/NET33_XI32/XI3/MM4_d N_XI32/XI3/NET34_XI32/XI3/MM4_g
+ N_VDD_XI32/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI3/MM10 N_XI32/XI3/NET35_XI32/XI3/MM10_d N_XI32/XI3/NET36_XI32/XI3/MM10_g
+ N_VDD_XI32/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI3/MM11 N_XI32/XI3/NET36_XI32/XI3/MM11_d N_XI32/XI3/NET35_XI32/XI3/MM11_g
+ N_VDD_XI32/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI4/MM2 N_XI32/XI4/NET34_XI32/XI4/MM2_d N_XI32/XI4/NET33_XI32/XI4/MM2_g
+ N_VSS_XI32/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI4/MM3 N_XI32/XI4/NET33_XI32/XI4/MM3_d N_WL<60>_XI32/XI4/MM3_g
+ N_BLN<11>_XI32/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI4/MM0 N_XI32/XI4/NET34_XI32/XI4/MM0_d N_WL<60>_XI32/XI4/MM0_g
+ N_BL<11>_XI32/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI4/MM1 N_XI32/XI4/NET33_XI32/XI4/MM1_d N_XI32/XI4/NET34_XI32/XI4/MM1_g
+ N_VSS_XI32/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI4/MM9 N_XI32/XI4/NET36_XI32/XI4/MM9_d N_WL<61>_XI32/XI4/MM9_g
+ N_BL<11>_XI32/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI4/MM6 N_XI32/XI4/NET35_XI32/XI4/MM6_d N_XI32/XI4/NET36_XI32/XI4/MM6_g
+ N_VSS_XI32/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI4/MM7 N_XI32/XI4/NET36_XI32/XI4/MM7_d N_XI32/XI4/NET35_XI32/XI4/MM7_g
+ N_VSS_XI32/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI4/MM8 N_XI32/XI4/NET35_XI32/XI4/MM8_d N_WL<61>_XI32/XI4/MM8_g
+ N_BLN<11>_XI32/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI4/MM5 N_XI32/XI4/NET34_XI32/XI4/MM5_d N_XI32/XI4/NET33_XI32/XI4/MM5_g
+ N_VDD_XI32/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI4/MM4 N_XI32/XI4/NET33_XI32/XI4/MM4_d N_XI32/XI4/NET34_XI32/XI4/MM4_g
+ N_VDD_XI32/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI4/MM10 N_XI32/XI4/NET35_XI32/XI4/MM10_d N_XI32/XI4/NET36_XI32/XI4/MM10_g
+ N_VDD_XI32/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI4/MM11 N_XI32/XI4/NET36_XI32/XI4/MM11_d N_XI32/XI4/NET35_XI32/XI4/MM11_g
+ N_VDD_XI32/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI5/MM2 N_XI32/XI5/NET34_XI32/XI5/MM2_d N_XI32/XI5/NET33_XI32/XI5/MM2_g
+ N_VSS_XI32/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI5/MM3 N_XI32/XI5/NET33_XI32/XI5/MM3_d N_WL<60>_XI32/XI5/MM3_g
+ N_BLN<10>_XI32/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI5/MM0 N_XI32/XI5/NET34_XI32/XI5/MM0_d N_WL<60>_XI32/XI5/MM0_g
+ N_BL<10>_XI32/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI5/MM1 N_XI32/XI5/NET33_XI32/XI5/MM1_d N_XI32/XI5/NET34_XI32/XI5/MM1_g
+ N_VSS_XI32/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI5/MM9 N_XI32/XI5/NET36_XI32/XI5/MM9_d N_WL<61>_XI32/XI5/MM9_g
+ N_BL<10>_XI32/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI5/MM6 N_XI32/XI5/NET35_XI32/XI5/MM6_d N_XI32/XI5/NET36_XI32/XI5/MM6_g
+ N_VSS_XI32/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI5/MM7 N_XI32/XI5/NET36_XI32/XI5/MM7_d N_XI32/XI5/NET35_XI32/XI5/MM7_g
+ N_VSS_XI32/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI5/MM8 N_XI32/XI5/NET35_XI32/XI5/MM8_d N_WL<61>_XI32/XI5/MM8_g
+ N_BLN<10>_XI32/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI5/MM5 N_XI32/XI5/NET34_XI32/XI5/MM5_d N_XI32/XI5/NET33_XI32/XI5/MM5_g
+ N_VDD_XI32/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI5/MM4 N_XI32/XI5/NET33_XI32/XI5/MM4_d N_XI32/XI5/NET34_XI32/XI5/MM4_g
+ N_VDD_XI32/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI5/MM10 N_XI32/XI5/NET35_XI32/XI5/MM10_d N_XI32/XI5/NET36_XI32/XI5/MM10_g
+ N_VDD_XI32/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI5/MM11 N_XI32/XI5/NET36_XI32/XI5/MM11_d N_XI32/XI5/NET35_XI32/XI5/MM11_g
+ N_VDD_XI32/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI6/MM2 N_XI32/XI6/NET34_XI32/XI6/MM2_d N_XI32/XI6/NET33_XI32/XI6/MM2_g
+ N_VSS_XI32/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM3 N_XI32/XI6/NET33_XI32/XI6/MM3_d N_WL<60>_XI32/XI6/MM3_g
+ N_BLN<9>_XI32/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM0 N_XI32/XI6/NET34_XI32/XI6/MM0_d N_WL<60>_XI32/XI6/MM0_g
+ N_BL<9>_XI32/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM1 N_XI32/XI6/NET33_XI32/XI6/MM1_d N_XI32/XI6/NET34_XI32/XI6/MM1_g
+ N_VSS_XI32/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM9 N_XI32/XI6/NET36_XI32/XI6/MM9_d N_WL<61>_XI32/XI6/MM9_g
+ N_BL<9>_XI32/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM6 N_XI32/XI6/NET35_XI32/XI6/MM6_d N_XI32/XI6/NET36_XI32/XI6/MM6_g
+ N_VSS_XI32/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM7 N_XI32/XI6/NET36_XI32/XI6/MM7_d N_XI32/XI6/NET35_XI32/XI6/MM7_g
+ N_VSS_XI32/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM8 N_XI32/XI6/NET35_XI32/XI6/MM8_d N_WL<61>_XI32/XI6/MM8_g
+ N_BLN<9>_XI32/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI6/MM5 N_XI32/XI6/NET34_XI32/XI6/MM5_d N_XI32/XI6/NET33_XI32/XI6/MM5_g
+ N_VDD_XI32/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI6/MM4 N_XI32/XI6/NET33_XI32/XI6/MM4_d N_XI32/XI6/NET34_XI32/XI6/MM4_g
+ N_VDD_XI32/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI6/MM10 N_XI32/XI6/NET35_XI32/XI6/MM10_d N_XI32/XI6/NET36_XI32/XI6/MM10_g
+ N_VDD_XI32/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI6/MM11 N_XI32/XI6/NET36_XI32/XI6/MM11_d N_XI32/XI6/NET35_XI32/XI6/MM11_g
+ N_VDD_XI32/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI7/MM2 N_XI32/XI7/NET34_XI32/XI7/MM2_d N_XI32/XI7/NET33_XI32/XI7/MM2_g
+ N_VSS_XI32/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM3 N_XI32/XI7/NET33_XI32/XI7/MM3_d N_WL<60>_XI32/XI7/MM3_g
+ N_BLN<8>_XI32/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM0 N_XI32/XI7/NET34_XI32/XI7/MM0_d N_WL<60>_XI32/XI7/MM0_g
+ N_BL<8>_XI32/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM1 N_XI32/XI7/NET33_XI32/XI7/MM1_d N_XI32/XI7/NET34_XI32/XI7/MM1_g
+ N_VSS_XI32/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM9 N_XI32/XI7/NET36_XI32/XI7/MM9_d N_WL<61>_XI32/XI7/MM9_g
+ N_BL<8>_XI32/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM6 N_XI32/XI7/NET35_XI32/XI7/MM6_d N_XI32/XI7/NET36_XI32/XI7/MM6_g
+ N_VSS_XI32/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM7 N_XI32/XI7/NET36_XI32/XI7/MM7_d N_XI32/XI7/NET35_XI32/XI7/MM7_g
+ N_VSS_XI32/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM8 N_XI32/XI7/NET35_XI32/XI7/MM8_d N_WL<61>_XI32/XI7/MM8_g
+ N_BLN<8>_XI32/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI7/MM5 N_XI32/XI7/NET34_XI32/XI7/MM5_d N_XI32/XI7/NET33_XI32/XI7/MM5_g
+ N_VDD_XI32/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI7/MM4 N_XI32/XI7/NET33_XI32/XI7/MM4_d N_XI32/XI7/NET34_XI32/XI7/MM4_g
+ N_VDD_XI32/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI7/MM10 N_XI32/XI7/NET35_XI32/XI7/MM10_d N_XI32/XI7/NET36_XI32/XI7/MM10_g
+ N_VDD_XI32/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI7/MM11 N_XI32/XI7/NET36_XI32/XI7/MM11_d N_XI32/XI7/NET35_XI32/XI7/MM11_g
+ N_VDD_XI32/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI8/MM2 N_XI32/XI8/NET34_XI32/XI8/MM2_d N_XI32/XI8/NET33_XI32/XI8/MM2_g
+ N_VSS_XI32/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM3 N_XI32/XI8/NET33_XI32/XI8/MM3_d N_WL<60>_XI32/XI8/MM3_g
+ N_BLN<7>_XI32/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM0 N_XI32/XI8/NET34_XI32/XI8/MM0_d N_WL<60>_XI32/XI8/MM0_g
+ N_BL<7>_XI32/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM1 N_XI32/XI8/NET33_XI32/XI8/MM1_d N_XI32/XI8/NET34_XI32/XI8/MM1_g
+ N_VSS_XI32/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM9 N_XI32/XI8/NET36_XI32/XI8/MM9_d N_WL<61>_XI32/XI8/MM9_g
+ N_BL<7>_XI32/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM6 N_XI32/XI8/NET35_XI32/XI8/MM6_d N_XI32/XI8/NET36_XI32/XI8/MM6_g
+ N_VSS_XI32/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM7 N_XI32/XI8/NET36_XI32/XI8/MM7_d N_XI32/XI8/NET35_XI32/XI8/MM7_g
+ N_VSS_XI32/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM8 N_XI32/XI8/NET35_XI32/XI8/MM8_d N_WL<61>_XI32/XI8/MM8_g
+ N_BLN<7>_XI32/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI8/MM5 N_XI32/XI8/NET34_XI32/XI8/MM5_d N_XI32/XI8/NET33_XI32/XI8/MM5_g
+ N_VDD_XI32/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI8/MM4 N_XI32/XI8/NET33_XI32/XI8/MM4_d N_XI32/XI8/NET34_XI32/XI8/MM4_g
+ N_VDD_XI32/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI8/MM10 N_XI32/XI8/NET35_XI32/XI8/MM10_d N_XI32/XI8/NET36_XI32/XI8/MM10_g
+ N_VDD_XI32/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI8/MM11 N_XI32/XI8/NET36_XI32/XI8/MM11_d N_XI32/XI8/NET35_XI32/XI8/MM11_g
+ N_VDD_XI32/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI9/MM2 N_XI32/XI9/NET34_XI32/XI9/MM2_d N_XI32/XI9/NET33_XI32/XI9/MM2_g
+ N_VSS_XI32/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM3 N_XI32/XI9/NET33_XI32/XI9/MM3_d N_WL<60>_XI32/XI9/MM3_g
+ N_BLN<6>_XI32/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM0 N_XI32/XI9/NET34_XI32/XI9/MM0_d N_WL<60>_XI32/XI9/MM0_g
+ N_BL<6>_XI32/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM1 N_XI32/XI9/NET33_XI32/XI9/MM1_d N_XI32/XI9/NET34_XI32/XI9/MM1_g
+ N_VSS_XI32/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM9 N_XI32/XI9/NET36_XI32/XI9/MM9_d N_WL<61>_XI32/XI9/MM9_g
+ N_BL<6>_XI32/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM6 N_XI32/XI9/NET35_XI32/XI9/MM6_d N_XI32/XI9/NET36_XI32/XI9/MM6_g
+ N_VSS_XI32/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM7 N_XI32/XI9/NET36_XI32/XI9/MM7_d N_XI32/XI9/NET35_XI32/XI9/MM7_g
+ N_VSS_XI32/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM8 N_XI32/XI9/NET35_XI32/XI9/MM8_d N_WL<61>_XI32/XI9/MM8_g
+ N_BLN<6>_XI32/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI9/MM5 N_XI32/XI9/NET34_XI32/XI9/MM5_d N_XI32/XI9/NET33_XI32/XI9/MM5_g
+ N_VDD_XI32/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI9/MM4 N_XI32/XI9/NET33_XI32/XI9/MM4_d N_XI32/XI9/NET34_XI32/XI9/MM4_g
+ N_VDD_XI32/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI9/MM10 N_XI32/XI9/NET35_XI32/XI9/MM10_d N_XI32/XI9/NET36_XI32/XI9/MM10_g
+ N_VDD_XI32/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI9/MM11 N_XI32/XI9/NET36_XI32/XI9/MM11_d N_XI32/XI9/NET35_XI32/XI9/MM11_g
+ N_VDD_XI32/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI10/MM2 N_XI32/XI10/NET34_XI32/XI10/MM2_d
+ N_XI32/XI10/NET33_XI32/XI10/MM2_g N_VSS_XI32/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI10/MM3 N_XI32/XI10/NET33_XI32/XI10/MM3_d N_WL<60>_XI32/XI10/MM3_g
+ N_BLN<5>_XI32/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI10/MM0 N_XI32/XI10/NET34_XI32/XI10/MM0_d N_WL<60>_XI32/XI10/MM0_g
+ N_BL<5>_XI32/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI10/MM1 N_XI32/XI10/NET33_XI32/XI10/MM1_d
+ N_XI32/XI10/NET34_XI32/XI10/MM1_g N_VSS_XI32/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI10/MM9 N_XI32/XI10/NET36_XI32/XI10/MM9_d N_WL<61>_XI32/XI10/MM9_g
+ N_BL<5>_XI32/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI10/MM6 N_XI32/XI10/NET35_XI32/XI10/MM6_d
+ N_XI32/XI10/NET36_XI32/XI10/MM6_g N_VSS_XI32/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI10/MM7 N_XI32/XI10/NET36_XI32/XI10/MM7_d
+ N_XI32/XI10/NET35_XI32/XI10/MM7_g N_VSS_XI32/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI10/MM8 N_XI32/XI10/NET35_XI32/XI10/MM8_d N_WL<61>_XI32/XI10/MM8_g
+ N_BLN<5>_XI32/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI10/MM5 N_XI32/XI10/NET34_XI32/XI10/MM5_d
+ N_XI32/XI10/NET33_XI32/XI10/MM5_g N_VDD_XI32/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI10/MM4 N_XI32/XI10/NET33_XI32/XI10/MM4_d
+ N_XI32/XI10/NET34_XI32/XI10/MM4_g N_VDD_XI32/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI10/MM10 N_XI32/XI10/NET35_XI32/XI10/MM10_d
+ N_XI32/XI10/NET36_XI32/XI10/MM10_g N_VDD_XI32/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI10/MM11 N_XI32/XI10/NET36_XI32/XI10/MM11_d
+ N_XI32/XI10/NET35_XI32/XI10/MM11_g N_VDD_XI32/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI11/MM2 N_XI32/XI11/NET34_XI32/XI11/MM2_d
+ N_XI32/XI11/NET33_XI32/XI11/MM2_g N_VSS_XI32/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI11/MM3 N_XI32/XI11/NET33_XI32/XI11/MM3_d N_WL<60>_XI32/XI11/MM3_g
+ N_BLN<4>_XI32/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI11/MM0 N_XI32/XI11/NET34_XI32/XI11/MM0_d N_WL<60>_XI32/XI11/MM0_g
+ N_BL<4>_XI32/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI11/MM1 N_XI32/XI11/NET33_XI32/XI11/MM1_d
+ N_XI32/XI11/NET34_XI32/XI11/MM1_g N_VSS_XI32/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI11/MM9 N_XI32/XI11/NET36_XI32/XI11/MM9_d N_WL<61>_XI32/XI11/MM9_g
+ N_BL<4>_XI32/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI11/MM6 N_XI32/XI11/NET35_XI32/XI11/MM6_d
+ N_XI32/XI11/NET36_XI32/XI11/MM6_g N_VSS_XI32/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI11/MM7 N_XI32/XI11/NET36_XI32/XI11/MM7_d
+ N_XI32/XI11/NET35_XI32/XI11/MM7_g N_VSS_XI32/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI11/MM8 N_XI32/XI11/NET35_XI32/XI11/MM8_d N_WL<61>_XI32/XI11/MM8_g
+ N_BLN<4>_XI32/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI11/MM5 N_XI32/XI11/NET34_XI32/XI11/MM5_d
+ N_XI32/XI11/NET33_XI32/XI11/MM5_g N_VDD_XI32/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI11/MM4 N_XI32/XI11/NET33_XI32/XI11/MM4_d
+ N_XI32/XI11/NET34_XI32/XI11/MM4_g N_VDD_XI32/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI11/MM10 N_XI32/XI11/NET35_XI32/XI11/MM10_d
+ N_XI32/XI11/NET36_XI32/XI11/MM10_g N_VDD_XI32/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI11/MM11 N_XI32/XI11/NET36_XI32/XI11/MM11_d
+ N_XI32/XI11/NET35_XI32/XI11/MM11_g N_VDD_XI32/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI12/MM2 N_XI32/XI12/NET34_XI32/XI12/MM2_d
+ N_XI32/XI12/NET33_XI32/XI12/MM2_g N_VSS_XI32/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI12/MM3 N_XI32/XI12/NET33_XI32/XI12/MM3_d N_WL<60>_XI32/XI12/MM3_g
+ N_BLN<3>_XI32/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI12/MM0 N_XI32/XI12/NET34_XI32/XI12/MM0_d N_WL<60>_XI32/XI12/MM0_g
+ N_BL<3>_XI32/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI12/MM1 N_XI32/XI12/NET33_XI32/XI12/MM1_d
+ N_XI32/XI12/NET34_XI32/XI12/MM1_g N_VSS_XI32/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI12/MM9 N_XI32/XI12/NET36_XI32/XI12/MM9_d N_WL<61>_XI32/XI12/MM9_g
+ N_BL<3>_XI32/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI12/MM6 N_XI32/XI12/NET35_XI32/XI12/MM6_d
+ N_XI32/XI12/NET36_XI32/XI12/MM6_g N_VSS_XI32/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI12/MM7 N_XI32/XI12/NET36_XI32/XI12/MM7_d
+ N_XI32/XI12/NET35_XI32/XI12/MM7_g N_VSS_XI32/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI12/MM8 N_XI32/XI12/NET35_XI32/XI12/MM8_d N_WL<61>_XI32/XI12/MM8_g
+ N_BLN<3>_XI32/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI12/MM5 N_XI32/XI12/NET34_XI32/XI12/MM5_d
+ N_XI32/XI12/NET33_XI32/XI12/MM5_g N_VDD_XI32/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI12/MM4 N_XI32/XI12/NET33_XI32/XI12/MM4_d
+ N_XI32/XI12/NET34_XI32/XI12/MM4_g N_VDD_XI32/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI12/MM10 N_XI32/XI12/NET35_XI32/XI12/MM10_d
+ N_XI32/XI12/NET36_XI32/XI12/MM10_g N_VDD_XI32/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI12/MM11 N_XI32/XI12/NET36_XI32/XI12/MM11_d
+ N_XI32/XI12/NET35_XI32/XI12/MM11_g N_VDD_XI32/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI13/MM2 N_XI32/XI13/NET34_XI32/XI13/MM2_d
+ N_XI32/XI13/NET33_XI32/XI13/MM2_g N_VSS_XI32/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI13/MM3 N_XI32/XI13/NET33_XI32/XI13/MM3_d N_WL<60>_XI32/XI13/MM3_g
+ N_BLN<2>_XI32/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI13/MM0 N_XI32/XI13/NET34_XI32/XI13/MM0_d N_WL<60>_XI32/XI13/MM0_g
+ N_BL<2>_XI32/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI13/MM1 N_XI32/XI13/NET33_XI32/XI13/MM1_d
+ N_XI32/XI13/NET34_XI32/XI13/MM1_g N_VSS_XI32/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI13/MM9 N_XI32/XI13/NET36_XI32/XI13/MM9_d N_WL<61>_XI32/XI13/MM9_g
+ N_BL<2>_XI32/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI13/MM6 N_XI32/XI13/NET35_XI32/XI13/MM6_d
+ N_XI32/XI13/NET36_XI32/XI13/MM6_g N_VSS_XI32/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI13/MM7 N_XI32/XI13/NET36_XI32/XI13/MM7_d
+ N_XI32/XI13/NET35_XI32/XI13/MM7_g N_VSS_XI32/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI13/MM8 N_XI32/XI13/NET35_XI32/XI13/MM8_d N_WL<61>_XI32/XI13/MM8_g
+ N_BLN<2>_XI32/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI13/MM5 N_XI32/XI13/NET34_XI32/XI13/MM5_d
+ N_XI32/XI13/NET33_XI32/XI13/MM5_g N_VDD_XI32/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI13/MM4 N_XI32/XI13/NET33_XI32/XI13/MM4_d
+ N_XI32/XI13/NET34_XI32/XI13/MM4_g N_VDD_XI32/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI13/MM10 N_XI32/XI13/NET35_XI32/XI13/MM10_d
+ N_XI32/XI13/NET36_XI32/XI13/MM10_g N_VDD_XI32/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI13/MM11 N_XI32/XI13/NET36_XI32/XI13/MM11_d
+ N_XI32/XI13/NET35_XI32/XI13/MM11_g N_VDD_XI32/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI14/MM2 N_XI32/XI14/NET34_XI32/XI14/MM2_d
+ N_XI32/XI14/NET33_XI32/XI14/MM2_g N_VSS_XI32/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI14/MM3 N_XI32/XI14/NET33_XI32/XI14/MM3_d N_WL<60>_XI32/XI14/MM3_g
+ N_BLN<1>_XI32/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI14/MM0 N_XI32/XI14/NET34_XI32/XI14/MM0_d N_WL<60>_XI32/XI14/MM0_g
+ N_BL<1>_XI32/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI14/MM1 N_XI32/XI14/NET33_XI32/XI14/MM1_d
+ N_XI32/XI14/NET34_XI32/XI14/MM1_g N_VSS_XI32/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI14/MM9 N_XI32/XI14/NET36_XI32/XI14/MM9_d N_WL<61>_XI32/XI14/MM9_g
+ N_BL<1>_XI32/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI14/MM6 N_XI32/XI14/NET35_XI32/XI14/MM6_d
+ N_XI32/XI14/NET36_XI32/XI14/MM6_g N_VSS_XI32/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI14/MM7 N_XI32/XI14/NET36_XI32/XI14/MM7_d
+ N_XI32/XI14/NET35_XI32/XI14/MM7_g N_VSS_XI32/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI14/MM8 N_XI32/XI14/NET35_XI32/XI14/MM8_d N_WL<61>_XI32/XI14/MM8_g
+ N_BLN<1>_XI32/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI14/MM5 N_XI32/XI14/NET34_XI32/XI14/MM5_d
+ N_XI32/XI14/NET33_XI32/XI14/MM5_g N_VDD_XI32/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI14/MM4 N_XI32/XI14/NET33_XI32/XI14/MM4_d
+ N_XI32/XI14/NET34_XI32/XI14/MM4_g N_VDD_XI32/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI14/MM10 N_XI32/XI14/NET35_XI32/XI14/MM10_d
+ N_XI32/XI14/NET36_XI32/XI14/MM10_g N_VDD_XI32/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI14/MM11 N_XI32/XI14/NET36_XI32/XI14/MM11_d
+ N_XI32/XI14/NET35_XI32/XI14/MM11_g N_VDD_XI32/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI15/MM2 N_XI32/XI15/NET34_XI32/XI15/MM2_d
+ N_XI32/XI15/NET33_XI32/XI15/MM2_g N_VSS_XI32/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI15/MM3 N_XI32/XI15/NET33_XI32/XI15/MM3_d N_WL<60>_XI32/XI15/MM3_g
+ N_BLN<0>_XI32/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI15/MM0 N_XI32/XI15/NET34_XI32/XI15/MM0_d N_WL<60>_XI32/XI15/MM0_g
+ N_BL<0>_XI32/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI15/MM1 N_XI32/XI15/NET33_XI32/XI15/MM1_d
+ N_XI32/XI15/NET34_XI32/XI15/MM1_g N_VSS_XI32/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI15/MM9 N_XI32/XI15/NET36_XI32/XI15/MM9_d N_WL<61>_XI32/XI15/MM9_g
+ N_BL<0>_XI32/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI15/MM6 N_XI32/XI15/NET35_XI32/XI15/MM6_d
+ N_XI32/XI15/NET36_XI32/XI15/MM6_g N_VSS_XI32/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI15/MM7 N_XI32/XI15/NET36_XI32/XI15/MM7_d
+ N_XI32/XI15/NET35_XI32/XI15/MM7_g N_VSS_XI32/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI32/XI15/MM8 N_XI32/XI15/NET35_XI32/XI15/MM8_d N_WL<61>_XI32/XI15/MM8_g
+ N_BLN<0>_XI32/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI32/XI15/MM5 N_XI32/XI15/NET34_XI32/XI15/MM5_d
+ N_XI32/XI15/NET33_XI32/XI15/MM5_g N_VDD_XI32/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI15/MM4 N_XI32/XI15/NET33_XI32/XI15/MM4_d
+ N_XI32/XI15/NET34_XI32/XI15/MM4_g N_VDD_XI32/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI15/MM10 N_XI32/XI15/NET35_XI32/XI15/MM10_d
+ N_XI32/XI15/NET36_XI32/XI15/MM10_g N_VDD_XI32/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI32/XI15/MM11 N_XI32/XI15/NET36_XI32/XI15/MM11_d
+ N_XI32/XI15/NET35_XI32/XI15/MM11_g N_VDD_XI32/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI0/MM2 N_XI33/XI0/NET34_XI33/XI0/MM2_d N_XI33/XI0/NET33_XI33/XI0/MM2_g
+ N_VSS_XI33/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI0/MM3 N_XI33/XI0/NET33_XI33/XI0/MM3_d N_WL<62>_XI33/XI0/MM3_g
+ N_BLN<15>_XI33/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI0/MM0 N_XI33/XI0/NET34_XI33/XI0/MM0_d N_WL<62>_XI33/XI0/MM0_g
+ N_BL<15>_XI33/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI0/MM1 N_XI33/XI0/NET33_XI33/XI0/MM1_d N_XI33/XI0/NET34_XI33/XI0/MM1_g
+ N_VSS_XI33/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI0/MM9 N_XI33/XI0/NET36_XI33/XI0/MM9_d N_WL<63>_XI33/XI0/MM9_g
+ N_BL<15>_XI33/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI0/MM6 N_XI33/XI0/NET35_XI33/XI0/MM6_d N_XI33/XI0/NET36_XI33/XI0/MM6_g
+ N_VSS_XI33/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI0/MM7 N_XI33/XI0/NET36_XI33/XI0/MM7_d N_XI33/XI0/NET35_XI33/XI0/MM7_g
+ N_VSS_XI33/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI0/MM8 N_XI33/XI0/NET35_XI33/XI0/MM8_d N_WL<63>_XI33/XI0/MM8_g
+ N_BLN<15>_XI33/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI0/MM5 N_XI33/XI0/NET34_XI33/XI0/MM5_d N_XI33/XI0/NET33_XI33/XI0/MM5_g
+ N_VDD_XI33/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI0/MM4 N_XI33/XI0/NET33_XI33/XI0/MM4_d N_XI33/XI0/NET34_XI33/XI0/MM4_g
+ N_VDD_XI33/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI0/MM10 N_XI33/XI0/NET35_XI33/XI0/MM10_d N_XI33/XI0/NET36_XI33/XI0/MM10_g
+ N_VDD_XI33/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI0/MM11 N_XI33/XI0/NET36_XI33/XI0/MM11_d N_XI33/XI0/NET35_XI33/XI0/MM11_g
+ N_VDD_XI33/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI1/MM2 N_XI33/XI1/NET34_XI33/XI1/MM2_d N_XI33/XI1/NET33_XI33/XI1/MM2_g
+ N_VSS_XI33/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI1/MM3 N_XI33/XI1/NET33_XI33/XI1/MM3_d N_WL<62>_XI33/XI1/MM3_g
+ N_BLN<14>_XI33/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI1/MM0 N_XI33/XI1/NET34_XI33/XI1/MM0_d N_WL<62>_XI33/XI1/MM0_g
+ N_BL<14>_XI33/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI1/MM1 N_XI33/XI1/NET33_XI33/XI1/MM1_d N_XI33/XI1/NET34_XI33/XI1/MM1_g
+ N_VSS_XI33/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI1/MM9 N_XI33/XI1/NET36_XI33/XI1/MM9_d N_WL<63>_XI33/XI1/MM9_g
+ N_BL<14>_XI33/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI1/MM6 N_XI33/XI1/NET35_XI33/XI1/MM6_d N_XI33/XI1/NET36_XI33/XI1/MM6_g
+ N_VSS_XI33/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI1/MM7 N_XI33/XI1/NET36_XI33/XI1/MM7_d N_XI33/XI1/NET35_XI33/XI1/MM7_g
+ N_VSS_XI33/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI1/MM8 N_XI33/XI1/NET35_XI33/XI1/MM8_d N_WL<63>_XI33/XI1/MM8_g
+ N_BLN<14>_XI33/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI1/MM5 N_XI33/XI1/NET34_XI33/XI1/MM5_d N_XI33/XI1/NET33_XI33/XI1/MM5_g
+ N_VDD_XI33/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI1/MM4 N_XI33/XI1/NET33_XI33/XI1/MM4_d N_XI33/XI1/NET34_XI33/XI1/MM4_g
+ N_VDD_XI33/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI1/MM10 N_XI33/XI1/NET35_XI33/XI1/MM10_d N_XI33/XI1/NET36_XI33/XI1/MM10_g
+ N_VDD_XI33/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI1/MM11 N_XI33/XI1/NET36_XI33/XI1/MM11_d N_XI33/XI1/NET35_XI33/XI1/MM11_g
+ N_VDD_XI33/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI2/MM2 N_XI33/XI2/NET34_XI33/XI2/MM2_d N_XI33/XI2/NET33_XI33/XI2/MM2_g
+ N_VSS_XI33/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI2/MM3 N_XI33/XI2/NET33_XI33/XI2/MM3_d N_WL<62>_XI33/XI2/MM3_g
+ N_BLN<13>_XI33/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI2/MM0 N_XI33/XI2/NET34_XI33/XI2/MM0_d N_WL<62>_XI33/XI2/MM0_g
+ N_BL<13>_XI33/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI2/MM1 N_XI33/XI2/NET33_XI33/XI2/MM1_d N_XI33/XI2/NET34_XI33/XI2/MM1_g
+ N_VSS_XI33/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI2/MM9 N_XI33/XI2/NET36_XI33/XI2/MM9_d N_WL<63>_XI33/XI2/MM9_g
+ N_BL<13>_XI33/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI2/MM6 N_XI33/XI2/NET35_XI33/XI2/MM6_d N_XI33/XI2/NET36_XI33/XI2/MM6_g
+ N_VSS_XI33/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI2/MM7 N_XI33/XI2/NET36_XI33/XI2/MM7_d N_XI33/XI2/NET35_XI33/XI2/MM7_g
+ N_VSS_XI33/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI2/MM8 N_XI33/XI2/NET35_XI33/XI2/MM8_d N_WL<63>_XI33/XI2/MM8_g
+ N_BLN<13>_XI33/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI2/MM5 N_XI33/XI2/NET34_XI33/XI2/MM5_d N_XI33/XI2/NET33_XI33/XI2/MM5_g
+ N_VDD_XI33/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI2/MM4 N_XI33/XI2/NET33_XI33/XI2/MM4_d N_XI33/XI2/NET34_XI33/XI2/MM4_g
+ N_VDD_XI33/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI2/MM10 N_XI33/XI2/NET35_XI33/XI2/MM10_d N_XI33/XI2/NET36_XI33/XI2/MM10_g
+ N_VDD_XI33/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI2/MM11 N_XI33/XI2/NET36_XI33/XI2/MM11_d N_XI33/XI2/NET35_XI33/XI2/MM11_g
+ N_VDD_XI33/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI3/MM2 N_XI33/XI3/NET34_XI33/XI3/MM2_d N_XI33/XI3/NET33_XI33/XI3/MM2_g
+ N_VSS_XI33/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI3/MM3 N_XI33/XI3/NET33_XI33/XI3/MM3_d N_WL<62>_XI33/XI3/MM3_g
+ N_BLN<12>_XI33/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI3/MM0 N_XI33/XI3/NET34_XI33/XI3/MM0_d N_WL<62>_XI33/XI3/MM0_g
+ N_BL<12>_XI33/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI3/MM1 N_XI33/XI3/NET33_XI33/XI3/MM1_d N_XI33/XI3/NET34_XI33/XI3/MM1_g
+ N_VSS_XI33/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI3/MM9 N_XI33/XI3/NET36_XI33/XI3/MM9_d N_WL<63>_XI33/XI3/MM9_g
+ N_BL<12>_XI33/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI3/MM6 N_XI33/XI3/NET35_XI33/XI3/MM6_d N_XI33/XI3/NET36_XI33/XI3/MM6_g
+ N_VSS_XI33/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI3/MM7 N_XI33/XI3/NET36_XI33/XI3/MM7_d N_XI33/XI3/NET35_XI33/XI3/MM7_g
+ N_VSS_XI33/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI3/MM8 N_XI33/XI3/NET35_XI33/XI3/MM8_d N_WL<63>_XI33/XI3/MM8_g
+ N_BLN<12>_XI33/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI3/MM5 N_XI33/XI3/NET34_XI33/XI3/MM5_d N_XI33/XI3/NET33_XI33/XI3/MM5_g
+ N_VDD_XI33/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI3/MM4 N_XI33/XI3/NET33_XI33/XI3/MM4_d N_XI33/XI3/NET34_XI33/XI3/MM4_g
+ N_VDD_XI33/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI3/MM10 N_XI33/XI3/NET35_XI33/XI3/MM10_d N_XI33/XI3/NET36_XI33/XI3/MM10_g
+ N_VDD_XI33/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI3/MM11 N_XI33/XI3/NET36_XI33/XI3/MM11_d N_XI33/XI3/NET35_XI33/XI3/MM11_g
+ N_VDD_XI33/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI4/MM2 N_XI33/XI4/NET34_XI33/XI4/MM2_d N_XI33/XI4/NET33_XI33/XI4/MM2_g
+ N_VSS_XI33/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI4/MM3 N_XI33/XI4/NET33_XI33/XI4/MM3_d N_WL<62>_XI33/XI4/MM3_g
+ N_BLN<11>_XI33/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI4/MM0 N_XI33/XI4/NET34_XI33/XI4/MM0_d N_WL<62>_XI33/XI4/MM0_g
+ N_BL<11>_XI33/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI4/MM1 N_XI33/XI4/NET33_XI33/XI4/MM1_d N_XI33/XI4/NET34_XI33/XI4/MM1_g
+ N_VSS_XI33/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI4/MM9 N_XI33/XI4/NET36_XI33/XI4/MM9_d N_WL<63>_XI33/XI4/MM9_g
+ N_BL<11>_XI33/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI4/MM6 N_XI33/XI4/NET35_XI33/XI4/MM6_d N_XI33/XI4/NET36_XI33/XI4/MM6_g
+ N_VSS_XI33/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI4/MM7 N_XI33/XI4/NET36_XI33/XI4/MM7_d N_XI33/XI4/NET35_XI33/XI4/MM7_g
+ N_VSS_XI33/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI4/MM8 N_XI33/XI4/NET35_XI33/XI4/MM8_d N_WL<63>_XI33/XI4/MM8_g
+ N_BLN<11>_XI33/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI4/MM5 N_XI33/XI4/NET34_XI33/XI4/MM5_d N_XI33/XI4/NET33_XI33/XI4/MM5_g
+ N_VDD_XI33/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI4/MM4 N_XI33/XI4/NET33_XI33/XI4/MM4_d N_XI33/XI4/NET34_XI33/XI4/MM4_g
+ N_VDD_XI33/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI4/MM10 N_XI33/XI4/NET35_XI33/XI4/MM10_d N_XI33/XI4/NET36_XI33/XI4/MM10_g
+ N_VDD_XI33/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI4/MM11 N_XI33/XI4/NET36_XI33/XI4/MM11_d N_XI33/XI4/NET35_XI33/XI4/MM11_g
+ N_VDD_XI33/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI5/MM2 N_XI33/XI5/NET34_XI33/XI5/MM2_d N_XI33/XI5/NET33_XI33/XI5/MM2_g
+ N_VSS_XI33/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI5/MM3 N_XI33/XI5/NET33_XI33/XI5/MM3_d N_WL<62>_XI33/XI5/MM3_g
+ N_BLN<10>_XI33/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI5/MM0 N_XI33/XI5/NET34_XI33/XI5/MM0_d N_WL<62>_XI33/XI5/MM0_g
+ N_BL<10>_XI33/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI5/MM1 N_XI33/XI5/NET33_XI33/XI5/MM1_d N_XI33/XI5/NET34_XI33/XI5/MM1_g
+ N_VSS_XI33/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI5/MM9 N_XI33/XI5/NET36_XI33/XI5/MM9_d N_WL<63>_XI33/XI5/MM9_g
+ N_BL<10>_XI33/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI5/MM6 N_XI33/XI5/NET35_XI33/XI5/MM6_d N_XI33/XI5/NET36_XI33/XI5/MM6_g
+ N_VSS_XI33/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI5/MM7 N_XI33/XI5/NET36_XI33/XI5/MM7_d N_XI33/XI5/NET35_XI33/XI5/MM7_g
+ N_VSS_XI33/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI5/MM8 N_XI33/XI5/NET35_XI33/XI5/MM8_d N_WL<63>_XI33/XI5/MM8_g
+ N_BLN<10>_XI33/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI5/MM5 N_XI33/XI5/NET34_XI33/XI5/MM5_d N_XI33/XI5/NET33_XI33/XI5/MM5_g
+ N_VDD_XI33/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI5/MM4 N_XI33/XI5/NET33_XI33/XI5/MM4_d N_XI33/XI5/NET34_XI33/XI5/MM4_g
+ N_VDD_XI33/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI5/MM10 N_XI33/XI5/NET35_XI33/XI5/MM10_d N_XI33/XI5/NET36_XI33/XI5/MM10_g
+ N_VDD_XI33/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI5/MM11 N_XI33/XI5/NET36_XI33/XI5/MM11_d N_XI33/XI5/NET35_XI33/XI5/MM11_g
+ N_VDD_XI33/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI6/MM2 N_XI33/XI6/NET34_XI33/XI6/MM2_d N_XI33/XI6/NET33_XI33/XI6/MM2_g
+ N_VSS_XI33/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM3 N_XI33/XI6/NET33_XI33/XI6/MM3_d N_WL<62>_XI33/XI6/MM3_g
+ N_BLN<9>_XI33/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM0 N_XI33/XI6/NET34_XI33/XI6/MM0_d N_WL<62>_XI33/XI6/MM0_g
+ N_BL<9>_XI33/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM1 N_XI33/XI6/NET33_XI33/XI6/MM1_d N_XI33/XI6/NET34_XI33/XI6/MM1_g
+ N_VSS_XI33/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM9 N_XI33/XI6/NET36_XI33/XI6/MM9_d N_WL<63>_XI33/XI6/MM9_g
+ N_BL<9>_XI33/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM6 N_XI33/XI6/NET35_XI33/XI6/MM6_d N_XI33/XI6/NET36_XI33/XI6/MM6_g
+ N_VSS_XI33/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM7 N_XI33/XI6/NET36_XI33/XI6/MM7_d N_XI33/XI6/NET35_XI33/XI6/MM7_g
+ N_VSS_XI33/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM8 N_XI33/XI6/NET35_XI33/XI6/MM8_d N_WL<63>_XI33/XI6/MM8_g
+ N_BLN<9>_XI33/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI6/MM5 N_XI33/XI6/NET34_XI33/XI6/MM5_d N_XI33/XI6/NET33_XI33/XI6/MM5_g
+ N_VDD_XI33/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI6/MM4 N_XI33/XI6/NET33_XI33/XI6/MM4_d N_XI33/XI6/NET34_XI33/XI6/MM4_g
+ N_VDD_XI33/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI6/MM10 N_XI33/XI6/NET35_XI33/XI6/MM10_d N_XI33/XI6/NET36_XI33/XI6/MM10_g
+ N_VDD_XI33/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI6/MM11 N_XI33/XI6/NET36_XI33/XI6/MM11_d N_XI33/XI6/NET35_XI33/XI6/MM11_g
+ N_VDD_XI33/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI7/MM2 N_XI33/XI7/NET34_XI33/XI7/MM2_d N_XI33/XI7/NET33_XI33/XI7/MM2_g
+ N_VSS_XI33/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM3 N_XI33/XI7/NET33_XI33/XI7/MM3_d N_WL<62>_XI33/XI7/MM3_g
+ N_BLN<8>_XI33/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM0 N_XI33/XI7/NET34_XI33/XI7/MM0_d N_WL<62>_XI33/XI7/MM0_g
+ N_BL<8>_XI33/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM1 N_XI33/XI7/NET33_XI33/XI7/MM1_d N_XI33/XI7/NET34_XI33/XI7/MM1_g
+ N_VSS_XI33/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM9 N_XI33/XI7/NET36_XI33/XI7/MM9_d N_WL<63>_XI33/XI7/MM9_g
+ N_BL<8>_XI33/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM6 N_XI33/XI7/NET35_XI33/XI7/MM6_d N_XI33/XI7/NET36_XI33/XI7/MM6_g
+ N_VSS_XI33/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM7 N_XI33/XI7/NET36_XI33/XI7/MM7_d N_XI33/XI7/NET35_XI33/XI7/MM7_g
+ N_VSS_XI33/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM8 N_XI33/XI7/NET35_XI33/XI7/MM8_d N_WL<63>_XI33/XI7/MM8_g
+ N_BLN<8>_XI33/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI7/MM5 N_XI33/XI7/NET34_XI33/XI7/MM5_d N_XI33/XI7/NET33_XI33/XI7/MM5_g
+ N_VDD_XI33/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI7/MM4 N_XI33/XI7/NET33_XI33/XI7/MM4_d N_XI33/XI7/NET34_XI33/XI7/MM4_g
+ N_VDD_XI33/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI7/MM10 N_XI33/XI7/NET35_XI33/XI7/MM10_d N_XI33/XI7/NET36_XI33/XI7/MM10_g
+ N_VDD_XI33/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI7/MM11 N_XI33/XI7/NET36_XI33/XI7/MM11_d N_XI33/XI7/NET35_XI33/XI7/MM11_g
+ N_VDD_XI33/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI8/MM2 N_XI33/XI8/NET34_XI33/XI8/MM2_d N_XI33/XI8/NET33_XI33/XI8/MM2_g
+ N_VSS_XI33/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM3 N_XI33/XI8/NET33_XI33/XI8/MM3_d N_WL<62>_XI33/XI8/MM3_g
+ N_BLN<7>_XI33/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM0 N_XI33/XI8/NET34_XI33/XI8/MM0_d N_WL<62>_XI33/XI8/MM0_g
+ N_BL<7>_XI33/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM1 N_XI33/XI8/NET33_XI33/XI8/MM1_d N_XI33/XI8/NET34_XI33/XI8/MM1_g
+ N_VSS_XI33/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM9 N_XI33/XI8/NET36_XI33/XI8/MM9_d N_WL<63>_XI33/XI8/MM9_g
+ N_BL<7>_XI33/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM6 N_XI33/XI8/NET35_XI33/XI8/MM6_d N_XI33/XI8/NET36_XI33/XI8/MM6_g
+ N_VSS_XI33/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM7 N_XI33/XI8/NET36_XI33/XI8/MM7_d N_XI33/XI8/NET35_XI33/XI8/MM7_g
+ N_VSS_XI33/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM8 N_XI33/XI8/NET35_XI33/XI8/MM8_d N_WL<63>_XI33/XI8/MM8_g
+ N_BLN<7>_XI33/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI8/MM5 N_XI33/XI8/NET34_XI33/XI8/MM5_d N_XI33/XI8/NET33_XI33/XI8/MM5_g
+ N_VDD_XI33/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI8/MM4 N_XI33/XI8/NET33_XI33/XI8/MM4_d N_XI33/XI8/NET34_XI33/XI8/MM4_g
+ N_VDD_XI33/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI8/MM10 N_XI33/XI8/NET35_XI33/XI8/MM10_d N_XI33/XI8/NET36_XI33/XI8/MM10_g
+ N_VDD_XI33/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI8/MM11 N_XI33/XI8/NET36_XI33/XI8/MM11_d N_XI33/XI8/NET35_XI33/XI8/MM11_g
+ N_VDD_XI33/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI9/MM2 N_XI33/XI9/NET34_XI33/XI9/MM2_d N_XI33/XI9/NET33_XI33/XI9/MM2_g
+ N_VSS_XI33/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM3 N_XI33/XI9/NET33_XI33/XI9/MM3_d N_WL<62>_XI33/XI9/MM3_g
+ N_BLN<6>_XI33/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM0 N_XI33/XI9/NET34_XI33/XI9/MM0_d N_WL<62>_XI33/XI9/MM0_g
+ N_BL<6>_XI33/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM1 N_XI33/XI9/NET33_XI33/XI9/MM1_d N_XI33/XI9/NET34_XI33/XI9/MM1_g
+ N_VSS_XI33/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM9 N_XI33/XI9/NET36_XI33/XI9/MM9_d N_WL<63>_XI33/XI9/MM9_g
+ N_BL<6>_XI33/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM6 N_XI33/XI9/NET35_XI33/XI9/MM6_d N_XI33/XI9/NET36_XI33/XI9/MM6_g
+ N_VSS_XI33/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM7 N_XI33/XI9/NET36_XI33/XI9/MM7_d N_XI33/XI9/NET35_XI33/XI9/MM7_g
+ N_VSS_XI33/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM8 N_XI33/XI9/NET35_XI33/XI9/MM8_d N_WL<63>_XI33/XI9/MM8_g
+ N_BLN<6>_XI33/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI9/MM5 N_XI33/XI9/NET34_XI33/XI9/MM5_d N_XI33/XI9/NET33_XI33/XI9/MM5_g
+ N_VDD_XI33/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI9/MM4 N_XI33/XI9/NET33_XI33/XI9/MM4_d N_XI33/XI9/NET34_XI33/XI9/MM4_g
+ N_VDD_XI33/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI9/MM10 N_XI33/XI9/NET35_XI33/XI9/MM10_d N_XI33/XI9/NET36_XI33/XI9/MM10_g
+ N_VDD_XI33/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI9/MM11 N_XI33/XI9/NET36_XI33/XI9/MM11_d N_XI33/XI9/NET35_XI33/XI9/MM11_g
+ N_VDD_XI33/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI10/MM2 N_XI33/XI10/NET34_XI33/XI10/MM2_d
+ N_XI33/XI10/NET33_XI33/XI10/MM2_g N_VSS_XI33/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI10/MM3 N_XI33/XI10/NET33_XI33/XI10/MM3_d N_WL<62>_XI33/XI10/MM3_g
+ N_BLN<5>_XI33/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI10/MM0 N_XI33/XI10/NET34_XI33/XI10/MM0_d N_WL<62>_XI33/XI10/MM0_g
+ N_BL<5>_XI33/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI10/MM1 N_XI33/XI10/NET33_XI33/XI10/MM1_d
+ N_XI33/XI10/NET34_XI33/XI10/MM1_g N_VSS_XI33/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI10/MM9 N_XI33/XI10/NET36_XI33/XI10/MM9_d N_WL<63>_XI33/XI10/MM9_g
+ N_BL<5>_XI33/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI10/MM6 N_XI33/XI10/NET35_XI33/XI10/MM6_d
+ N_XI33/XI10/NET36_XI33/XI10/MM6_g N_VSS_XI33/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI10/MM7 N_XI33/XI10/NET36_XI33/XI10/MM7_d
+ N_XI33/XI10/NET35_XI33/XI10/MM7_g N_VSS_XI33/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI10/MM8 N_XI33/XI10/NET35_XI33/XI10/MM8_d N_WL<63>_XI33/XI10/MM8_g
+ N_BLN<5>_XI33/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI10/MM5 N_XI33/XI10/NET34_XI33/XI10/MM5_d
+ N_XI33/XI10/NET33_XI33/XI10/MM5_g N_VDD_XI33/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI10/MM4 N_XI33/XI10/NET33_XI33/XI10/MM4_d
+ N_XI33/XI10/NET34_XI33/XI10/MM4_g N_VDD_XI33/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI10/MM10 N_XI33/XI10/NET35_XI33/XI10/MM10_d
+ N_XI33/XI10/NET36_XI33/XI10/MM10_g N_VDD_XI33/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI10/MM11 N_XI33/XI10/NET36_XI33/XI10/MM11_d
+ N_XI33/XI10/NET35_XI33/XI10/MM11_g N_VDD_XI33/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI11/MM2 N_XI33/XI11/NET34_XI33/XI11/MM2_d
+ N_XI33/XI11/NET33_XI33/XI11/MM2_g N_VSS_XI33/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI11/MM3 N_XI33/XI11/NET33_XI33/XI11/MM3_d N_WL<62>_XI33/XI11/MM3_g
+ N_BLN<4>_XI33/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI11/MM0 N_XI33/XI11/NET34_XI33/XI11/MM0_d N_WL<62>_XI33/XI11/MM0_g
+ N_BL<4>_XI33/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI11/MM1 N_XI33/XI11/NET33_XI33/XI11/MM1_d
+ N_XI33/XI11/NET34_XI33/XI11/MM1_g N_VSS_XI33/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI11/MM9 N_XI33/XI11/NET36_XI33/XI11/MM9_d N_WL<63>_XI33/XI11/MM9_g
+ N_BL<4>_XI33/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI11/MM6 N_XI33/XI11/NET35_XI33/XI11/MM6_d
+ N_XI33/XI11/NET36_XI33/XI11/MM6_g N_VSS_XI33/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI11/MM7 N_XI33/XI11/NET36_XI33/XI11/MM7_d
+ N_XI33/XI11/NET35_XI33/XI11/MM7_g N_VSS_XI33/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI11/MM8 N_XI33/XI11/NET35_XI33/XI11/MM8_d N_WL<63>_XI33/XI11/MM8_g
+ N_BLN<4>_XI33/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI11/MM5 N_XI33/XI11/NET34_XI33/XI11/MM5_d
+ N_XI33/XI11/NET33_XI33/XI11/MM5_g N_VDD_XI33/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI11/MM4 N_XI33/XI11/NET33_XI33/XI11/MM4_d
+ N_XI33/XI11/NET34_XI33/XI11/MM4_g N_VDD_XI33/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI11/MM10 N_XI33/XI11/NET35_XI33/XI11/MM10_d
+ N_XI33/XI11/NET36_XI33/XI11/MM10_g N_VDD_XI33/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI11/MM11 N_XI33/XI11/NET36_XI33/XI11/MM11_d
+ N_XI33/XI11/NET35_XI33/XI11/MM11_g N_VDD_XI33/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI12/MM2 N_XI33/XI12/NET34_XI33/XI12/MM2_d
+ N_XI33/XI12/NET33_XI33/XI12/MM2_g N_VSS_XI33/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI12/MM3 N_XI33/XI12/NET33_XI33/XI12/MM3_d N_WL<62>_XI33/XI12/MM3_g
+ N_BLN<3>_XI33/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI12/MM0 N_XI33/XI12/NET34_XI33/XI12/MM0_d N_WL<62>_XI33/XI12/MM0_g
+ N_BL<3>_XI33/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI12/MM1 N_XI33/XI12/NET33_XI33/XI12/MM1_d
+ N_XI33/XI12/NET34_XI33/XI12/MM1_g N_VSS_XI33/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI12/MM9 N_XI33/XI12/NET36_XI33/XI12/MM9_d N_WL<63>_XI33/XI12/MM9_g
+ N_BL<3>_XI33/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI12/MM6 N_XI33/XI12/NET35_XI33/XI12/MM6_d
+ N_XI33/XI12/NET36_XI33/XI12/MM6_g N_VSS_XI33/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI12/MM7 N_XI33/XI12/NET36_XI33/XI12/MM7_d
+ N_XI33/XI12/NET35_XI33/XI12/MM7_g N_VSS_XI33/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI12/MM8 N_XI33/XI12/NET35_XI33/XI12/MM8_d N_WL<63>_XI33/XI12/MM8_g
+ N_BLN<3>_XI33/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI12/MM5 N_XI33/XI12/NET34_XI33/XI12/MM5_d
+ N_XI33/XI12/NET33_XI33/XI12/MM5_g N_VDD_XI33/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI12/MM4 N_XI33/XI12/NET33_XI33/XI12/MM4_d
+ N_XI33/XI12/NET34_XI33/XI12/MM4_g N_VDD_XI33/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI12/MM10 N_XI33/XI12/NET35_XI33/XI12/MM10_d
+ N_XI33/XI12/NET36_XI33/XI12/MM10_g N_VDD_XI33/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI12/MM11 N_XI33/XI12/NET36_XI33/XI12/MM11_d
+ N_XI33/XI12/NET35_XI33/XI12/MM11_g N_VDD_XI33/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI13/MM2 N_XI33/XI13/NET34_XI33/XI13/MM2_d
+ N_XI33/XI13/NET33_XI33/XI13/MM2_g N_VSS_XI33/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI13/MM3 N_XI33/XI13/NET33_XI33/XI13/MM3_d N_WL<62>_XI33/XI13/MM3_g
+ N_BLN<2>_XI33/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI13/MM0 N_XI33/XI13/NET34_XI33/XI13/MM0_d N_WL<62>_XI33/XI13/MM0_g
+ N_BL<2>_XI33/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI13/MM1 N_XI33/XI13/NET33_XI33/XI13/MM1_d
+ N_XI33/XI13/NET34_XI33/XI13/MM1_g N_VSS_XI33/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI13/MM9 N_XI33/XI13/NET36_XI33/XI13/MM9_d N_WL<63>_XI33/XI13/MM9_g
+ N_BL<2>_XI33/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI13/MM6 N_XI33/XI13/NET35_XI33/XI13/MM6_d
+ N_XI33/XI13/NET36_XI33/XI13/MM6_g N_VSS_XI33/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI13/MM7 N_XI33/XI13/NET36_XI33/XI13/MM7_d
+ N_XI33/XI13/NET35_XI33/XI13/MM7_g N_VSS_XI33/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI13/MM8 N_XI33/XI13/NET35_XI33/XI13/MM8_d N_WL<63>_XI33/XI13/MM8_g
+ N_BLN<2>_XI33/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI13/MM5 N_XI33/XI13/NET34_XI33/XI13/MM5_d
+ N_XI33/XI13/NET33_XI33/XI13/MM5_g N_VDD_XI33/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI13/MM4 N_XI33/XI13/NET33_XI33/XI13/MM4_d
+ N_XI33/XI13/NET34_XI33/XI13/MM4_g N_VDD_XI33/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI13/MM10 N_XI33/XI13/NET35_XI33/XI13/MM10_d
+ N_XI33/XI13/NET36_XI33/XI13/MM10_g N_VDD_XI33/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI13/MM11 N_XI33/XI13/NET36_XI33/XI13/MM11_d
+ N_XI33/XI13/NET35_XI33/XI13/MM11_g N_VDD_XI33/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI14/MM2 N_XI33/XI14/NET34_XI33/XI14/MM2_d
+ N_XI33/XI14/NET33_XI33/XI14/MM2_g N_VSS_XI33/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI14/MM3 N_XI33/XI14/NET33_XI33/XI14/MM3_d N_WL<62>_XI33/XI14/MM3_g
+ N_BLN<1>_XI33/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI14/MM0 N_XI33/XI14/NET34_XI33/XI14/MM0_d N_WL<62>_XI33/XI14/MM0_g
+ N_BL<1>_XI33/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI14/MM1 N_XI33/XI14/NET33_XI33/XI14/MM1_d
+ N_XI33/XI14/NET34_XI33/XI14/MM1_g N_VSS_XI33/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI14/MM9 N_XI33/XI14/NET36_XI33/XI14/MM9_d N_WL<63>_XI33/XI14/MM9_g
+ N_BL<1>_XI33/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI14/MM6 N_XI33/XI14/NET35_XI33/XI14/MM6_d
+ N_XI33/XI14/NET36_XI33/XI14/MM6_g N_VSS_XI33/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI14/MM7 N_XI33/XI14/NET36_XI33/XI14/MM7_d
+ N_XI33/XI14/NET35_XI33/XI14/MM7_g N_VSS_XI33/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI14/MM8 N_XI33/XI14/NET35_XI33/XI14/MM8_d N_WL<63>_XI33/XI14/MM8_g
+ N_BLN<1>_XI33/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI14/MM5 N_XI33/XI14/NET34_XI33/XI14/MM5_d
+ N_XI33/XI14/NET33_XI33/XI14/MM5_g N_VDD_XI33/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI14/MM4 N_XI33/XI14/NET33_XI33/XI14/MM4_d
+ N_XI33/XI14/NET34_XI33/XI14/MM4_g N_VDD_XI33/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI14/MM10 N_XI33/XI14/NET35_XI33/XI14/MM10_d
+ N_XI33/XI14/NET36_XI33/XI14/MM10_g N_VDD_XI33/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI14/MM11 N_XI33/XI14/NET36_XI33/XI14/MM11_d
+ N_XI33/XI14/NET35_XI33/XI14/MM11_g N_VDD_XI33/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI15/MM2 N_XI33/XI15/NET34_XI33/XI15/MM2_d
+ N_XI33/XI15/NET33_XI33/XI15/MM2_g N_VSS_XI33/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI15/MM3 N_XI33/XI15/NET33_XI33/XI15/MM3_d N_WL<62>_XI33/XI15/MM3_g
+ N_BLN<0>_XI33/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI15/MM0 N_XI33/XI15/NET34_XI33/XI15/MM0_d N_WL<62>_XI33/XI15/MM0_g
+ N_BL<0>_XI33/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI15/MM1 N_XI33/XI15/NET33_XI33/XI15/MM1_d
+ N_XI33/XI15/NET34_XI33/XI15/MM1_g N_VSS_XI33/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI15/MM9 N_XI33/XI15/NET36_XI33/XI15/MM9_d N_WL<63>_XI33/XI15/MM9_g
+ N_BL<0>_XI33/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI15/MM6 N_XI33/XI15/NET35_XI33/XI15/MM6_d
+ N_XI33/XI15/NET36_XI33/XI15/MM6_g N_VSS_XI33/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI15/MM7 N_XI33/XI15/NET36_XI33/XI15/MM7_d
+ N_XI33/XI15/NET35_XI33/XI15/MM7_g N_VSS_XI33/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI33/XI15/MM8 N_XI33/XI15/NET35_XI33/XI15/MM8_d N_WL<63>_XI33/XI15/MM8_g
+ N_BLN<0>_XI33/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI33/XI15/MM5 N_XI33/XI15/NET34_XI33/XI15/MM5_d
+ N_XI33/XI15/NET33_XI33/XI15/MM5_g N_VDD_XI33/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI15/MM4 N_XI33/XI15/NET33_XI33/XI15/MM4_d
+ N_XI33/XI15/NET34_XI33/XI15/MM4_g N_VDD_XI33/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI15/MM10 N_XI33/XI15/NET35_XI33/XI15/MM10_d
+ N_XI33/XI15/NET36_XI33/XI15/MM10_g N_VDD_XI33/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI33/XI15/MM11 N_XI33/XI15/NET36_XI33/XI15/MM11_d
+ N_XI33/XI15/NET35_XI33/XI15/MM11_g N_VDD_XI33/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI0/MM2 N_XI34/XI0/NET34_XI34/XI0/MM2_d N_XI34/XI0/NET33_XI34/XI0/MM2_g
+ N_VSS_XI34/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI0/MM3 N_XI34/XI0/NET33_XI34/XI0/MM3_d N_WL<64>_XI34/XI0/MM3_g
+ N_BLN<15>_XI34/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI0/MM0 N_XI34/XI0/NET34_XI34/XI0/MM0_d N_WL<64>_XI34/XI0/MM0_g
+ N_BL<15>_XI34/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI0/MM1 N_XI34/XI0/NET33_XI34/XI0/MM1_d N_XI34/XI0/NET34_XI34/XI0/MM1_g
+ N_VSS_XI34/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI0/MM9 N_XI34/XI0/NET36_XI34/XI0/MM9_d N_WL<65>_XI34/XI0/MM9_g
+ N_BL<15>_XI34/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI0/MM6 N_XI34/XI0/NET35_XI34/XI0/MM6_d N_XI34/XI0/NET36_XI34/XI0/MM6_g
+ N_VSS_XI34/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI0/MM7 N_XI34/XI0/NET36_XI34/XI0/MM7_d N_XI34/XI0/NET35_XI34/XI0/MM7_g
+ N_VSS_XI34/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI0/MM8 N_XI34/XI0/NET35_XI34/XI0/MM8_d N_WL<65>_XI34/XI0/MM8_g
+ N_BLN<15>_XI34/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI0/MM5 N_XI34/XI0/NET34_XI34/XI0/MM5_d N_XI34/XI0/NET33_XI34/XI0/MM5_g
+ N_VDD_XI34/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI0/MM4 N_XI34/XI0/NET33_XI34/XI0/MM4_d N_XI34/XI0/NET34_XI34/XI0/MM4_g
+ N_VDD_XI34/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI0/MM10 N_XI34/XI0/NET35_XI34/XI0/MM10_d N_XI34/XI0/NET36_XI34/XI0/MM10_g
+ N_VDD_XI34/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI0/MM11 N_XI34/XI0/NET36_XI34/XI0/MM11_d N_XI34/XI0/NET35_XI34/XI0/MM11_g
+ N_VDD_XI34/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI1/MM2 N_XI34/XI1/NET34_XI34/XI1/MM2_d N_XI34/XI1/NET33_XI34/XI1/MM2_g
+ N_VSS_XI34/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI1/MM3 N_XI34/XI1/NET33_XI34/XI1/MM3_d N_WL<64>_XI34/XI1/MM3_g
+ N_BLN<14>_XI34/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI1/MM0 N_XI34/XI1/NET34_XI34/XI1/MM0_d N_WL<64>_XI34/XI1/MM0_g
+ N_BL<14>_XI34/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI1/MM1 N_XI34/XI1/NET33_XI34/XI1/MM1_d N_XI34/XI1/NET34_XI34/XI1/MM1_g
+ N_VSS_XI34/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI1/MM9 N_XI34/XI1/NET36_XI34/XI1/MM9_d N_WL<65>_XI34/XI1/MM9_g
+ N_BL<14>_XI34/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI1/MM6 N_XI34/XI1/NET35_XI34/XI1/MM6_d N_XI34/XI1/NET36_XI34/XI1/MM6_g
+ N_VSS_XI34/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI1/MM7 N_XI34/XI1/NET36_XI34/XI1/MM7_d N_XI34/XI1/NET35_XI34/XI1/MM7_g
+ N_VSS_XI34/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI1/MM8 N_XI34/XI1/NET35_XI34/XI1/MM8_d N_WL<65>_XI34/XI1/MM8_g
+ N_BLN<14>_XI34/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI1/MM5 N_XI34/XI1/NET34_XI34/XI1/MM5_d N_XI34/XI1/NET33_XI34/XI1/MM5_g
+ N_VDD_XI34/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI1/MM4 N_XI34/XI1/NET33_XI34/XI1/MM4_d N_XI34/XI1/NET34_XI34/XI1/MM4_g
+ N_VDD_XI34/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI1/MM10 N_XI34/XI1/NET35_XI34/XI1/MM10_d N_XI34/XI1/NET36_XI34/XI1/MM10_g
+ N_VDD_XI34/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI1/MM11 N_XI34/XI1/NET36_XI34/XI1/MM11_d N_XI34/XI1/NET35_XI34/XI1/MM11_g
+ N_VDD_XI34/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI2/MM2 N_XI34/XI2/NET34_XI34/XI2/MM2_d N_XI34/XI2/NET33_XI34/XI2/MM2_g
+ N_VSS_XI34/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI2/MM3 N_XI34/XI2/NET33_XI34/XI2/MM3_d N_WL<64>_XI34/XI2/MM3_g
+ N_BLN<13>_XI34/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI2/MM0 N_XI34/XI2/NET34_XI34/XI2/MM0_d N_WL<64>_XI34/XI2/MM0_g
+ N_BL<13>_XI34/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI2/MM1 N_XI34/XI2/NET33_XI34/XI2/MM1_d N_XI34/XI2/NET34_XI34/XI2/MM1_g
+ N_VSS_XI34/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI2/MM9 N_XI34/XI2/NET36_XI34/XI2/MM9_d N_WL<65>_XI34/XI2/MM9_g
+ N_BL<13>_XI34/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI2/MM6 N_XI34/XI2/NET35_XI34/XI2/MM6_d N_XI34/XI2/NET36_XI34/XI2/MM6_g
+ N_VSS_XI34/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI2/MM7 N_XI34/XI2/NET36_XI34/XI2/MM7_d N_XI34/XI2/NET35_XI34/XI2/MM7_g
+ N_VSS_XI34/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI2/MM8 N_XI34/XI2/NET35_XI34/XI2/MM8_d N_WL<65>_XI34/XI2/MM8_g
+ N_BLN<13>_XI34/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI2/MM5 N_XI34/XI2/NET34_XI34/XI2/MM5_d N_XI34/XI2/NET33_XI34/XI2/MM5_g
+ N_VDD_XI34/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI2/MM4 N_XI34/XI2/NET33_XI34/XI2/MM4_d N_XI34/XI2/NET34_XI34/XI2/MM4_g
+ N_VDD_XI34/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI2/MM10 N_XI34/XI2/NET35_XI34/XI2/MM10_d N_XI34/XI2/NET36_XI34/XI2/MM10_g
+ N_VDD_XI34/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI2/MM11 N_XI34/XI2/NET36_XI34/XI2/MM11_d N_XI34/XI2/NET35_XI34/XI2/MM11_g
+ N_VDD_XI34/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI3/MM2 N_XI34/XI3/NET34_XI34/XI3/MM2_d N_XI34/XI3/NET33_XI34/XI3/MM2_g
+ N_VSS_XI34/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI3/MM3 N_XI34/XI3/NET33_XI34/XI3/MM3_d N_WL<64>_XI34/XI3/MM3_g
+ N_BLN<12>_XI34/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI3/MM0 N_XI34/XI3/NET34_XI34/XI3/MM0_d N_WL<64>_XI34/XI3/MM0_g
+ N_BL<12>_XI34/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI3/MM1 N_XI34/XI3/NET33_XI34/XI3/MM1_d N_XI34/XI3/NET34_XI34/XI3/MM1_g
+ N_VSS_XI34/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI3/MM9 N_XI34/XI3/NET36_XI34/XI3/MM9_d N_WL<65>_XI34/XI3/MM9_g
+ N_BL<12>_XI34/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI3/MM6 N_XI34/XI3/NET35_XI34/XI3/MM6_d N_XI34/XI3/NET36_XI34/XI3/MM6_g
+ N_VSS_XI34/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI3/MM7 N_XI34/XI3/NET36_XI34/XI3/MM7_d N_XI34/XI3/NET35_XI34/XI3/MM7_g
+ N_VSS_XI34/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI3/MM8 N_XI34/XI3/NET35_XI34/XI3/MM8_d N_WL<65>_XI34/XI3/MM8_g
+ N_BLN<12>_XI34/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI3/MM5 N_XI34/XI3/NET34_XI34/XI3/MM5_d N_XI34/XI3/NET33_XI34/XI3/MM5_g
+ N_VDD_XI34/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI3/MM4 N_XI34/XI3/NET33_XI34/XI3/MM4_d N_XI34/XI3/NET34_XI34/XI3/MM4_g
+ N_VDD_XI34/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI3/MM10 N_XI34/XI3/NET35_XI34/XI3/MM10_d N_XI34/XI3/NET36_XI34/XI3/MM10_g
+ N_VDD_XI34/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI3/MM11 N_XI34/XI3/NET36_XI34/XI3/MM11_d N_XI34/XI3/NET35_XI34/XI3/MM11_g
+ N_VDD_XI34/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI4/MM2 N_XI34/XI4/NET34_XI34/XI4/MM2_d N_XI34/XI4/NET33_XI34/XI4/MM2_g
+ N_VSS_XI34/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI4/MM3 N_XI34/XI4/NET33_XI34/XI4/MM3_d N_WL<64>_XI34/XI4/MM3_g
+ N_BLN<11>_XI34/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI4/MM0 N_XI34/XI4/NET34_XI34/XI4/MM0_d N_WL<64>_XI34/XI4/MM0_g
+ N_BL<11>_XI34/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI4/MM1 N_XI34/XI4/NET33_XI34/XI4/MM1_d N_XI34/XI4/NET34_XI34/XI4/MM1_g
+ N_VSS_XI34/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI4/MM9 N_XI34/XI4/NET36_XI34/XI4/MM9_d N_WL<65>_XI34/XI4/MM9_g
+ N_BL<11>_XI34/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI4/MM6 N_XI34/XI4/NET35_XI34/XI4/MM6_d N_XI34/XI4/NET36_XI34/XI4/MM6_g
+ N_VSS_XI34/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI4/MM7 N_XI34/XI4/NET36_XI34/XI4/MM7_d N_XI34/XI4/NET35_XI34/XI4/MM7_g
+ N_VSS_XI34/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI4/MM8 N_XI34/XI4/NET35_XI34/XI4/MM8_d N_WL<65>_XI34/XI4/MM8_g
+ N_BLN<11>_XI34/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI4/MM5 N_XI34/XI4/NET34_XI34/XI4/MM5_d N_XI34/XI4/NET33_XI34/XI4/MM5_g
+ N_VDD_XI34/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI4/MM4 N_XI34/XI4/NET33_XI34/XI4/MM4_d N_XI34/XI4/NET34_XI34/XI4/MM4_g
+ N_VDD_XI34/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI4/MM10 N_XI34/XI4/NET35_XI34/XI4/MM10_d N_XI34/XI4/NET36_XI34/XI4/MM10_g
+ N_VDD_XI34/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI4/MM11 N_XI34/XI4/NET36_XI34/XI4/MM11_d N_XI34/XI4/NET35_XI34/XI4/MM11_g
+ N_VDD_XI34/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI5/MM2 N_XI34/XI5/NET34_XI34/XI5/MM2_d N_XI34/XI5/NET33_XI34/XI5/MM2_g
+ N_VSS_XI34/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI5/MM3 N_XI34/XI5/NET33_XI34/XI5/MM3_d N_WL<64>_XI34/XI5/MM3_g
+ N_BLN<10>_XI34/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI5/MM0 N_XI34/XI5/NET34_XI34/XI5/MM0_d N_WL<64>_XI34/XI5/MM0_g
+ N_BL<10>_XI34/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI5/MM1 N_XI34/XI5/NET33_XI34/XI5/MM1_d N_XI34/XI5/NET34_XI34/XI5/MM1_g
+ N_VSS_XI34/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI5/MM9 N_XI34/XI5/NET36_XI34/XI5/MM9_d N_WL<65>_XI34/XI5/MM9_g
+ N_BL<10>_XI34/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI5/MM6 N_XI34/XI5/NET35_XI34/XI5/MM6_d N_XI34/XI5/NET36_XI34/XI5/MM6_g
+ N_VSS_XI34/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI5/MM7 N_XI34/XI5/NET36_XI34/XI5/MM7_d N_XI34/XI5/NET35_XI34/XI5/MM7_g
+ N_VSS_XI34/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI5/MM8 N_XI34/XI5/NET35_XI34/XI5/MM8_d N_WL<65>_XI34/XI5/MM8_g
+ N_BLN<10>_XI34/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI5/MM5 N_XI34/XI5/NET34_XI34/XI5/MM5_d N_XI34/XI5/NET33_XI34/XI5/MM5_g
+ N_VDD_XI34/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI5/MM4 N_XI34/XI5/NET33_XI34/XI5/MM4_d N_XI34/XI5/NET34_XI34/XI5/MM4_g
+ N_VDD_XI34/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI5/MM10 N_XI34/XI5/NET35_XI34/XI5/MM10_d N_XI34/XI5/NET36_XI34/XI5/MM10_g
+ N_VDD_XI34/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI5/MM11 N_XI34/XI5/NET36_XI34/XI5/MM11_d N_XI34/XI5/NET35_XI34/XI5/MM11_g
+ N_VDD_XI34/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI6/MM2 N_XI34/XI6/NET34_XI34/XI6/MM2_d N_XI34/XI6/NET33_XI34/XI6/MM2_g
+ N_VSS_XI34/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM3 N_XI34/XI6/NET33_XI34/XI6/MM3_d N_WL<64>_XI34/XI6/MM3_g
+ N_BLN<9>_XI34/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM0 N_XI34/XI6/NET34_XI34/XI6/MM0_d N_WL<64>_XI34/XI6/MM0_g
+ N_BL<9>_XI34/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM1 N_XI34/XI6/NET33_XI34/XI6/MM1_d N_XI34/XI6/NET34_XI34/XI6/MM1_g
+ N_VSS_XI34/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM9 N_XI34/XI6/NET36_XI34/XI6/MM9_d N_WL<65>_XI34/XI6/MM9_g
+ N_BL<9>_XI34/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM6 N_XI34/XI6/NET35_XI34/XI6/MM6_d N_XI34/XI6/NET36_XI34/XI6/MM6_g
+ N_VSS_XI34/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM7 N_XI34/XI6/NET36_XI34/XI6/MM7_d N_XI34/XI6/NET35_XI34/XI6/MM7_g
+ N_VSS_XI34/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM8 N_XI34/XI6/NET35_XI34/XI6/MM8_d N_WL<65>_XI34/XI6/MM8_g
+ N_BLN<9>_XI34/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI6/MM5 N_XI34/XI6/NET34_XI34/XI6/MM5_d N_XI34/XI6/NET33_XI34/XI6/MM5_g
+ N_VDD_XI34/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI6/MM4 N_XI34/XI6/NET33_XI34/XI6/MM4_d N_XI34/XI6/NET34_XI34/XI6/MM4_g
+ N_VDD_XI34/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI6/MM10 N_XI34/XI6/NET35_XI34/XI6/MM10_d N_XI34/XI6/NET36_XI34/XI6/MM10_g
+ N_VDD_XI34/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI6/MM11 N_XI34/XI6/NET36_XI34/XI6/MM11_d N_XI34/XI6/NET35_XI34/XI6/MM11_g
+ N_VDD_XI34/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI7/MM2 N_XI34/XI7/NET34_XI34/XI7/MM2_d N_XI34/XI7/NET33_XI34/XI7/MM2_g
+ N_VSS_XI34/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM3 N_XI34/XI7/NET33_XI34/XI7/MM3_d N_WL<64>_XI34/XI7/MM3_g
+ N_BLN<8>_XI34/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM0 N_XI34/XI7/NET34_XI34/XI7/MM0_d N_WL<64>_XI34/XI7/MM0_g
+ N_BL<8>_XI34/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM1 N_XI34/XI7/NET33_XI34/XI7/MM1_d N_XI34/XI7/NET34_XI34/XI7/MM1_g
+ N_VSS_XI34/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM9 N_XI34/XI7/NET36_XI34/XI7/MM9_d N_WL<65>_XI34/XI7/MM9_g
+ N_BL<8>_XI34/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM6 N_XI34/XI7/NET35_XI34/XI7/MM6_d N_XI34/XI7/NET36_XI34/XI7/MM6_g
+ N_VSS_XI34/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM7 N_XI34/XI7/NET36_XI34/XI7/MM7_d N_XI34/XI7/NET35_XI34/XI7/MM7_g
+ N_VSS_XI34/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM8 N_XI34/XI7/NET35_XI34/XI7/MM8_d N_WL<65>_XI34/XI7/MM8_g
+ N_BLN<8>_XI34/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI7/MM5 N_XI34/XI7/NET34_XI34/XI7/MM5_d N_XI34/XI7/NET33_XI34/XI7/MM5_g
+ N_VDD_XI34/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI7/MM4 N_XI34/XI7/NET33_XI34/XI7/MM4_d N_XI34/XI7/NET34_XI34/XI7/MM4_g
+ N_VDD_XI34/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI7/MM10 N_XI34/XI7/NET35_XI34/XI7/MM10_d N_XI34/XI7/NET36_XI34/XI7/MM10_g
+ N_VDD_XI34/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI7/MM11 N_XI34/XI7/NET36_XI34/XI7/MM11_d N_XI34/XI7/NET35_XI34/XI7/MM11_g
+ N_VDD_XI34/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI8/MM2 N_XI34/XI8/NET34_XI34/XI8/MM2_d N_XI34/XI8/NET33_XI34/XI8/MM2_g
+ N_VSS_XI34/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM3 N_XI34/XI8/NET33_XI34/XI8/MM3_d N_WL<64>_XI34/XI8/MM3_g
+ N_BLN<7>_XI34/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM0 N_XI34/XI8/NET34_XI34/XI8/MM0_d N_WL<64>_XI34/XI8/MM0_g
+ N_BL<7>_XI34/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM1 N_XI34/XI8/NET33_XI34/XI8/MM1_d N_XI34/XI8/NET34_XI34/XI8/MM1_g
+ N_VSS_XI34/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM9 N_XI34/XI8/NET36_XI34/XI8/MM9_d N_WL<65>_XI34/XI8/MM9_g
+ N_BL<7>_XI34/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM6 N_XI34/XI8/NET35_XI34/XI8/MM6_d N_XI34/XI8/NET36_XI34/XI8/MM6_g
+ N_VSS_XI34/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM7 N_XI34/XI8/NET36_XI34/XI8/MM7_d N_XI34/XI8/NET35_XI34/XI8/MM7_g
+ N_VSS_XI34/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM8 N_XI34/XI8/NET35_XI34/XI8/MM8_d N_WL<65>_XI34/XI8/MM8_g
+ N_BLN<7>_XI34/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI8/MM5 N_XI34/XI8/NET34_XI34/XI8/MM5_d N_XI34/XI8/NET33_XI34/XI8/MM5_g
+ N_VDD_XI34/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI8/MM4 N_XI34/XI8/NET33_XI34/XI8/MM4_d N_XI34/XI8/NET34_XI34/XI8/MM4_g
+ N_VDD_XI34/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI8/MM10 N_XI34/XI8/NET35_XI34/XI8/MM10_d N_XI34/XI8/NET36_XI34/XI8/MM10_g
+ N_VDD_XI34/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI8/MM11 N_XI34/XI8/NET36_XI34/XI8/MM11_d N_XI34/XI8/NET35_XI34/XI8/MM11_g
+ N_VDD_XI34/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI9/MM2 N_XI34/XI9/NET34_XI34/XI9/MM2_d N_XI34/XI9/NET33_XI34/XI9/MM2_g
+ N_VSS_XI34/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM3 N_XI34/XI9/NET33_XI34/XI9/MM3_d N_WL<64>_XI34/XI9/MM3_g
+ N_BLN<6>_XI34/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM0 N_XI34/XI9/NET34_XI34/XI9/MM0_d N_WL<64>_XI34/XI9/MM0_g
+ N_BL<6>_XI34/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM1 N_XI34/XI9/NET33_XI34/XI9/MM1_d N_XI34/XI9/NET34_XI34/XI9/MM1_g
+ N_VSS_XI34/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM9 N_XI34/XI9/NET36_XI34/XI9/MM9_d N_WL<65>_XI34/XI9/MM9_g
+ N_BL<6>_XI34/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM6 N_XI34/XI9/NET35_XI34/XI9/MM6_d N_XI34/XI9/NET36_XI34/XI9/MM6_g
+ N_VSS_XI34/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM7 N_XI34/XI9/NET36_XI34/XI9/MM7_d N_XI34/XI9/NET35_XI34/XI9/MM7_g
+ N_VSS_XI34/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM8 N_XI34/XI9/NET35_XI34/XI9/MM8_d N_WL<65>_XI34/XI9/MM8_g
+ N_BLN<6>_XI34/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI9/MM5 N_XI34/XI9/NET34_XI34/XI9/MM5_d N_XI34/XI9/NET33_XI34/XI9/MM5_g
+ N_VDD_XI34/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI9/MM4 N_XI34/XI9/NET33_XI34/XI9/MM4_d N_XI34/XI9/NET34_XI34/XI9/MM4_g
+ N_VDD_XI34/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI9/MM10 N_XI34/XI9/NET35_XI34/XI9/MM10_d N_XI34/XI9/NET36_XI34/XI9/MM10_g
+ N_VDD_XI34/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI9/MM11 N_XI34/XI9/NET36_XI34/XI9/MM11_d N_XI34/XI9/NET35_XI34/XI9/MM11_g
+ N_VDD_XI34/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI10/MM2 N_XI34/XI10/NET34_XI34/XI10/MM2_d
+ N_XI34/XI10/NET33_XI34/XI10/MM2_g N_VSS_XI34/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI10/MM3 N_XI34/XI10/NET33_XI34/XI10/MM3_d N_WL<64>_XI34/XI10/MM3_g
+ N_BLN<5>_XI34/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI10/MM0 N_XI34/XI10/NET34_XI34/XI10/MM0_d N_WL<64>_XI34/XI10/MM0_g
+ N_BL<5>_XI34/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI10/MM1 N_XI34/XI10/NET33_XI34/XI10/MM1_d
+ N_XI34/XI10/NET34_XI34/XI10/MM1_g N_VSS_XI34/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI10/MM9 N_XI34/XI10/NET36_XI34/XI10/MM9_d N_WL<65>_XI34/XI10/MM9_g
+ N_BL<5>_XI34/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI10/MM6 N_XI34/XI10/NET35_XI34/XI10/MM6_d
+ N_XI34/XI10/NET36_XI34/XI10/MM6_g N_VSS_XI34/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI10/MM7 N_XI34/XI10/NET36_XI34/XI10/MM7_d
+ N_XI34/XI10/NET35_XI34/XI10/MM7_g N_VSS_XI34/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI10/MM8 N_XI34/XI10/NET35_XI34/XI10/MM8_d N_WL<65>_XI34/XI10/MM8_g
+ N_BLN<5>_XI34/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI10/MM5 N_XI34/XI10/NET34_XI34/XI10/MM5_d
+ N_XI34/XI10/NET33_XI34/XI10/MM5_g N_VDD_XI34/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI10/MM4 N_XI34/XI10/NET33_XI34/XI10/MM4_d
+ N_XI34/XI10/NET34_XI34/XI10/MM4_g N_VDD_XI34/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI10/MM10 N_XI34/XI10/NET35_XI34/XI10/MM10_d
+ N_XI34/XI10/NET36_XI34/XI10/MM10_g N_VDD_XI34/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI10/MM11 N_XI34/XI10/NET36_XI34/XI10/MM11_d
+ N_XI34/XI10/NET35_XI34/XI10/MM11_g N_VDD_XI34/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI11/MM2 N_XI34/XI11/NET34_XI34/XI11/MM2_d
+ N_XI34/XI11/NET33_XI34/XI11/MM2_g N_VSS_XI34/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI11/MM3 N_XI34/XI11/NET33_XI34/XI11/MM3_d N_WL<64>_XI34/XI11/MM3_g
+ N_BLN<4>_XI34/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI11/MM0 N_XI34/XI11/NET34_XI34/XI11/MM0_d N_WL<64>_XI34/XI11/MM0_g
+ N_BL<4>_XI34/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI11/MM1 N_XI34/XI11/NET33_XI34/XI11/MM1_d
+ N_XI34/XI11/NET34_XI34/XI11/MM1_g N_VSS_XI34/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI11/MM9 N_XI34/XI11/NET36_XI34/XI11/MM9_d N_WL<65>_XI34/XI11/MM9_g
+ N_BL<4>_XI34/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI11/MM6 N_XI34/XI11/NET35_XI34/XI11/MM6_d
+ N_XI34/XI11/NET36_XI34/XI11/MM6_g N_VSS_XI34/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI11/MM7 N_XI34/XI11/NET36_XI34/XI11/MM7_d
+ N_XI34/XI11/NET35_XI34/XI11/MM7_g N_VSS_XI34/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI11/MM8 N_XI34/XI11/NET35_XI34/XI11/MM8_d N_WL<65>_XI34/XI11/MM8_g
+ N_BLN<4>_XI34/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI11/MM5 N_XI34/XI11/NET34_XI34/XI11/MM5_d
+ N_XI34/XI11/NET33_XI34/XI11/MM5_g N_VDD_XI34/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI11/MM4 N_XI34/XI11/NET33_XI34/XI11/MM4_d
+ N_XI34/XI11/NET34_XI34/XI11/MM4_g N_VDD_XI34/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI11/MM10 N_XI34/XI11/NET35_XI34/XI11/MM10_d
+ N_XI34/XI11/NET36_XI34/XI11/MM10_g N_VDD_XI34/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI11/MM11 N_XI34/XI11/NET36_XI34/XI11/MM11_d
+ N_XI34/XI11/NET35_XI34/XI11/MM11_g N_VDD_XI34/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI12/MM2 N_XI34/XI12/NET34_XI34/XI12/MM2_d
+ N_XI34/XI12/NET33_XI34/XI12/MM2_g N_VSS_XI34/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI12/MM3 N_XI34/XI12/NET33_XI34/XI12/MM3_d N_WL<64>_XI34/XI12/MM3_g
+ N_BLN<3>_XI34/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI12/MM0 N_XI34/XI12/NET34_XI34/XI12/MM0_d N_WL<64>_XI34/XI12/MM0_g
+ N_BL<3>_XI34/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI12/MM1 N_XI34/XI12/NET33_XI34/XI12/MM1_d
+ N_XI34/XI12/NET34_XI34/XI12/MM1_g N_VSS_XI34/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI12/MM9 N_XI34/XI12/NET36_XI34/XI12/MM9_d N_WL<65>_XI34/XI12/MM9_g
+ N_BL<3>_XI34/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI12/MM6 N_XI34/XI12/NET35_XI34/XI12/MM6_d
+ N_XI34/XI12/NET36_XI34/XI12/MM6_g N_VSS_XI34/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI12/MM7 N_XI34/XI12/NET36_XI34/XI12/MM7_d
+ N_XI34/XI12/NET35_XI34/XI12/MM7_g N_VSS_XI34/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI12/MM8 N_XI34/XI12/NET35_XI34/XI12/MM8_d N_WL<65>_XI34/XI12/MM8_g
+ N_BLN<3>_XI34/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI12/MM5 N_XI34/XI12/NET34_XI34/XI12/MM5_d
+ N_XI34/XI12/NET33_XI34/XI12/MM5_g N_VDD_XI34/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI12/MM4 N_XI34/XI12/NET33_XI34/XI12/MM4_d
+ N_XI34/XI12/NET34_XI34/XI12/MM4_g N_VDD_XI34/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI12/MM10 N_XI34/XI12/NET35_XI34/XI12/MM10_d
+ N_XI34/XI12/NET36_XI34/XI12/MM10_g N_VDD_XI34/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI12/MM11 N_XI34/XI12/NET36_XI34/XI12/MM11_d
+ N_XI34/XI12/NET35_XI34/XI12/MM11_g N_VDD_XI34/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI13/MM2 N_XI34/XI13/NET34_XI34/XI13/MM2_d
+ N_XI34/XI13/NET33_XI34/XI13/MM2_g N_VSS_XI34/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI13/MM3 N_XI34/XI13/NET33_XI34/XI13/MM3_d N_WL<64>_XI34/XI13/MM3_g
+ N_BLN<2>_XI34/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI13/MM0 N_XI34/XI13/NET34_XI34/XI13/MM0_d N_WL<64>_XI34/XI13/MM0_g
+ N_BL<2>_XI34/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI13/MM1 N_XI34/XI13/NET33_XI34/XI13/MM1_d
+ N_XI34/XI13/NET34_XI34/XI13/MM1_g N_VSS_XI34/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI13/MM9 N_XI34/XI13/NET36_XI34/XI13/MM9_d N_WL<65>_XI34/XI13/MM9_g
+ N_BL<2>_XI34/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI13/MM6 N_XI34/XI13/NET35_XI34/XI13/MM6_d
+ N_XI34/XI13/NET36_XI34/XI13/MM6_g N_VSS_XI34/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI13/MM7 N_XI34/XI13/NET36_XI34/XI13/MM7_d
+ N_XI34/XI13/NET35_XI34/XI13/MM7_g N_VSS_XI34/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI13/MM8 N_XI34/XI13/NET35_XI34/XI13/MM8_d N_WL<65>_XI34/XI13/MM8_g
+ N_BLN<2>_XI34/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI13/MM5 N_XI34/XI13/NET34_XI34/XI13/MM5_d
+ N_XI34/XI13/NET33_XI34/XI13/MM5_g N_VDD_XI34/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI13/MM4 N_XI34/XI13/NET33_XI34/XI13/MM4_d
+ N_XI34/XI13/NET34_XI34/XI13/MM4_g N_VDD_XI34/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI13/MM10 N_XI34/XI13/NET35_XI34/XI13/MM10_d
+ N_XI34/XI13/NET36_XI34/XI13/MM10_g N_VDD_XI34/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI13/MM11 N_XI34/XI13/NET36_XI34/XI13/MM11_d
+ N_XI34/XI13/NET35_XI34/XI13/MM11_g N_VDD_XI34/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI14/MM2 N_XI34/XI14/NET34_XI34/XI14/MM2_d
+ N_XI34/XI14/NET33_XI34/XI14/MM2_g N_VSS_XI34/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI14/MM3 N_XI34/XI14/NET33_XI34/XI14/MM3_d N_WL<64>_XI34/XI14/MM3_g
+ N_BLN<1>_XI34/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI14/MM0 N_XI34/XI14/NET34_XI34/XI14/MM0_d N_WL<64>_XI34/XI14/MM0_g
+ N_BL<1>_XI34/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI14/MM1 N_XI34/XI14/NET33_XI34/XI14/MM1_d
+ N_XI34/XI14/NET34_XI34/XI14/MM1_g N_VSS_XI34/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI14/MM9 N_XI34/XI14/NET36_XI34/XI14/MM9_d N_WL<65>_XI34/XI14/MM9_g
+ N_BL<1>_XI34/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI14/MM6 N_XI34/XI14/NET35_XI34/XI14/MM6_d
+ N_XI34/XI14/NET36_XI34/XI14/MM6_g N_VSS_XI34/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI14/MM7 N_XI34/XI14/NET36_XI34/XI14/MM7_d
+ N_XI34/XI14/NET35_XI34/XI14/MM7_g N_VSS_XI34/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI14/MM8 N_XI34/XI14/NET35_XI34/XI14/MM8_d N_WL<65>_XI34/XI14/MM8_g
+ N_BLN<1>_XI34/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI14/MM5 N_XI34/XI14/NET34_XI34/XI14/MM5_d
+ N_XI34/XI14/NET33_XI34/XI14/MM5_g N_VDD_XI34/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI14/MM4 N_XI34/XI14/NET33_XI34/XI14/MM4_d
+ N_XI34/XI14/NET34_XI34/XI14/MM4_g N_VDD_XI34/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI14/MM10 N_XI34/XI14/NET35_XI34/XI14/MM10_d
+ N_XI34/XI14/NET36_XI34/XI14/MM10_g N_VDD_XI34/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI14/MM11 N_XI34/XI14/NET36_XI34/XI14/MM11_d
+ N_XI34/XI14/NET35_XI34/XI14/MM11_g N_VDD_XI34/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI15/MM2 N_XI34/XI15/NET34_XI34/XI15/MM2_d
+ N_XI34/XI15/NET33_XI34/XI15/MM2_g N_VSS_XI34/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI15/MM3 N_XI34/XI15/NET33_XI34/XI15/MM3_d N_WL<64>_XI34/XI15/MM3_g
+ N_BLN<0>_XI34/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI15/MM0 N_XI34/XI15/NET34_XI34/XI15/MM0_d N_WL<64>_XI34/XI15/MM0_g
+ N_BL<0>_XI34/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI15/MM1 N_XI34/XI15/NET33_XI34/XI15/MM1_d
+ N_XI34/XI15/NET34_XI34/XI15/MM1_g N_VSS_XI34/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI15/MM9 N_XI34/XI15/NET36_XI34/XI15/MM9_d N_WL<65>_XI34/XI15/MM9_g
+ N_BL<0>_XI34/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI15/MM6 N_XI34/XI15/NET35_XI34/XI15/MM6_d
+ N_XI34/XI15/NET36_XI34/XI15/MM6_g N_VSS_XI34/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI15/MM7 N_XI34/XI15/NET36_XI34/XI15/MM7_d
+ N_XI34/XI15/NET35_XI34/XI15/MM7_g N_VSS_XI34/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI34/XI15/MM8 N_XI34/XI15/NET35_XI34/XI15/MM8_d N_WL<65>_XI34/XI15/MM8_g
+ N_BLN<0>_XI34/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI34/XI15/MM5 N_XI34/XI15/NET34_XI34/XI15/MM5_d
+ N_XI34/XI15/NET33_XI34/XI15/MM5_g N_VDD_XI34/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI15/MM4 N_XI34/XI15/NET33_XI34/XI15/MM4_d
+ N_XI34/XI15/NET34_XI34/XI15/MM4_g N_VDD_XI34/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI15/MM10 N_XI34/XI15/NET35_XI34/XI15/MM10_d
+ N_XI34/XI15/NET36_XI34/XI15/MM10_g N_VDD_XI34/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI34/XI15/MM11 N_XI34/XI15/NET36_XI34/XI15/MM11_d
+ N_XI34/XI15/NET35_XI34/XI15/MM11_g N_VDD_XI34/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI0/MM2 N_XI35/XI0/NET34_XI35/XI0/MM2_d N_XI35/XI0/NET33_XI35/XI0/MM2_g
+ N_VSS_XI35/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI0/MM3 N_XI35/XI0/NET33_XI35/XI0/MM3_d N_WL<66>_XI35/XI0/MM3_g
+ N_BLN<15>_XI35/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI0/MM0 N_XI35/XI0/NET34_XI35/XI0/MM0_d N_WL<66>_XI35/XI0/MM0_g
+ N_BL<15>_XI35/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI0/MM1 N_XI35/XI0/NET33_XI35/XI0/MM1_d N_XI35/XI0/NET34_XI35/XI0/MM1_g
+ N_VSS_XI35/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI0/MM9 N_XI35/XI0/NET36_XI35/XI0/MM9_d N_WL<67>_XI35/XI0/MM9_g
+ N_BL<15>_XI35/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI0/MM6 N_XI35/XI0/NET35_XI35/XI0/MM6_d N_XI35/XI0/NET36_XI35/XI0/MM6_g
+ N_VSS_XI35/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI0/MM7 N_XI35/XI0/NET36_XI35/XI0/MM7_d N_XI35/XI0/NET35_XI35/XI0/MM7_g
+ N_VSS_XI35/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI0/MM8 N_XI35/XI0/NET35_XI35/XI0/MM8_d N_WL<67>_XI35/XI0/MM8_g
+ N_BLN<15>_XI35/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI0/MM5 N_XI35/XI0/NET34_XI35/XI0/MM5_d N_XI35/XI0/NET33_XI35/XI0/MM5_g
+ N_VDD_XI35/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI0/MM4 N_XI35/XI0/NET33_XI35/XI0/MM4_d N_XI35/XI0/NET34_XI35/XI0/MM4_g
+ N_VDD_XI35/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI0/MM10 N_XI35/XI0/NET35_XI35/XI0/MM10_d N_XI35/XI0/NET36_XI35/XI0/MM10_g
+ N_VDD_XI35/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI0/MM11 N_XI35/XI0/NET36_XI35/XI0/MM11_d N_XI35/XI0/NET35_XI35/XI0/MM11_g
+ N_VDD_XI35/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI1/MM2 N_XI35/XI1/NET34_XI35/XI1/MM2_d N_XI35/XI1/NET33_XI35/XI1/MM2_g
+ N_VSS_XI35/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI1/MM3 N_XI35/XI1/NET33_XI35/XI1/MM3_d N_WL<66>_XI35/XI1/MM3_g
+ N_BLN<14>_XI35/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI1/MM0 N_XI35/XI1/NET34_XI35/XI1/MM0_d N_WL<66>_XI35/XI1/MM0_g
+ N_BL<14>_XI35/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI1/MM1 N_XI35/XI1/NET33_XI35/XI1/MM1_d N_XI35/XI1/NET34_XI35/XI1/MM1_g
+ N_VSS_XI35/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI1/MM9 N_XI35/XI1/NET36_XI35/XI1/MM9_d N_WL<67>_XI35/XI1/MM9_g
+ N_BL<14>_XI35/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI1/MM6 N_XI35/XI1/NET35_XI35/XI1/MM6_d N_XI35/XI1/NET36_XI35/XI1/MM6_g
+ N_VSS_XI35/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI1/MM7 N_XI35/XI1/NET36_XI35/XI1/MM7_d N_XI35/XI1/NET35_XI35/XI1/MM7_g
+ N_VSS_XI35/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI1/MM8 N_XI35/XI1/NET35_XI35/XI1/MM8_d N_WL<67>_XI35/XI1/MM8_g
+ N_BLN<14>_XI35/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI1/MM5 N_XI35/XI1/NET34_XI35/XI1/MM5_d N_XI35/XI1/NET33_XI35/XI1/MM5_g
+ N_VDD_XI35/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI1/MM4 N_XI35/XI1/NET33_XI35/XI1/MM4_d N_XI35/XI1/NET34_XI35/XI1/MM4_g
+ N_VDD_XI35/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI1/MM10 N_XI35/XI1/NET35_XI35/XI1/MM10_d N_XI35/XI1/NET36_XI35/XI1/MM10_g
+ N_VDD_XI35/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI1/MM11 N_XI35/XI1/NET36_XI35/XI1/MM11_d N_XI35/XI1/NET35_XI35/XI1/MM11_g
+ N_VDD_XI35/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI2/MM2 N_XI35/XI2/NET34_XI35/XI2/MM2_d N_XI35/XI2/NET33_XI35/XI2/MM2_g
+ N_VSS_XI35/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI2/MM3 N_XI35/XI2/NET33_XI35/XI2/MM3_d N_WL<66>_XI35/XI2/MM3_g
+ N_BLN<13>_XI35/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI2/MM0 N_XI35/XI2/NET34_XI35/XI2/MM0_d N_WL<66>_XI35/XI2/MM0_g
+ N_BL<13>_XI35/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI2/MM1 N_XI35/XI2/NET33_XI35/XI2/MM1_d N_XI35/XI2/NET34_XI35/XI2/MM1_g
+ N_VSS_XI35/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI2/MM9 N_XI35/XI2/NET36_XI35/XI2/MM9_d N_WL<67>_XI35/XI2/MM9_g
+ N_BL<13>_XI35/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI2/MM6 N_XI35/XI2/NET35_XI35/XI2/MM6_d N_XI35/XI2/NET36_XI35/XI2/MM6_g
+ N_VSS_XI35/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI2/MM7 N_XI35/XI2/NET36_XI35/XI2/MM7_d N_XI35/XI2/NET35_XI35/XI2/MM7_g
+ N_VSS_XI35/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI2/MM8 N_XI35/XI2/NET35_XI35/XI2/MM8_d N_WL<67>_XI35/XI2/MM8_g
+ N_BLN<13>_XI35/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI2/MM5 N_XI35/XI2/NET34_XI35/XI2/MM5_d N_XI35/XI2/NET33_XI35/XI2/MM5_g
+ N_VDD_XI35/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI2/MM4 N_XI35/XI2/NET33_XI35/XI2/MM4_d N_XI35/XI2/NET34_XI35/XI2/MM4_g
+ N_VDD_XI35/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI2/MM10 N_XI35/XI2/NET35_XI35/XI2/MM10_d N_XI35/XI2/NET36_XI35/XI2/MM10_g
+ N_VDD_XI35/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI2/MM11 N_XI35/XI2/NET36_XI35/XI2/MM11_d N_XI35/XI2/NET35_XI35/XI2/MM11_g
+ N_VDD_XI35/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI3/MM2 N_XI35/XI3/NET34_XI35/XI3/MM2_d N_XI35/XI3/NET33_XI35/XI3/MM2_g
+ N_VSS_XI35/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI3/MM3 N_XI35/XI3/NET33_XI35/XI3/MM3_d N_WL<66>_XI35/XI3/MM3_g
+ N_BLN<12>_XI35/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI3/MM0 N_XI35/XI3/NET34_XI35/XI3/MM0_d N_WL<66>_XI35/XI3/MM0_g
+ N_BL<12>_XI35/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI3/MM1 N_XI35/XI3/NET33_XI35/XI3/MM1_d N_XI35/XI3/NET34_XI35/XI3/MM1_g
+ N_VSS_XI35/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI3/MM9 N_XI35/XI3/NET36_XI35/XI3/MM9_d N_WL<67>_XI35/XI3/MM9_g
+ N_BL<12>_XI35/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI3/MM6 N_XI35/XI3/NET35_XI35/XI3/MM6_d N_XI35/XI3/NET36_XI35/XI3/MM6_g
+ N_VSS_XI35/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI3/MM7 N_XI35/XI3/NET36_XI35/XI3/MM7_d N_XI35/XI3/NET35_XI35/XI3/MM7_g
+ N_VSS_XI35/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI3/MM8 N_XI35/XI3/NET35_XI35/XI3/MM8_d N_WL<67>_XI35/XI3/MM8_g
+ N_BLN<12>_XI35/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI3/MM5 N_XI35/XI3/NET34_XI35/XI3/MM5_d N_XI35/XI3/NET33_XI35/XI3/MM5_g
+ N_VDD_XI35/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI3/MM4 N_XI35/XI3/NET33_XI35/XI3/MM4_d N_XI35/XI3/NET34_XI35/XI3/MM4_g
+ N_VDD_XI35/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI3/MM10 N_XI35/XI3/NET35_XI35/XI3/MM10_d N_XI35/XI3/NET36_XI35/XI3/MM10_g
+ N_VDD_XI35/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI3/MM11 N_XI35/XI3/NET36_XI35/XI3/MM11_d N_XI35/XI3/NET35_XI35/XI3/MM11_g
+ N_VDD_XI35/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI4/MM2 N_XI35/XI4/NET34_XI35/XI4/MM2_d N_XI35/XI4/NET33_XI35/XI4/MM2_g
+ N_VSS_XI35/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI4/MM3 N_XI35/XI4/NET33_XI35/XI4/MM3_d N_WL<66>_XI35/XI4/MM3_g
+ N_BLN<11>_XI35/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI4/MM0 N_XI35/XI4/NET34_XI35/XI4/MM0_d N_WL<66>_XI35/XI4/MM0_g
+ N_BL<11>_XI35/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI4/MM1 N_XI35/XI4/NET33_XI35/XI4/MM1_d N_XI35/XI4/NET34_XI35/XI4/MM1_g
+ N_VSS_XI35/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI4/MM9 N_XI35/XI4/NET36_XI35/XI4/MM9_d N_WL<67>_XI35/XI4/MM9_g
+ N_BL<11>_XI35/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI4/MM6 N_XI35/XI4/NET35_XI35/XI4/MM6_d N_XI35/XI4/NET36_XI35/XI4/MM6_g
+ N_VSS_XI35/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI4/MM7 N_XI35/XI4/NET36_XI35/XI4/MM7_d N_XI35/XI4/NET35_XI35/XI4/MM7_g
+ N_VSS_XI35/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI4/MM8 N_XI35/XI4/NET35_XI35/XI4/MM8_d N_WL<67>_XI35/XI4/MM8_g
+ N_BLN<11>_XI35/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI4/MM5 N_XI35/XI4/NET34_XI35/XI4/MM5_d N_XI35/XI4/NET33_XI35/XI4/MM5_g
+ N_VDD_XI35/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI4/MM4 N_XI35/XI4/NET33_XI35/XI4/MM4_d N_XI35/XI4/NET34_XI35/XI4/MM4_g
+ N_VDD_XI35/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI4/MM10 N_XI35/XI4/NET35_XI35/XI4/MM10_d N_XI35/XI4/NET36_XI35/XI4/MM10_g
+ N_VDD_XI35/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI4/MM11 N_XI35/XI4/NET36_XI35/XI4/MM11_d N_XI35/XI4/NET35_XI35/XI4/MM11_g
+ N_VDD_XI35/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI5/MM2 N_XI35/XI5/NET34_XI35/XI5/MM2_d N_XI35/XI5/NET33_XI35/XI5/MM2_g
+ N_VSS_XI35/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI5/MM3 N_XI35/XI5/NET33_XI35/XI5/MM3_d N_WL<66>_XI35/XI5/MM3_g
+ N_BLN<10>_XI35/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI5/MM0 N_XI35/XI5/NET34_XI35/XI5/MM0_d N_WL<66>_XI35/XI5/MM0_g
+ N_BL<10>_XI35/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI5/MM1 N_XI35/XI5/NET33_XI35/XI5/MM1_d N_XI35/XI5/NET34_XI35/XI5/MM1_g
+ N_VSS_XI35/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI5/MM9 N_XI35/XI5/NET36_XI35/XI5/MM9_d N_WL<67>_XI35/XI5/MM9_g
+ N_BL<10>_XI35/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI5/MM6 N_XI35/XI5/NET35_XI35/XI5/MM6_d N_XI35/XI5/NET36_XI35/XI5/MM6_g
+ N_VSS_XI35/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI5/MM7 N_XI35/XI5/NET36_XI35/XI5/MM7_d N_XI35/XI5/NET35_XI35/XI5/MM7_g
+ N_VSS_XI35/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI5/MM8 N_XI35/XI5/NET35_XI35/XI5/MM8_d N_WL<67>_XI35/XI5/MM8_g
+ N_BLN<10>_XI35/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI5/MM5 N_XI35/XI5/NET34_XI35/XI5/MM5_d N_XI35/XI5/NET33_XI35/XI5/MM5_g
+ N_VDD_XI35/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI5/MM4 N_XI35/XI5/NET33_XI35/XI5/MM4_d N_XI35/XI5/NET34_XI35/XI5/MM4_g
+ N_VDD_XI35/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI5/MM10 N_XI35/XI5/NET35_XI35/XI5/MM10_d N_XI35/XI5/NET36_XI35/XI5/MM10_g
+ N_VDD_XI35/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI5/MM11 N_XI35/XI5/NET36_XI35/XI5/MM11_d N_XI35/XI5/NET35_XI35/XI5/MM11_g
+ N_VDD_XI35/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI6/MM2 N_XI35/XI6/NET34_XI35/XI6/MM2_d N_XI35/XI6/NET33_XI35/XI6/MM2_g
+ N_VSS_XI35/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM3 N_XI35/XI6/NET33_XI35/XI6/MM3_d N_WL<66>_XI35/XI6/MM3_g
+ N_BLN<9>_XI35/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM0 N_XI35/XI6/NET34_XI35/XI6/MM0_d N_WL<66>_XI35/XI6/MM0_g
+ N_BL<9>_XI35/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM1 N_XI35/XI6/NET33_XI35/XI6/MM1_d N_XI35/XI6/NET34_XI35/XI6/MM1_g
+ N_VSS_XI35/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM9 N_XI35/XI6/NET36_XI35/XI6/MM9_d N_WL<67>_XI35/XI6/MM9_g
+ N_BL<9>_XI35/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM6 N_XI35/XI6/NET35_XI35/XI6/MM6_d N_XI35/XI6/NET36_XI35/XI6/MM6_g
+ N_VSS_XI35/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM7 N_XI35/XI6/NET36_XI35/XI6/MM7_d N_XI35/XI6/NET35_XI35/XI6/MM7_g
+ N_VSS_XI35/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM8 N_XI35/XI6/NET35_XI35/XI6/MM8_d N_WL<67>_XI35/XI6/MM8_g
+ N_BLN<9>_XI35/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI6/MM5 N_XI35/XI6/NET34_XI35/XI6/MM5_d N_XI35/XI6/NET33_XI35/XI6/MM5_g
+ N_VDD_XI35/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI6/MM4 N_XI35/XI6/NET33_XI35/XI6/MM4_d N_XI35/XI6/NET34_XI35/XI6/MM4_g
+ N_VDD_XI35/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI6/MM10 N_XI35/XI6/NET35_XI35/XI6/MM10_d N_XI35/XI6/NET36_XI35/XI6/MM10_g
+ N_VDD_XI35/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI6/MM11 N_XI35/XI6/NET36_XI35/XI6/MM11_d N_XI35/XI6/NET35_XI35/XI6/MM11_g
+ N_VDD_XI35/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI7/MM2 N_XI35/XI7/NET34_XI35/XI7/MM2_d N_XI35/XI7/NET33_XI35/XI7/MM2_g
+ N_VSS_XI35/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM3 N_XI35/XI7/NET33_XI35/XI7/MM3_d N_WL<66>_XI35/XI7/MM3_g
+ N_BLN<8>_XI35/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM0 N_XI35/XI7/NET34_XI35/XI7/MM0_d N_WL<66>_XI35/XI7/MM0_g
+ N_BL<8>_XI35/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM1 N_XI35/XI7/NET33_XI35/XI7/MM1_d N_XI35/XI7/NET34_XI35/XI7/MM1_g
+ N_VSS_XI35/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM9 N_XI35/XI7/NET36_XI35/XI7/MM9_d N_WL<67>_XI35/XI7/MM9_g
+ N_BL<8>_XI35/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM6 N_XI35/XI7/NET35_XI35/XI7/MM6_d N_XI35/XI7/NET36_XI35/XI7/MM6_g
+ N_VSS_XI35/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM7 N_XI35/XI7/NET36_XI35/XI7/MM7_d N_XI35/XI7/NET35_XI35/XI7/MM7_g
+ N_VSS_XI35/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM8 N_XI35/XI7/NET35_XI35/XI7/MM8_d N_WL<67>_XI35/XI7/MM8_g
+ N_BLN<8>_XI35/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI7/MM5 N_XI35/XI7/NET34_XI35/XI7/MM5_d N_XI35/XI7/NET33_XI35/XI7/MM5_g
+ N_VDD_XI35/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI7/MM4 N_XI35/XI7/NET33_XI35/XI7/MM4_d N_XI35/XI7/NET34_XI35/XI7/MM4_g
+ N_VDD_XI35/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI7/MM10 N_XI35/XI7/NET35_XI35/XI7/MM10_d N_XI35/XI7/NET36_XI35/XI7/MM10_g
+ N_VDD_XI35/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI7/MM11 N_XI35/XI7/NET36_XI35/XI7/MM11_d N_XI35/XI7/NET35_XI35/XI7/MM11_g
+ N_VDD_XI35/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI8/MM2 N_XI35/XI8/NET34_XI35/XI8/MM2_d N_XI35/XI8/NET33_XI35/XI8/MM2_g
+ N_VSS_XI35/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM3 N_XI35/XI8/NET33_XI35/XI8/MM3_d N_WL<66>_XI35/XI8/MM3_g
+ N_BLN<7>_XI35/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM0 N_XI35/XI8/NET34_XI35/XI8/MM0_d N_WL<66>_XI35/XI8/MM0_g
+ N_BL<7>_XI35/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM1 N_XI35/XI8/NET33_XI35/XI8/MM1_d N_XI35/XI8/NET34_XI35/XI8/MM1_g
+ N_VSS_XI35/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM9 N_XI35/XI8/NET36_XI35/XI8/MM9_d N_WL<67>_XI35/XI8/MM9_g
+ N_BL<7>_XI35/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM6 N_XI35/XI8/NET35_XI35/XI8/MM6_d N_XI35/XI8/NET36_XI35/XI8/MM6_g
+ N_VSS_XI35/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM7 N_XI35/XI8/NET36_XI35/XI8/MM7_d N_XI35/XI8/NET35_XI35/XI8/MM7_g
+ N_VSS_XI35/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM8 N_XI35/XI8/NET35_XI35/XI8/MM8_d N_WL<67>_XI35/XI8/MM8_g
+ N_BLN<7>_XI35/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI8/MM5 N_XI35/XI8/NET34_XI35/XI8/MM5_d N_XI35/XI8/NET33_XI35/XI8/MM5_g
+ N_VDD_XI35/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI8/MM4 N_XI35/XI8/NET33_XI35/XI8/MM4_d N_XI35/XI8/NET34_XI35/XI8/MM4_g
+ N_VDD_XI35/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI8/MM10 N_XI35/XI8/NET35_XI35/XI8/MM10_d N_XI35/XI8/NET36_XI35/XI8/MM10_g
+ N_VDD_XI35/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI8/MM11 N_XI35/XI8/NET36_XI35/XI8/MM11_d N_XI35/XI8/NET35_XI35/XI8/MM11_g
+ N_VDD_XI35/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI9/MM2 N_XI35/XI9/NET34_XI35/XI9/MM2_d N_XI35/XI9/NET33_XI35/XI9/MM2_g
+ N_VSS_XI35/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM3 N_XI35/XI9/NET33_XI35/XI9/MM3_d N_WL<66>_XI35/XI9/MM3_g
+ N_BLN<6>_XI35/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM0 N_XI35/XI9/NET34_XI35/XI9/MM0_d N_WL<66>_XI35/XI9/MM0_g
+ N_BL<6>_XI35/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM1 N_XI35/XI9/NET33_XI35/XI9/MM1_d N_XI35/XI9/NET34_XI35/XI9/MM1_g
+ N_VSS_XI35/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM9 N_XI35/XI9/NET36_XI35/XI9/MM9_d N_WL<67>_XI35/XI9/MM9_g
+ N_BL<6>_XI35/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM6 N_XI35/XI9/NET35_XI35/XI9/MM6_d N_XI35/XI9/NET36_XI35/XI9/MM6_g
+ N_VSS_XI35/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM7 N_XI35/XI9/NET36_XI35/XI9/MM7_d N_XI35/XI9/NET35_XI35/XI9/MM7_g
+ N_VSS_XI35/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM8 N_XI35/XI9/NET35_XI35/XI9/MM8_d N_WL<67>_XI35/XI9/MM8_g
+ N_BLN<6>_XI35/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI9/MM5 N_XI35/XI9/NET34_XI35/XI9/MM5_d N_XI35/XI9/NET33_XI35/XI9/MM5_g
+ N_VDD_XI35/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI9/MM4 N_XI35/XI9/NET33_XI35/XI9/MM4_d N_XI35/XI9/NET34_XI35/XI9/MM4_g
+ N_VDD_XI35/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI9/MM10 N_XI35/XI9/NET35_XI35/XI9/MM10_d N_XI35/XI9/NET36_XI35/XI9/MM10_g
+ N_VDD_XI35/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI9/MM11 N_XI35/XI9/NET36_XI35/XI9/MM11_d N_XI35/XI9/NET35_XI35/XI9/MM11_g
+ N_VDD_XI35/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI10/MM2 N_XI35/XI10/NET34_XI35/XI10/MM2_d
+ N_XI35/XI10/NET33_XI35/XI10/MM2_g N_VSS_XI35/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI10/MM3 N_XI35/XI10/NET33_XI35/XI10/MM3_d N_WL<66>_XI35/XI10/MM3_g
+ N_BLN<5>_XI35/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI10/MM0 N_XI35/XI10/NET34_XI35/XI10/MM0_d N_WL<66>_XI35/XI10/MM0_g
+ N_BL<5>_XI35/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI10/MM1 N_XI35/XI10/NET33_XI35/XI10/MM1_d
+ N_XI35/XI10/NET34_XI35/XI10/MM1_g N_VSS_XI35/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI10/MM9 N_XI35/XI10/NET36_XI35/XI10/MM9_d N_WL<67>_XI35/XI10/MM9_g
+ N_BL<5>_XI35/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI10/MM6 N_XI35/XI10/NET35_XI35/XI10/MM6_d
+ N_XI35/XI10/NET36_XI35/XI10/MM6_g N_VSS_XI35/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI10/MM7 N_XI35/XI10/NET36_XI35/XI10/MM7_d
+ N_XI35/XI10/NET35_XI35/XI10/MM7_g N_VSS_XI35/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI10/MM8 N_XI35/XI10/NET35_XI35/XI10/MM8_d N_WL<67>_XI35/XI10/MM8_g
+ N_BLN<5>_XI35/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI10/MM5 N_XI35/XI10/NET34_XI35/XI10/MM5_d
+ N_XI35/XI10/NET33_XI35/XI10/MM5_g N_VDD_XI35/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI10/MM4 N_XI35/XI10/NET33_XI35/XI10/MM4_d
+ N_XI35/XI10/NET34_XI35/XI10/MM4_g N_VDD_XI35/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI10/MM10 N_XI35/XI10/NET35_XI35/XI10/MM10_d
+ N_XI35/XI10/NET36_XI35/XI10/MM10_g N_VDD_XI35/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI10/MM11 N_XI35/XI10/NET36_XI35/XI10/MM11_d
+ N_XI35/XI10/NET35_XI35/XI10/MM11_g N_VDD_XI35/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI11/MM2 N_XI35/XI11/NET34_XI35/XI11/MM2_d
+ N_XI35/XI11/NET33_XI35/XI11/MM2_g N_VSS_XI35/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI11/MM3 N_XI35/XI11/NET33_XI35/XI11/MM3_d N_WL<66>_XI35/XI11/MM3_g
+ N_BLN<4>_XI35/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI11/MM0 N_XI35/XI11/NET34_XI35/XI11/MM0_d N_WL<66>_XI35/XI11/MM0_g
+ N_BL<4>_XI35/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI11/MM1 N_XI35/XI11/NET33_XI35/XI11/MM1_d
+ N_XI35/XI11/NET34_XI35/XI11/MM1_g N_VSS_XI35/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI11/MM9 N_XI35/XI11/NET36_XI35/XI11/MM9_d N_WL<67>_XI35/XI11/MM9_g
+ N_BL<4>_XI35/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI11/MM6 N_XI35/XI11/NET35_XI35/XI11/MM6_d
+ N_XI35/XI11/NET36_XI35/XI11/MM6_g N_VSS_XI35/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI11/MM7 N_XI35/XI11/NET36_XI35/XI11/MM7_d
+ N_XI35/XI11/NET35_XI35/XI11/MM7_g N_VSS_XI35/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI11/MM8 N_XI35/XI11/NET35_XI35/XI11/MM8_d N_WL<67>_XI35/XI11/MM8_g
+ N_BLN<4>_XI35/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI11/MM5 N_XI35/XI11/NET34_XI35/XI11/MM5_d
+ N_XI35/XI11/NET33_XI35/XI11/MM5_g N_VDD_XI35/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI11/MM4 N_XI35/XI11/NET33_XI35/XI11/MM4_d
+ N_XI35/XI11/NET34_XI35/XI11/MM4_g N_VDD_XI35/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI11/MM10 N_XI35/XI11/NET35_XI35/XI11/MM10_d
+ N_XI35/XI11/NET36_XI35/XI11/MM10_g N_VDD_XI35/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI11/MM11 N_XI35/XI11/NET36_XI35/XI11/MM11_d
+ N_XI35/XI11/NET35_XI35/XI11/MM11_g N_VDD_XI35/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI12/MM2 N_XI35/XI12/NET34_XI35/XI12/MM2_d
+ N_XI35/XI12/NET33_XI35/XI12/MM2_g N_VSS_XI35/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI12/MM3 N_XI35/XI12/NET33_XI35/XI12/MM3_d N_WL<66>_XI35/XI12/MM3_g
+ N_BLN<3>_XI35/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI12/MM0 N_XI35/XI12/NET34_XI35/XI12/MM0_d N_WL<66>_XI35/XI12/MM0_g
+ N_BL<3>_XI35/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI12/MM1 N_XI35/XI12/NET33_XI35/XI12/MM1_d
+ N_XI35/XI12/NET34_XI35/XI12/MM1_g N_VSS_XI35/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI12/MM9 N_XI35/XI12/NET36_XI35/XI12/MM9_d N_WL<67>_XI35/XI12/MM9_g
+ N_BL<3>_XI35/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI12/MM6 N_XI35/XI12/NET35_XI35/XI12/MM6_d
+ N_XI35/XI12/NET36_XI35/XI12/MM6_g N_VSS_XI35/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI12/MM7 N_XI35/XI12/NET36_XI35/XI12/MM7_d
+ N_XI35/XI12/NET35_XI35/XI12/MM7_g N_VSS_XI35/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI12/MM8 N_XI35/XI12/NET35_XI35/XI12/MM8_d N_WL<67>_XI35/XI12/MM8_g
+ N_BLN<3>_XI35/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI12/MM5 N_XI35/XI12/NET34_XI35/XI12/MM5_d
+ N_XI35/XI12/NET33_XI35/XI12/MM5_g N_VDD_XI35/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI12/MM4 N_XI35/XI12/NET33_XI35/XI12/MM4_d
+ N_XI35/XI12/NET34_XI35/XI12/MM4_g N_VDD_XI35/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI12/MM10 N_XI35/XI12/NET35_XI35/XI12/MM10_d
+ N_XI35/XI12/NET36_XI35/XI12/MM10_g N_VDD_XI35/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI12/MM11 N_XI35/XI12/NET36_XI35/XI12/MM11_d
+ N_XI35/XI12/NET35_XI35/XI12/MM11_g N_VDD_XI35/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI13/MM2 N_XI35/XI13/NET34_XI35/XI13/MM2_d
+ N_XI35/XI13/NET33_XI35/XI13/MM2_g N_VSS_XI35/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI13/MM3 N_XI35/XI13/NET33_XI35/XI13/MM3_d N_WL<66>_XI35/XI13/MM3_g
+ N_BLN<2>_XI35/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI13/MM0 N_XI35/XI13/NET34_XI35/XI13/MM0_d N_WL<66>_XI35/XI13/MM0_g
+ N_BL<2>_XI35/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI13/MM1 N_XI35/XI13/NET33_XI35/XI13/MM1_d
+ N_XI35/XI13/NET34_XI35/XI13/MM1_g N_VSS_XI35/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI13/MM9 N_XI35/XI13/NET36_XI35/XI13/MM9_d N_WL<67>_XI35/XI13/MM9_g
+ N_BL<2>_XI35/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI13/MM6 N_XI35/XI13/NET35_XI35/XI13/MM6_d
+ N_XI35/XI13/NET36_XI35/XI13/MM6_g N_VSS_XI35/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI13/MM7 N_XI35/XI13/NET36_XI35/XI13/MM7_d
+ N_XI35/XI13/NET35_XI35/XI13/MM7_g N_VSS_XI35/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI13/MM8 N_XI35/XI13/NET35_XI35/XI13/MM8_d N_WL<67>_XI35/XI13/MM8_g
+ N_BLN<2>_XI35/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI13/MM5 N_XI35/XI13/NET34_XI35/XI13/MM5_d
+ N_XI35/XI13/NET33_XI35/XI13/MM5_g N_VDD_XI35/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI13/MM4 N_XI35/XI13/NET33_XI35/XI13/MM4_d
+ N_XI35/XI13/NET34_XI35/XI13/MM4_g N_VDD_XI35/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI13/MM10 N_XI35/XI13/NET35_XI35/XI13/MM10_d
+ N_XI35/XI13/NET36_XI35/XI13/MM10_g N_VDD_XI35/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI13/MM11 N_XI35/XI13/NET36_XI35/XI13/MM11_d
+ N_XI35/XI13/NET35_XI35/XI13/MM11_g N_VDD_XI35/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI14/MM2 N_XI35/XI14/NET34_XI35/XI14/MM2_d
+ N_XI35/XI14/NET33_XI35/XI14/MM2_g N_VSS_XI35/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI14/MM3 N_XI35/XI14/NET33_XI35/XI14/MM3_d N_WL<66>_XI35/XI14/MM3_g
+ N_BLN<1>_XI35/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI14/MM0 N_XI35/XI14/NET34_XI35/XI14/MM0_d N_WL<66>_XI35/XI14/MM0_g
+ N_BL<1>_XI35/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI14/MM1 N_XI35/XI14/NET33_XI35/XI14/MM1_d
+ N_XI35/XI14/NET34_XI35/XI14/MM1_g N_VSS_XI35/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI14/MM9 N_XI35/XI14/NET36_XI35/XI14/MM9_d N_WL<67>_XI35/XI14/MM9_g
+ N_BL<1>_XI35/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI14/MM6 N_XI35/XI14/NET35_XI35/XI14/MM6_d
+ N_XI35/XI14/NET36_XI35/XI14/MM6_g N_VSS_XI35/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI14/MM7 N_XI35/XI14/NET36_XI35/XI14/MM7_d
+ N_XI35/XI14/NET35_XI35/XI14/MM7_g N_VSS_XI35/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI14/MM8 N_XI35/XI14/NET35_XI35/XI14/MM8_d N_WL<67>_XI35/XI14/MM8_g
+ N_BLN<1>_XI35/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI14/MM5 N_XI35/XI14/NET34_XI35/XI14/MM5_d
+ N_XI35/XI14/NET33_XI35/XI14/MM5_g N_VDD_XI35/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI14/MM4 N_XI35/XI14/NET33_XI35/XI14/MM4_d
+ N_XI35/XI14/NET34_XI35/XI14/MM4_g N_VDD_XI35/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI14/MM10 N_XI35/XI14/NET35_XI35/XI14/MM10_d
+ N_XI35/XI14/NET36_XI35/XI14/MM10_g N_VDD_XI35/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI14/MM11 N_XI35/XI14/NET36_XI35/XI14/MM11_d
+ N_XI35/XI14/NET35_XI35/XI14/MM11_g N_VDD_XI35/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI15/MM2 N_XI35/XI15/NET34_XI35/XI15/MM2_d
+ N_XI35/XI15/NET33_XI35/XI15/MM2_g N_VSS_XI35/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI15/MM3 N_XI35/XI15/NET33_XI35/XI15/MM3_d N_WL<66>_XI35/XI15/MM3_g
+ N_BLN<0>_XI35/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI15/MM0 N_XI35/XI15/NET34_XI35/XI15/MM0_d N_WL<66>_XI35/XI15/MM0_g
+ N_BL<0>_XI35/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI15/MM1 N_XI35/XI15/NET33_XI35/XI15/MM1_d
+ N_XI35/XI15/NET34_XI35/XI15/MM1_g N_VSS_XI35/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI15/MM9 N_XI35/XI15/NET36_XI35/XI15/MM9_d N_WL<67>_XI35/XI15/MM9_g
+ N_BL<0>_XI35/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI15/MM6 N_XI35/XI15/NET35_XI35/XI15/MM6_d
+ N_XI35/XI15/NET36_XI35/XI15/MM6_g N_VSS_XI35/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI15/MM7 N_XI35/XI15/NET36_XI35/XI15/MM7_d
+ N_XI35/XI15/NET35_XI35/XI15/MM7_g N_VSS_XI35/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI35/XI15/MM8 N_XI35/XI15/NET35_XI35/XI15/MM8_d N_WL<67>_XI35/XI15/MM8_g
+ N_BLN<0>_XI35/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI35/XI15/MM5 N_XI35/XI15/NET34_XI35/XI15/MM5_d
+ N_XI35/XI15/NET33_XI35/XI15/MM5_g N_VDD_XI35/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI15/MM4 N_XI35/XI15/NET33_XI35/XI15/MM4_d
+ N_XI35/XI15/NET34_XI35/XI15/MM4_g N_VDD_XI35/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI15/MM10 N_XI35/XI15/NET35_XI35/XI15/MM10_d
+ N_XI35/XI15/NET36_XI35/XI15/MM10_g N_VDD_XI35/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI35/XI15/MM11 N_XI35/XI15/NET36_XI35/XI15/MM11_d
+ N_XI35/XI15/NET35_XI35/XI15/MM11_g N_VDD_XI35/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI0/MM2 N_XI36/XI0/NET34_XI36/XI0/MM2_d N_XI36/XI0/NET33_XI36/XI0/MM2_g
+ N_VSS_XI36/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI0/MM3 N_XI36/XI0/NET33_XI36/XI0/MM3_d N_WL<68>_XI36/XI0/MM3_g
+ N_BLN<15>_XI36/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI0/MM0 N_XI36/XI0/NET34_XI36/XI0/MM0_d N_WL<68>_XI36/XI0/MM0_g
+ N_BL<15>_XI36/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI0/MM1 N_XI36/XI0/NET33_XI36/XI0/MM1_d N_XI36/XI0/NET34_XI36/XI0/MM1_g
+ N_VSS_XI36/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI0/MM9 N_XI36/XI0/NET36_XI36/XI0/MM9_d N_WL<69>_XI36/XI0/MM9_g
+ N_BL<15>_XI36/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI0/MM6 N_XI36/XI0/NET35_XI36/XI0/MM6_d N_XI36/XI0/NET36_XI36/XI0/MM6_g
+ N_VSS_XI36/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI0/MM7 N_XI36/XI0/NET36_XI36/XI0/MM7_d N_XI36/XI0/NET35_XI36/XI0/MM7_g
+ N_VSS_XI36/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI0/MM8 N_XI36/XI0/NET35_XI36/XI0/MM8_d N_WL<69>_XI36/XI0/MM8_g
+ N_BLN<15>_XI36/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI0/MM5 N_XI36/XI0/NET34_XI36/XI0/MM5_d N_XI36/XI0/NET33_XI36/XI0/MM5_g
+ N_VDD_XI36/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI0/MM4 N_XI36/XI0/NET33_XI36/XI0/MM4_d N_XI36/XI0/NET34_XI36/XI0/MM4_g
+ N_VDD_XI36/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI0/MM10 N_XI36/XI0/NET35_XI36/XI0/MM10_d N_XI36/XI0/NET36_XI36/XI0/MM10_g
+ N_VDD_XI36/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI0/MM11 N_XI36/XI0/NET36_XI36/XI0/MM11_d N_XI36/XI0/NET35_XI36/XI0/MM11_g
+ N_VDD_XI36/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI1/MM2 N_XI36/XI1/NET34_XI36/XI1/MM2_d N_XI36/XI1/NET33_XI36/XI1/MM2_g
+ N_VSS_XI36/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI1/MM3 N_XI36/XI1/NET33_XI36/XI1/MM3_d N_WL<68>_XI36/XI1/MM3_g
+ N_BLN<14>_XI36/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI1/MM0 N_XI36/XI1/NET34_XI36/XI1/MM0_d N_WL<68>_XI36/XI1/MM0_g
+ N_BL<14>_XI36/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI1/MM1 N_XI36/XI1/NET33_XI36/XI1/MM1_d N_XI36/XI1/NET34_XI36/XI1/MM1_g
+ N_VSS_XI36/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI1/MM9 N_XI36/XI1/NET36_XI36/XI1/MM9_d N_WL<69>_XI36/XI1/MM9_g
+ N_BL<14>_XI36/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI1/MM6 N_XI36/XI1/NET35_XI36/XI1/MM6_d N_XI36/XI1/NET36_XI36/XI1/MM6_g
+ N_VSS_XI36/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI1/MM7 N_XI36/XI1/NET36_XI36/XI1/MM7_d N_XI36/XI1/NET35_XI36/XI1/MM7_g
+ N_VSS_XI36/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI1/MM8 N_XI36/XI1/NET35_XI36/XI1/MM8_d N_WL<69>_XI36/XI1/MM8_g
+ N_BLN<14>_XI36/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI1/MM5 N_XI36/XI1/NET34_XI36/XI1/MM5_d N_XI36/XI1/NET33_XI36/XI1/MM5_g
+ N_VDD_XI36/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI1/MM4 N_XI36/XI1/NET33_XI36/XI1/MM4_d N_XI36/XI1/NET34_XI36/XI1/MM4_g
+ N_VDD_XI36/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI1/MM10 N_XI36/XI1/NET35_XI36/XI1/MM10_d N_XI36/XI1/NET36_XI36/XI1/MM10_g
+ N_VDD_XI36/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI1/MM11 N_XI36/XI1/NET36_XI36/XI1/MM11_d N_XI36/XI1/NET35_XI36/XI1/MM11_g
+ N_VDD_XI36/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI2/MM2 N_XI36/XI2/NET34_XI36/XI2/MM2_d N_XI36/XI2/NET33_XI36/XI2/MM2_g
+ N_VSS_XI36/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI2/MM3 N_XI36/XI2/NET33_XI36/XI2/MM3_d N_WL<68>_XI36/XI2/MM3_g
+ N_BLN<13>_XI36/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI2/MM0 N_XI36/XI2/NET34_XI36/XI2/MM0_d N_WL<68>_XI36/XI2/MM0_g
+ N_BL<13>_XI36/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI2/MM1 N_XI36/XI2/NET33_XI36/XI2/MM1_d N_XI36/XI2/NET34_XI36/XI2/MM1_g
+ N_VSS_XI36/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI2/MM9 N_XI36/XI2/NET36_XI36/XI2/MM9_d N_WL<69>_XI36/XI2/MM9_g
+ N_BL<13>_XI36/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI2/MM6 N_XI36/XI2/NET35_XI36/XI2/MM6_d N_XI36/XI2/NET36_XI36/XI2/MM6_g
+ N_VSS_XI36/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI2/MM7 N_XI36/XI2/NET36_XI36/XI2/MM7_d N_XI36/XI2/NET35_XI36/XI2/MM7_g
+ N_VSS_XI36/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI2/MM8 N_XI36/XI2/NET35_XI36/XI2/MM8_d N_WL<69>_XI36/XI2/MM8_g
+ N_BLN<13>_XI36/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI2/MM5 N_XI36/XI2/NET34_XI36/XI2/MM5_d N_XI36/XI2/NET33_XI36/XI2/MM5_g
+ N_VDD_XI36/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI2/MM4 N_XI36/XI2/NET33_XI36/XI2/MM4_d N_XI36/XI2/NET34_XI36/XI2/MM4_g
+ N_VDD_XI36/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI2/MM10 N_XI36/XI2/NET35_XI36/XI2/MM10_d N_XI36/XI2/NET36_XI36/XI2/MM10_g
+ N_VDD_XI36/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI2/MM11 N_XI36/XI2/NET36_XI36/XI2/MM11_d N_XI36/XI2/NET35_XI36/XI2/MM11_g
+ N_VDD_XI36/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI3/MM2 N_XI36/XI3/NET34_XI36/XI3/MM2_d N_XI36/XI3/NET33_XI36/XI3/MM2_g
+ N_VSS_XI36/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI3/MM3 N_XI36/XI3/NET33_XI36/XI3/MM3_d N_WL<68>_XI36/XI3/MM3_g
+ N_BLN<12>_XI36/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI3/MM0 N_XI36/XI3/NET34_XI36/XI3/MM0_d N_WL<68>_XI36/XI3/MM0_g
+ N_BL<12>_XI36/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI3/MM1 N_XI36/XI3/NET33_XI36/XI3/MM1_d N_XI36/XI3/NET34_XI36/XI3/MM1_g
+ N_VSS_XI36/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI3/MM9 N_XI36/XI3/NET36_XI36/XI3/MM9_d N_WL<69>_XI36/XI3/MM9_g
+ N_BL<12>_XI36/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI3/MM6 N_XI36/XI3/NET35_XI36/XI3/MM6_d N_XI36/XI3/NET36_XI36/XI3/MM6_g
+ N_VSS_XI36/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI3/MM7 N_XI36/XI3/NET36_XI36/XI3/MM7_d N_XI36/XI3/NET35_XI36/XI3/MM7_g
+ N_VSS_XI36/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI3/MM8 N_XI36/XI3/NET35_XI36/XI3/MM8_d N_WL<69>_XI36/XI3/MM8_g
+ N_BLN<12>_XI36/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI3/MM5 N_XI36/XI3/NET34_XI36/XI3/MM5_d N_XI36/XI3/NET33_XI36/XI3/MM5_g
+ N_VDD_XI36/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI3/MM4 N_XI36/XI3/NET33_XI36/XI3/MM4_d N_XI36/XI3/NET34_XI36/XI3/MM4_g
+ N_VDD_XI36/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI3/MM10 N_XI36/XI3/NET35_XI36/XI3/MM10_d N_XI36/XI3/NET36_XI36/XI3/MM10_g
+ N_VDD_XI36/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI3/MM11 N_XI36/XI3/NET36_XI36/XI3/MM11_d N_XI36/XI3/NET35_XI36/XI3/MM11_g
+ N_VDD_XI36/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI4/MM2 N_XI36/XI4/NET34_XI36/XI4/MM2_d N_XI36/XI4/NET33_XI36/XI4/MM2_g
+ N_VSS_XI36/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI4/MM3 N_XI36/XI4/NET33_XI36/XI4/MM3_d N_WL<68>_XI36/XI4/MM3_g
+ N_BLN<11>_XI36/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI4/MM0 N_XI36/XI4/NET34_XI36/XI4/MM0_d N_WL<68>_XI36/XI4/MM0_g
+ N_BL<11>_XI36/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI4/MM1 N_XI36/XI4/NET33_XI36/XI4/MM1_d N_XI36/XI4/NET34_XI36/XI4/MM1_g
+ N_VSS_XI36/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI4/MM9 N_XI36/XI4/NET36_XI36/XI4/MM9_d N_WL<69>_XI36/XI4/MM9_g
+ N_BL<11>_XI36/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI4/MM6 N_XI36/XI4/NET35_XI36/XI4/MM6_d N_XI36/XI4/NET36_XI36/XI4/MM6_g
+ N_VSS_XI36/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI4/MM7 N_XI36/XI4/NET36_XI36/XI4/MM7_d N_XI36/XI4/NET35_XI36/XI4/MM7_g
+ N_VSS_XI36/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI4/MM8 N_XI36/XI4/NET35_XI36/XI4/MM8_d N_WL<69>_XI36/XI4/MM8_g
+ N_BLN<11>_XI36/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI4/MM5 N_XI36/XI4/NET34_XI36/XI4/MM5_d N_XI36/XI4/NET33_XI36/XI4/MM5_g
+ N_VDD_XI36/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI4/MM4 N_XI36/XI4/NET33_XI36/XI4/MM4_d N_XI36/XI4/NET34_XI36/XI4/MM4_g
+ N_VDD_XI36/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI4/MM10 N_XI36/XI4/NET35_XI36/XI4/MM10_d N_XI36/XI4/NET36_XI36/XI4/MM10_g
+ N_VDD_XI36/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI4/MM11 N_XI36/XI4/NET36_XI36/XI4/MM11_d N_XI36/XI4/NET35_XI36/XI4/MM11_g
+ N_VDD_XI36/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI5/MM2 N_XI36/XI5/NET34_XI36/XI5/MM2_d N_XI36/XI5/NET33_XI36/XI5/MM2_g
+ N_VSS_XI36/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI5/MM3 N_XI36/XI5/NET33_XI36/XI5/MM3_d N_WL<68>_XI36/XI5/MM3_g
+ N_BLN<10>_XI36/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI5/MM0 N_XI36/XI5/NET34_XI36/XI5/MM0_d N_WL<68>_XI36/XI5/MM0_g
+ N_BL<10>_XI36/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI5/MM1 N_XI36/XI5/NET33_XI36/XI5/MM1_d N_XI36/XI5/NET34_XI36/XI5/MM1_g
+ N_VSS_XI36/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI5/MM9 N_XI36/XI5/NET36_XI36/XI5/MM9_d N_WL<69>_XI36/XI5/MM9_g
+ N_BL<10>_XI36/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI5/MM6 N_XI36/XI5/NET35_XI36/XI5/MM6_d N_XI36/XI5/NET36_XI36/XI5/MM6_g
+ N_VSS_XI36/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI5/MM7 N_XI36/XI5/NET36_XI36/XI5/MM7_d N_XI36/XI5/NET35_XI36/XI5/MM7_g
+ N_VSS_XI36/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI5/MM8 N_XI36/XI5/NET35_XI36/XI5/MM8_d N_WL<69>_XI36/XI5/MM8_g
+ N_BLN<10>_XI36/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI5/MM5 N_XI36/XI5/NET34_XI36/XI5/MM5_d N_XI36/XI5/NET33_XI36/XI5/MM5_g
+ N_VDD_XI36/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI5/MM4 N_XI36/XI5/NET33_XI36/XI5/MM4_d N_XI36/XI5/NET34_XI36/XI5/MM4_g
+ N_VDD_XI36/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI5/MM10 N_XI36/XI5/NET35_XI36/XI5/MM10_d N_XI36/XI5/NET36_XI36/XI5/MM10_g
+ N_VDD_XI36/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI5/MM11 N_XI36/XI5/NET36_XI36/XI5/MM11_d N_XI36/XI5/NET35_XI36/XI5/MM11_g
+ N_VDD_XI36/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI6/MM2 N_XI36/XI6/NET34_XI36/XI6/MM2_d N_XI36/XI6/NET33_XI36/XI6/MM2_g
+ N_VSS_XI36/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM3 N_XI36/XI6/NET33_XI36/XI6/MM3_d N_WL<68>_XI36/XI6/MM3_g
+ N_BLN<9>_XI36/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM0 N_XI36/XI6/NET34_XI36/XI6/MM0_d N_WL<68>_XI36/XI6/MM0_g
+ N_BL<9>_XI36/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM1 N_XI36/XI6/NET33_XI36/XI6/MM1_d N_XI36/XI6/NET34_XI36/XI6/MM1_g
+ N_VSS_XI36/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM9 N_XI36/XI6/NET36_XI36/XI6/MM9_d N_WL<69>_XI36/XI6/MM9_g
+ N_BL<9>_XI36/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM6 N_XI36/XI6/NET35_XI36/XI6/MM6_d N_XI36/XI6/NET36_XI36/XI6/MM6_g
+ N_VSS_XI36/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM7 N_XI36/XI6/NET36_XI36/XI6/MM7_d N_XI36/XI6/NET35_XI36/XI6/MM7_g
+ N_VSS_XI36/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM8 N_XI36/XI6/NET35_XI36/XI6/MM8_d N_WL<69>_XI36/XI6/MM8_g
+ N_BLN<9>_XI36/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI6/MM5 N_XI36/XI6/NET34_XI36/XI6/MM5_d N_XI36/XI6/NET33_XI36/XI6/MM5_g
+ N_VDD_XI36/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI6/MM4 N_XI36/XI6/NET33_XI36/XI6/MM4_d N_XI36/XI6/NET34_XI36/XI6/MM4_g
+ N_VDD_XI36/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI6/MM10 N_XI36/XI6/NET35_XI36/XI6/MM10_d N_XI36/XI6/NET36_XI36/XI6/MM10_g
+ N_VDD_XI36/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI6/MM11 N_XI36/XI6/NET36_XI36/XI6/MM11_d N_XI36/XI6/NET35_XI36/XI6/MM11_g
+ N_VDD_XI36/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI7/MM2 N_XI36/XI7/NET34_XI36/XI7/MM2_d N_XI36/XI7/NET33_XI36/XI7/MM2_g
+ N_VSS_XI36/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM3 N_XI36/XI7/NET33_XI36/XI7/MM3_d N_WL<68>_XI36/XI7/MM3_g
+ N_BLN<8>_XI36/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM0 N_XI36/XI7/NET34_XI36/XI7/MM0_d N_WL<68>_XI36/XI7/MM0_g
+ N_BL<8>_XI36/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM1 N_XI36/XI7/NET33_XI36/XI7/MM1_d N_XI36/XI7/NET34_XI36/XI7/MM1_g
+ N_VSS_XI36/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM9 N_XI36/XI7/NET36_XI36/XI7/MM9_d N_WL<69>_XI36/XI7/MM9_g
+ N_BL<8>_XI36/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM6 N_XI36/XI7/NET35_XI36/XI7/MM6_d N_XI36/XI7/NET36_XI36/XI7/MM6_g
+ N_VSS_XI36/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM7 N_XI36/XI7/NET36_XI36/XI7/MM7_d N_XI36/XI7/NET35_XI36/XI7/MM7_g
+ N_VSS_XI36/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM8 N_XI36/XI7/NET35_XI36/XI7/MM8_d N_WL<69>_XI36/XI7/MM8_g
+ N_BLN<8>_XI36/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI7/MM5 N_XI36/XI7/NET34_XI36/XI7/MM5_d N_XI36/XI7/NET33_XI36/XI7/MM5_g
+ N_VDD_XI36/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI7/MM4 N_XI36/XI7/NET33_XI36/XI7/MM4_d N_XI36/XI7/NET34_XI36/XI7/MM4_g
+ N_VDD_XI36/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI7/MM10 N_XI36/XI7/NET35_XI36/XI7/MM10_d N_XI36/XI7/NET36_XI36/XI7/MM10_g
+ N_VDD_XI36/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI7/MM11 N_XI36/XI7/NET36_XI36/XI7/MM11_d N_XI36/XI7/NET35_XI36/XI7/MM11_g
+ N_VDD_XI36/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI8/MM2 N_XI36/XI8/NET34_XI36/XI8/MM2_d N_XI36/XI8/NET33_XI36/XI8/MM2_g
+ N_VSS_XI36/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM3 N_XI36/XI8/NET33_XI36/XI8/MM3_d N_WL<68>_XI36/XI8/MM3_g
+ N_BLN<7>_XI36/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM0 N_XI36/XI8/NET34_XI36/XI8/MM0_d N_WL<68>_XI36/XI8/MM0_g
+ N_BL<7>_XI36/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM1 N_XI36/XI8/NET33_XI36/XI8/MM1_d N_XI36/XI8/NET34_XI36/XI8/MM1_g
+ N_VSS_XI36/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM9 N_XI36/XI8/NET36_XI36/XI8/MM9_d N_WL<69>_XI36/XI8/MM9_g
+ N_BL<7>_XI36/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM6 N_XI36/XI8/NET35_XI36/XI8/MM6_d N_XI36/XI8/NET36_XI36/XI8/MM6_g
+ N_VSS_XI36/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM7 N_XI36/XI8/NET36_XI36/XI8/MM7_d N_XI36/XI8/NET35_XI36/XI8/MM7_g
+ N_VSS_XI36/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM8 N_XI36/XI8/NET35_XI36/XI8/MM8_d N_WL<69>_XI36/XI8/MM8_g
+ N_BLN<7>_XI36/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI8/MM5 N_XI36/XI8/NET34_XI36/XI8/MM5_d N_XI36/XI8/NET33_XI36/XI8/MM5_g
+ N_VDD_XI36/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI8/MM4 N_XI36/XI8/NET33_XI36/XI8/MM4_d N_XI36/XI8/NET34_XI36/XI8/MM4_g
+ N_VDD_XI36/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI8/MM10 N_XI36/XI8/NET35_XI36/XI8/MM10_d N_XI36/XI8/NET36_XI36/XI8/MM10_g
+ N_VDD_XI36/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI8/MM11 N_XI36/XI8/NET36_XI36/XI8/MM11_d N_XI36/XI8/NET35_XI36/XI8/MM11_g
+ N_VDD_XI36/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI9/MM2 N_XI36/XI9/NET34_XI36/XI9/MM2_d N_XI36/XI9/NET33_XI36/XI9/MM2_g
+ N_VSS_XI36/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM3 N_XI36/XI9/NET33_XI36/XI9/MM3_d N_WL<68>_XI36/XI9/MM3_g
+ N_BLN<6>_XI36/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM0 N_XI36/XI9/NET34_XI36/XI9/MM0_d N_WL<68>_XI36/XI9/MM0_g
+ N_BL<6>_XI36/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM1 N_XI36/XI9/NET33_XI36/XI9/MM1_d N_XI36/XI9/NET34_XI36/XI9/MM1_g
+ N_VSS_XI36/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM9 N_XI36/XI9/NET36_XI36/XI9/MM9_d N_WL<69>_XI36/XI9/MM9_g
+ N_BL<6>_XI36/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM6 N_XI36/XI9/NET35_XI36/XI9/MM6_d N_XI36/XI9/NET36_XI36/XI9/MM6_g
+ N_VSS_XI36/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM7 N_XI36/XI9/NET36_XI36/XI9/MM7_d N_XI36/XI9/NET35_XI36/XI9/MM7_g
+ N_VSS_XI36/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM8 N_XI36/XI9/NET35_XI36/XI9/MM8_d N_WL<69>_XI36/XI9/MM8_g
+ N_BLN<6>_XI36/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI9/MM5 N_XI36/XI9/NET34_XI36/XI9/MM5_d N_XI36/XI9/NET33_XI36/XI9/MM5_g
+ N_VDD_XI36/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI9/MM4 N_XI36/XI9/NET33_XI36/XI9/MM4_d N_XI36/XI9/NET34_XI36/XI9/MM4_g
+ N_VDD_XI36/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI9/MM10 N_XI36/XI9/NET35_XI36/XI9/MM10_d N_XI36/XI9/NET36_XI36/XI9/MM10_g
+ N_VDD_XI36/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI9/MM11 N_XI36/XI9/NET36_XI36/XI9/MM11_d N_XI36/XI9/NET35_XI36/XI9/MM11_g
+ N_VDD_XI36/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI10/MM2 N_XI36/XI10/NET34_XI36/XI10/MM2_d
+ N_XI36/XI10/NET33_XI36/XI10/MM2_g N_VSS_XI36/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI10/MM3 N_XI36/XI10/NET33_XI36/XI10/MM3_d N_WL<68>_XI36/XI10/MM3_g
+ N_BLN<5>_XI36/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI10/MM0 N_XI36/XI10/NET34_XI36/XI10/MM0_d N_WL<68>_XI36/XI10/MM0_g
+ N_BL<5>_XI36/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI10/MM1 N_XI36/XI10/NET33_XI36/XI10/MM1_d
+ N_XI36/XI10/NET34_XI36/XI10/MM1_g N_VSS_XI36/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI10/MM9 N_XI36/XI10/NET36_XI36/XI10/MM9_d N_WL<69>_XI36/XI10/MM9_g
+ N_BL<5>_XI36/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI10/MM6 N_XI36/XI10/NET35_XI36/XI10/MM6_d
+ N_XI36/XI10/NET36_XI36/XI10/MM6_g N_VSS_XI36/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI10/MM7 N_XI36/XI10/NET36_XI36/XI10/MM7_d
+ N_XI36/XI10/NET35_XI36/XI10/MM7_g N_VSS_XI36/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI10/MM8 N_XI36/XI10/NET35_XI36/XI10/MM8_d N_WL<69>_XI36/XI10/MM8_g
+ N_BLN<5>_XI36/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI10/MM5 N_XI36/XI10/NET34_XI36/XI10/MM5_d
+ N_XI36/XI10/NET33_XI36/XI10/MM5_g N_VDD_XI36/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI10/MM4 N_XI36/XI10/NET33_XI36/XI10/MM4_d
+ N_XI36/XI10/NET34_XI36/XI10/MM4_g N_VDD_XI36/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI10/MM10 N_XI36/XI10/NET35_XI36/XI10/MM10_d
+ N_XI36/XI10/NET36_XI36/XI10/MM10_g N_VDD_XI36/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI10/MM11 N_XI36/XI10/NET36_XI36/XI10/MM11_d
+ N_XI36/XI10/NET35_XI36/XI10/MM11_g N_VDD_XI36/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI11/MM2 N_XI36/XI11/NET34_XI36/XI11/MM2_d
+ N_XI36/XI11/NET33_XI36/XI11/MM2_g N_VSS_XI36/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI11/MM3 N_XI36/XI11/NET33_XI36/XI11/MM3_d N_WL<68>_XI36/XI11/MM3_g
+ N_BLN<4>_XI36/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI11/MM0 N_XI36/XI11/NET34_XI36/XI11/MM0_d N_WL<68>_XI36/XI11/MM0_g
+ N_BL<4>_XI36/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI11/MM1 N_XI36/XI11/NET33_XI36/XI11/MM1_d
+ N_XI36/XI11/NET34_XI36/XI11/MM1_g N_VSS_XI36/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI11/MM9 N_XI36/XI11/NET36_XI36/XI11/MM9_d N_WL<69>_XI36/XI11/MM9_g
+ N_BL<4>_XI36/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI11/MM6 N_XI36/XI11/NET35_XI36/XI11/MM6_d
+ N_XI36/XI11/NET36_XI36/XI11/MM6_g N_VSS_XI36/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI11/MM7 N_XI36/XI11/NET36_XI36/XI11/MM7_d
+ N_XI36/XI11/NET35_XI36/XI11/MM7_g N_VSS_XI36/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI11/MM8 N_XI36/XI11/NET35_XI36/XI11/MM8_d N_WL<69>_XI36/XI11/MM8_g
+ N_BLN<4>_XI36/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI11/MM5 N_XI36/XI11/NET34_XI36/XI11/MM5_d
+ N_XI36/XI11/NET33_XI36/XI11/MM5_g N_VDD_XI36/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI11/MM4 N_XI36/XI11/NET33_XI36/XI11/MM4_d
+ N_XI36/XI11/NET34_XI36/XI11/MM4_g N_VDD_XI36/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI11/MM10 N_XI36/XI11/NET35_XI36/XI11/MM10_d
+ N_XI36/XI11/NET36_XI36/XI11/MM10_g N_VDD_XI36/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI11/MM11 N_XI36/XI11/NET36_XI36/XI11/MM11_d
+ N_XI36/XI11/NET35_XI36/XI11/MM11_g N_VDD_XI36/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI12/MM2 N_XI36/XI12/NET34_XI36/XI12/MM2_d
+ N_XI36/XI12/NET33_XI36/XI12/MM2_g N_VSS_XI36/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI12/MM3 N_XI36/XI12/NET33_XI36/XI12/MM3_d N_WL<68>_XI36/XI12/MM3_g
+ N_BLN<3>_XI36/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI12/MM0 N_XI36/XI12/NET34_XI36/XI12/MM0_d N_WL<68>_XI36/XI12/MM0_g
+ N_BL<3>_XI36/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI12/MM1 N_XI36/XI12/NET33_XI36/XI12/MM1_d
+ N_XI36/XI12/NET34_XI36/XI12/MM1_g N_VSS_XI36/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI12/MM9 N_XI36/XI12/NET36_XI36/XI12/MM9_d N_WL<69>_XI36/XI12/MM9_g
+ N_BL<3>_XI36/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI12/MM6 N_XI36/XI12/NET35_XI36/XI12/MM6_d
+ N_XI36/XI12/NET36_XI36/XI12/MM6_g N_VSS_XI36/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI12/MM7 N_XI36/XI12/NET36_XI36/XI12/MM7_d
+ N_XI36/XI12/NET35_XI36/XI12/MM7_g N_VSS_XI36/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI12/MM8 N_XI36/XI12/NET35_XI36/XI12/MM8_d N_WL<69>_XI36/XI12/MM8_g
+ N_BLN<3>_XI36/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI12/MM5 N_XI36/XI12/NET34_XI36/XI12/MM5_d
+ N_XI36/XI12/NET33_XI36/XI12/MM5_g N_VDD_XI36/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI12/MM4 N_XI36/XI12/NET33_XI36/XI12/MM4_d
+ N_XI36/XI12/NET34_XI36/XI12/MM4_g N_VDD_XI36/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI12/MM10 N_XI36/XI12/NET35_XI36/XI12/MM10_d
+ N_XI36/XI12/NET36_XI36/XI12/MM10_g N_VDD_XI36/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI12/MM11 N_XI36/XI12/NET36_XI36/XI12/MM11_d
+ N_XI36/XI12/NET35_XI36/XI12/MM11_g N_VDD_XI36/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI13/MM2 N_XI36/XI13/NET34_XI36/XI13/MM2_d
+ N_XI36/XI13/NET33_XI36/XI13/MM2_g N_VSS_XI36/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI13/MM3 N_XI36/XI13/NET33_XI36/XI13/MM3_d N_WL<68>_XI36/XI13/MM3_g
+ N_BLN<2>_XI36/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI13/MM0 N_XI36/XI13/NET34_XI36/XI13/MM0_d N_WL<68>_XI36/XI13/MM0_g
+ N_BL<2>_XI36/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI13/MM1 N_XI36/XI13/NET33_XI36/XI13/MM1_d
+ N_XI36/XI13/NET34_XI36/XI13/MM1_g N_VSS_XI36/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI13/MM9 N_XI36/XI13/NET36_XI36/XI13/MM9_d N_WL<69>_XI36/XI13/MM9_g
+ N_BL<2>_XI36/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI13/MM6 N_XI36/XI13/NET35_XI36/XI13/MM6_d
+ N_XI36/XI13/NET36_XI36/XI13/MM6_g N_VSS_XI36/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI13/MM7 N_XI36/XI13/NET36_XI36/XI13/MM7_d
+ N_XI36/XI13/NET35_XI36/XI13/MM7_g N_VSS_XI36/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI13/MM8 N_XI36/XI13/NET35_XI36/XI13/MM8_d N_WL<69>_XI36/XI13/MM8_g
+ N_BLN<2>_XI36/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI13/MM5 N_XI36/XI13/NET34_XI36/XI13/MM5_d
+ N_XI36/XI13/NET33_XI36/XI13/MM5_g N_VDD_XI36/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI13/MM4 N_XI36/XI13/NET33_XI36/XI13/MM4_d
+ N_XI36/XI13/NET34_XI36/XI13/MM4_g N_VDD_XI36/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI13/MM10 N_XI36/XI13/NET35_XI36/XI13/MM10_d
+ N_XI36/XI13/NET36_XI36/XI13/MM10_g N_VDD_XI36/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI13/MM11 N_XI36/XI13/NET36_XI36/XI13/MM11_d
+ N_XI36/XI13/NET35_XI36/XI13/MM11_g N_VDD_XI36/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI14/MM2 N_XI36/XI14/NET34_XI36/XI14/MM2_d
+ N_XI36/XI14/NET33_XI36/XI14/MM2_g N_VSS_XI36/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI14/MM3 N_XI36/XI14/NET33_XI36/XI14/MM3_d N_WL<68>_XI36/XI14/MM3_g
+ N_BLN<1>_XI36/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI14/MM0 N_XI36/XI14/NET34_XI36/XI14/MM0_d N_WL<68>_XI36/XI14/MM0_g
+ N_BL<1>_XI36/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI14/MM1 N_XI36/XI14/NET33_XI36/XI14/MM1_d
+ N_XI36/XI14/NET34_XI36/XI14/MM1_g N_VSS_XI36/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI14/MM9 N_XI36/XI14/NET36_XI36/XI14/MM9_d N_WL<69>_XI36/XI14/MM9_g
+ N_BL<1>_XI36/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI14/MM6 N_XI36/XI14/NET35_XI36/XI14/MM6_d
+ N_XI36/XI14/NET36_XI36/XI14/MM6_g N_VSS_XI36/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI14/MM7 N_XI36/XI14/NET36_XI36/XI14/MM7_d
+ N_XI36/XI14/NET35_XI36/XI14/MM7_g N_VSS_XI36/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI14/MM8 N_XI36/XI14/NET35_XI36/XI14/MM8_d N_WL<69>_XI36/XI14/MM8_g
+ N_BLN<1>_XI36/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI14/MM5 N_XI36/XI14/NET34_XI36/XI14/MM5_d
+ N_XI36/XI14/NET33_XI36/XI14/MM5_g N_VDD_XI36/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI14/MM4 N_XI36/XI14/NET33_XI36/XI14/MM4_d
+ N_XI36/XI14/NET34_XI36/XI14/MM4_g N_VDD_XI36/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI14/MM10 N_XI36/XI14/NET35_XI36/XI14/MM10_d
+ N_XI36/XI14/NET36_XI36/XI14/MM10_g N_VDD_XI36/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI14/MM11 N_XI36/XI14/NET36_XI36/XI14/MM11_d
+ N_XI36/XI14/NET35_XI36/XI14/MM11_g N_VDD_XI36/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI15/MM2 N_XI36/XI15/NET34_XI36/XI15/MM2_d
+ N_XI36/XI15/NET33_XI36/XI15/MM2_g N_VSS_XI36/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI15/MM3 N_XI36/XI15/NET33_XI36/XI15/MM3_d N_WL<68>_XI36/XI15/MM3_g
+ N_BLN<0>_XI36/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI15/MM0 N_XI36/XI15/NET34_XI36/XI15/MM0_d N_WL<68>_XI36/XI15/MM0_g
+ N_BL<0>_XI36/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI15/MM1 N_XI36/XI15/NET33_XI36/XI15/MM1_d
+ N_XI36/XI15/NET34_XI36/XI15/MM1_g N_VSS_XI36/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI15/MM9 N_XI36/XI15/NET36_XI36/XI15/MM9_d N_WL<69>_XI36/XI15/MM9_g
+ N_BL<0>_XI36/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI15/MM6 N_XI36/XI15/NET35_XI36/XI15/MM6_d
+ N_XI36/XI15/NET36_XI36/XI15/MM6_g N_VSS_XI36/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI15/MM7 N_XI36/XI15/NET36_XI36/XI15/MM7_d
+ N_XI36/XI15/NET35_XI36/XI15/MM7_g N_VSS_XI36/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI36/XI15/MM8 N_XI36/XI15/NET35_XI36/XI15/MM8_d N_WL<69>_XI36/XI15/MM8_g
+ N_BLN<0>_XI36/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI36/XI15/MM5 N_XI36/XI15/NET34_XI36/XI15/MM5_d
+ N_XI36/XI15/NET33_XI36/XI15/MM5_g N_VDD_XI36/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI15/MM4 N_XI36/XI15/NET33_XI36/XI15/MM4_d
+ N_XI36/XI15/NET34_XI36/XI15/MM4_g N_VDD_XI36/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI15/MM10 N_XI36/XI15/NET35_XI36/XI15/MM10_d
+ N_XI36/XI15/NET36_XI36/XI15/MM10_g N_VDD_XI36/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI36/XI15/MM11 N_XI36/XI15/NET36_XI36/XI15/MM11_d
+ N_XI36/XI15/NET35_XI36/XI15/MM11_g N_VDD_XI36/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI0/MM2 N_XI37/XI0/NET34_XI37/XI0/MM2_d N_XI37/XI0/NET33_XI37/XI0/MM2_g
+ N_VSS_XI37/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI0/MM3 N_XI37/XI0/NET33_XI37/XI0/MM3_d N_WL<70>_XI37/XI0/MM3_g
+ N_BLN<15>_XI37/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI0/MM0 N_XI37/XI0/NET34_XI37/XI0/MM0_d N_WL<70>_XI37/XI0/MM0_g
+ N_BL<15>_XI37/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI0/MM1 N_XI37/XI0/NET33_XI37/XI0/MM1_d N_XI37/XI0/NET34_XI37/XI0/MM1_g
+ N_VSS_XI37/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI0/MM9 N_XI37/XI0/NET36_XI37/XI0/MM9_d N_WL<71>_XI37/XI0/MM9_g
+ N_BL<15>_XI37/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI0/MM6 N_XI37/XI0/NET35_XI37/XI0/MM6_d N_XI37/XI0/NET36_XI37/XI0/MM6_g
+ N_VSS_XI37/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI0/MM7 N_XI37/XI0/NET36_XI37/XI0/MM7_d N_XI37/XI0/NET35_XI37/XI0/MM7_g
+ N_VSS_XI37/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI0/MM8 N_XI37/XI0/NET35_XI37/XI0/MM8_d N_WL<71>_XI37/XI0/MM8_g
+ N_BLN<15>_XI37/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI0/MM5 N_XI37/XI0/NET34_XI37/XI0/MM5_d N_XI37/XI0/NET33_XI37/XI0/MM5_g
+ N_VDD_XI37/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI0/MM4 N_XI37/XI0/NET33_XI37/XI0/MM4_d N_XI37/XI0/NET34_XI37/XI0/MM4_g
+ N_VDD_XI37/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI0/MM10 N_XI37/XI0/NET35_XI37/XI0/MM10_d N_XI37/XI0/NET36_XI37/XI0/MM10_g
+ N_VDD_XI37/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI0/MM11 N_XI37/XI0/NET36_XI37/XI0/MM11_d N_XI37/XI0/NET35_XI37/XI0/MM11_g
+ N_VDD_XI37/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI1/MM2 N_XI37/XI1/NET34_XI37/XI1/MM2_d N_XI37/XI1/NET33_XI37/XI1/MM2_g
+ N_VSS_XI37/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI1/MM3 N_XI37/XI1/NET33_XI37/XI1/MM3_d N_WL<70>_XI37/XI1/MM3_g
+ N_BLN<14>_XI37/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI1/MM0 N_XI37/XI1/NET34_XI37/XI1/MM0_d N_WL<70>_XI37/XI1/MM0_g
+ N_BL<14>_XI37/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI1/MM1 N_XI37/XI1/NET33_XI37/XI1/MM1_d N_XI37/XI1/NET34_XI37/XI1/MM1_g
+ N_VSS_XI37/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI1/MM9 N_XI37/XI1/NET36_XI37/XI1/MM9_d N_WL<71>_XI37/XI1/MM9_g
+ N_BL<14>_XI37/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI1/MM6 N_XI37/XI1/NET35_XI37/XI1/MM6_d N_XI37/XI1/NET36_XI37/XI1/MM6_g
+ N_VSS_XI37/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI1/MM7 N_XI37/XI1/NET36_XI37/XI1/MM7_d N_XI37/XI1/NET35_XI37/XI1/MM7_g
+ N_VSS_XI37/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI1/MM8 N_XI37/XI1/NET35_XI37/XI1/MM8_d N_WL<71>_XI37/XI1/MM8_g
+ N_BLN<14>_XI37/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI1/MM5 N_XI37/XI1/NET34_XI37/XI1/MM5_d N_XI37/XI1/NET33_XI37/XI1/MM5_g
+ N_VDD_XI37/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI1/MM4 N_XI37/XI1/NET33_XI37/XI1/MM4_d N_XI37/XI1/NET34_XI37/XI1/MM4_g
+ N_VDD_XI37/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI1/MM10 N_XI37/XI1/NET35_XI37/XI1/MM10_d N_XI37/XI1/NET36_XI37/XI1/MM10_g
+ N_VDD_XI37/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI1/MM11 N_XI37/XI1/NET36_XI37/XI1/MM11_d N_XI37/XI1/NET35_XI37/XI1/MM11_g
+ N_VDD_XI37/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI2/MM2 N_XI37/XI2/NET34_XI37/XI2/MM2_d N_XI37/XI2/NET33_XI37/XI2/MM2_g
+ N_VSS_XI37/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI2/MM3 N_XI37/XI2/NET33_XI37/XI2/MM3_d N_WL<70>_XI37/XI2/MM3_g
+ N_BLN<13>_XI37/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI2/MM0 N_XI37/XI2/NET34_XI37/XI2/MM0_d N_WL<70>_XI37/XI2/MM0_g
+ N_BL<13>_XI37/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI2/MM1 N_XI37/XI2/NET33_XI37/XI2/MM1_d N_XI37/XI2/NET34_XI37/XI2/MM1_g
+ N_VSS_XI37/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI2/MM9 N_XI37/XI2/NET36_XI37/XI2/MM9_d N_WL<71>_XI37/XI2/MM9_g
+ N_BL<13>_XI37/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI2/MM6 N_XI37/XI2/NET35_XI37/XI2/MM6_d N_XI37/XI2/NET36_XI37/XI2/MM6_g
+ N_VSS_XI37/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI2/MM7 N_XI37/XI2/NET36_XI37/XI2/MM7_d N_XI37/XI2/NET35_XI37/XI2/MM7_g
+ N_VSS_XI37/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI2/MM8 N_XI37/XI2/NET35_XI37/XI2/MM8_d N_WL<71>_XI37/XI2/MM8_g
+ N_BLN<13>_XI37/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI2/MM5 N_XI37/XI2/NET34_XI37/XI2/MM5_d N_XI37/XI2/NET33_XI37/XI2/MM5_g
+ N_VDD_XI37/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI2/MM4 N_XI37/XI2/NET33_XI37/XI2/MM4_d N_XI37/XI2/NET34_XI37/XI2/MM4_g
+ N_VDD_XI37/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI2/MM10 N_XI37/XI2/NET35_XI37/XI2/MM10_d N_XI37/XI2/NET36_XI37/XI2/MM10_g
+ N_VDD_XI37/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI2/MM11 N_XI37/XI2/NET36_XI37/XI2/MM11_d N_XI37/XI2/NET35_XI37/XI2/MM11_g
+ N_VDD_XI37/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI3/MM2 N_XI37/XI3/NET34_XI37/XI3/MM2_d N_XI37/XI3/NET33_XI37/XI3/MM2_g
+ N_VSS_XI37/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI3/MM3 N_XI37/XI3/NET33_XI37/XI3/MM3_d N_WL<70>_XI37/XI3/MM3_g
+ N_BLN<12>_XI37/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI3/MM0 N_XI37/XI3/NET34_XI37/XI3/MM0_d N_WL<70>_XI37/XI3/MM0_g
+ N_BL<12>_XI37/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI3/MM1 N_XI37/XI3/NET33_XI37/XI3/MM1_d N_XI37/XI3/NET34_XI37/XI3/MM1_g
+ N_VSS_XI37/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI3/MM9 N_XI37/XI3/NET36_XI37/XI3/MM9_d N_WL<71>_XI37/XI3/MM9_g
+ N_BL<12>_XI37/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI3/MM6 N_XI37/XI3/NET35_XI37/XI3/MM6_d N_XI37/XI3/NET36_XI37/XI3/MM6_g
+ N_VSS_XI37/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI3/MM7 N_XI37/XI3/NET36_XI37/XI3/MM7_d N_XI37/XI3/NET35_XI37/XI3/MM7_g
+ N_VSS_XI37/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI3/MM8 N_XI37/XI3/NET35_XI37/XI3/MM8_d N_WL<71>_XI37/XI3/MM8_g
+ N_BLN<12>_XI37/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI3/MM5 N_XI37/XI3/NET34_XI37/XI3/MM5_d N_XI37/XI3/NET33_XI37/XI3/MM5_g
+ N_VDD_XI37/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI3/MM4 N_XI37/XI3/NET33_XI37/XI3/MM4_d N_XI37/XI3/NET34_XI37/XI3/MM4_g
+ N_VDD_XI37/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI3/MM10 N_XI37/XI3/NET35_XI37/XI3/MM10_d N_XI37/XI3/NET36_XI37/XI3/MM10_g
+ N_VDD_XI37/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI3/MM11 N_XI37/XI3/NET36_XI37/XI3/MM11_d N_XI37/XI3/NET35_XI37/XI3/MM11_g
+ N_VDD_XI37/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI4/MM2 N_XI37/XI4/NET34_XI37/XI4/MM2_d N_XI37/XI4/NET33_XI37/XI4/MM2_g
+ N_VSS_XI37/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI4/MM3 N_XI37/XI4/NET33_XI37/XI4/MM3_d N_WL<70>_XI37/XI4/MM3_g
+ N_BLN<11>_XI37/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI4/MM0 N_XI37/XI4/NET34_XI37/XI4/MM0_d N_WL<70>_XI37/XI4/MM0_g
+ N_BL<11>_XI37/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI4/MM1 N_XI37/XI4/NET33_XI37/XI4/MM1_d N_XI37/XI4/NET34_XI37/XI4/MM1_g
+ N_VSS_XI37/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI4/MM9 N_XI37/XI4/NET36_XI37/XI4/MM9_d N_WL<71>_XI37/XI4/MM9_g
+ N_BL<11>_XI37/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI4/MM6 N_XI37/XI4/NET35_XI37/XI4/MM6_d N_XI37/XI4/NET36_XI37/XI4/MM6_g
+ N_VSS_XI37/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI4/MM7 N_XI37/XI4/NET36_XI37/XI4/MM7_d N_XI37/XI4/NET35_XI37/XI4/MM7_g
+ N_VSS_XI37/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI4/MM8 N_XI37/XI4/NET35_XI37/XI4/MM8_d N_WL<71>_XI37/XI4/MM8_g
+ N_BLN<11>_XI37/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI4/MM5 N_XI37/XI4/NET34_XI37/XI4/MM5_d N_XI37/XI4/NET33_XI37/XI4/MM5_g
+ N_VDD_XI37/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI4/MM4 N_XI37/XI4/NET33_XI37/XI4/MM4_d N_XI37/XI4/NET34_XI37/XI4/MM4_g
+ N_VDD_XI37/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI4/MM10 N_XI37/XI4/NET35_XI37/XI4/MM10_d N_XI37/XI4/NET36_XI37/XI4/MM10_g
+ N_VDD_XI37/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI4/MM11 N_XI37/XI4/NET36_XI37/XI4/MM11_d N_XI37/XI4/NET35_XI37/XI4/MM11_g
+ N_VDD_XI37/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI5/MM2 N_XI37/XI5/NET34_XI37/XI5/MM2_d N_XI37/XI5/NET33_XI37/XI5/MM2_g
+ N_VSS_XI37/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI5/MM3 N_XI37/XI5/NET33_XI37/XI5/MM3_d N_WL<70>_XI37/XI5/MM3_g
+ N_BLN<10>_XI37/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI5/MM0 N_XI37/XI5/NET34_XI37/XI5/MM0_d N_WL<70>_XI37/XI5/MM0_g
+ N_BL<10>_XI37/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI5/MM1 N_XI37/XI5/NET33_XI37/XI5/MM1_d N_XI37/XI5/NET34_XI37/XI5/MM1_g
+ N_VSS_XI37/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI5/MM9 N_XI37/XI5/NET36_XI37/XI5/MM9_d N_WL<71>_XI37/XI5/MM9_g
+ N_BL<10>_XI37/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI5/MM6 N_XI37/XI5/NET35_XI37/XI5/MM6_d N_XI37/XI5/NET36_XI37/XI5/MM6_g
+ N_VSS_XI37/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI5/MM7 N_XI37/XI5/NET36_XI37/XI5/MM7_d N_XI37/XI5/NET35_XI37/XI5/MM7_g
+ N_VSS_XI37/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI5/MM8 N_XI37/XI5/NET35_XI37/XI5/MM8_d N_WL<71>_XI37/XI5/MM8_g
+ N_BLN<10>_XI37/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI5/MM5 N_XI37/XI5/NET34_XI37/XI5/MM5_d N_XI37/XI5/NET33_XI37/XI5/MM5_g
+ N_VDD_XI37/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI5/MM4 N_XI37/XI5/NET33_XI37/XI5/MM4_d N_XI37/XI5/NET34_XI37/XI5/MM4_g
+ N_VDD_XI37/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI5/MM10 N_XI37/XI5/NET35_XI37/XI5/MM10_d N_XI37/XI5/NET36_XI37/XI5/MM10_g
+ N_VDD_XI37/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI5/MM11 N_XI37/XI5/NET36_XI37/XI5/MM11_d N_XI37/XI5/NET35_XI37/XI5/MM11_g
+ N_VDD_XI37/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI6/MM2 N_XI37/XI6/NET34_XI37/XI6/MM2_d N_XI37/XI6/NET33_XI37/XI6/MM2_g
+ N_VSS_XI37/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM3 N_XI37/XI6/NET33_XI37/XI6/MM3_d N_WL<70>_XI37/XI6/MM3_g
+ N_BLN<9>_XI37/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM0 N_XI37/XI6/NET34_XI37/XI6/MM0_d N_WL<70>_XI37/XI6/MM0_g
+ N_BL<9>_XI37/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM1 N_XI37/XI6/NET33_XI37/XI6/MM1_d N_XI37/XI6/NET34_XI37/XI6/MM1_g
+ N_VSS_XI37/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM9 N_XI37/XI6/NET36_XI37/XI6/MM9_d N_WL<71>_XI37/XI6/MM9_g
+ N_BL<9>_XI37/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM6 N_XI37/XI6/NET35_XI37/XI6/MM6_d N_XI37/XI6/NET36_XI37/XI6/MM6_g
+ N_VSS_XI37/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM7 N_XI37/XI6/NET36_XI37/XI6/MM7_d N_XI37/XI6/NET35_XI37/XI6/MM7_g
+ N_VSS_XI37/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM8 N_XI37/XI6/NET35_XI37/XI6/MM8_d N_WL<71>_XI37/XI6/MM8_g
+ N_BLN<9>_XI37/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI6/MM5 N_XI37/XI6/NET34_XI37/XI6/MM5_d N_XI37/XI6/NET33_XI37/XI6/MM5_g
+ N_VDD_XI37/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI6/MM4 N_XI37/XI6/NET33_XI37/XI6/MM4_d N_XI37/XI6/NET34_XI37/XI6/MM4_g
+ N_VDD_XI37/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI6/MM10 N_XI37/XI6/NET35_XI37/XI6/MM10_d N_XI37/XI6/NET36_XI37/XI6/MM10_g
+ N_VDD_XI37/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI6/MM11 N_XI37/XI6/NET36_XI37/XI6/MM11_d N_XI37/XI6/NET35_XI37/XI6/MM11_g
+ N_VDD_XI37/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI7/MM2 N_XI37/XI7/NET34_XI37/XI7/MM2_d N_XI37/XI7/NET33_XI37/XI7/MM2_g
+ N_VSS_XI37/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM3 N_XI37/XI7/NET33_XI37/XI7/MM3_d N_WL<70>_XI37/XI7/MM3_g
+ N_BLN<8>_XI37/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM0 N_XI37/XI7/NET34_XI37/XI7/MM0_d N_WL<70>_XI37/XI7/MM0_g
+ N_BL<8>_XI37/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM1 N_XI37/XI7/NET33_XI37/XI7/MM1_d N_XI37/XI7/NET34_XI37/XI7/MM1_g
+ N_VSS_XI37/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM9 N_XI37/XI7/NET36_XI37/XI7/MM9_d N_WL<71>_XI37/XI7/MM9_g
+ N_BL<8>_XI37/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM6 N_XI37/XI7/NET35_XI37/XI7/MM6_d N_XI37/XI7/NET36_XI37/XI7/MM6_g
+ N_VSS_XI37/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM7 N_XI37/XI7/NET36_XI37/XI7/MM7_d N_XI37/XI7/NET35_XI37/XI7/MM7_g
+ N_VSS_XI37/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM8 N_XI37/XI7/NET35_XI37/XI7/MM8_d N_WL<71>_XI37/XI7/MM8_g
+ N_BLN<8>_XI37/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI7/MM5 N_XI37/XI7/NET34_XI37/XI7/MM5_d N_XI37/XI7/NET33_XI37/XI7/MM5_g
+ N_VDD_XI37/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI7/MM4 N_XI37/XI7/NET33_XI37/XI7/MM4_d N_XI37/XI7/NET34_XI37/XI7/MM4_g
+ N_VDD_XI37/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI7/MM10 N_XI37/XI7/NET35_XI37/XI7/MM10_d N_XI37/XI7/NET36_XI37/XI7/MM10_g
+ N_VDD_XI37/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI7/MM11 N_XI37/XI7/NET36_XI37/XI7/MM11_d N_XI37/XI7/NET35_XI37/XI7/MM11_g
+ N_VDD_XI37/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI8/MM2 N_XI37/XI8/NET34_XI37/XI8/MM2_d N_XI37/XI8/NET33_XI37/XI8/MM2_g
+ N_VSS_XI37/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM3 N_XI37/XI8/NET33_XI37/XI8/MM3_d N_WL<70>_XI37/XI8/MM3_g
+ N_BLN<7>_XI37/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM0 N_XI37/XI8/NET34_XI37/XI8/MM0_d N_WL<70>_XI37/XI8/MM0_g
+ N_BL<7>_XI37/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM1 N_XI37/XI8/NET33_XI37/XI8/MM1_d N_XI37/XI8/NET34_XI37/XI8/MM1_g
+ N_VSS_XI37/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM9 N_XI37/XI8/NET36_XI37/XI8/MM9_d N_WL<71>_XI37/XI8/MM9_g
+ N_BL<7>_XI37/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM6 N_XI37/XI8/NET35_XI37/XI8/MM6_d N_XI37/XI8/NET36_XI37/XI8/MM6_g
+ N_VSS_XI37/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM7 N_XI37/XI8/NET36_XI37/XI8/MM7_d N_XI37/XI8/NET35_XI37/XI8/MM7_g
+ N_VSS_XI37/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM8 N_XI37/XI8/NET35_XI37/XI8/MM8_d N_WL<71>_XI37/XI8/MM8_g
+ N_BLN<7>_XI37/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI8/MM5 N_XI37/XI8/NET34_XI37/XI8/MM5_d N_XI37/XI8/NET33_XI37/XI8/MM5_g
+ N_VDD_XI37/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI8/MM4 N_XI37/XI8/NET33_XI37/XI8/MM4_d N_XI37/XI8/NET34_XI37/XI8/MM4_g
+ N_VDD_XI37/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI8/MM10 N_XI37/XI8/NET35_XI37/XI8/MM10_d N_XI37/XI8/NET36_XI37/XI8/MM10_g
+ N_VDD_XI37/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI8/MM11 N_XI37/XI8/NET36_XI37/XI8/MM11_d N_XI37/XI8/NET35_XI37/XI8/MM11_g
+ N_VDD_XI37/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI9/MM2 N_XI37/XI9/NET34_XI37/XI9/MM2_d N_XI37/XI9/NET33_XI37/XI9/MM2_g
+ N_VSS_XI37/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM3 N_XI37/XI9/NET33_XI37/XI9/MM3_d N_WL<70>_XI37/XI9/MM3_g
+ N_BLN<6>_XI37/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM0 N_XI37/XI9/NET34_XI37/XI9/MM0_d N_WL<70>_XI37/XI9/MM0_g
+ N_BL<6>_XI37/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM1 N_XI37/XI9/NET33_XI37/XI9/MM1_d N_XI37/XI9/NET34_XI37/XI9/MM1_g
+ N_VSS_XI37/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM9 N_XI37/XI9/NET36_XI37/XI9/MM9_d N_WL<71>_XI37/XI9/MM9_g
+ N_BL<6>_XI37/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM6 N_XI37/XI9/NET35_XI37/XI9/MM6_d N_XI37/XI9/NET36_XI37/XI9/MM6_g
+ N_VSS_XI37/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM7 N_XI37/XI9/NET36_XI37/XI9/MM7_d N_XI37/XI9/NET35_XI37/XI9/MM7_g
+ N_VSS_XI37/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM8 N_XI37/XI9/NET35_XI37/XI9/MM8_d N_WL<71>_XI37/XI9/MM8_g
+ N_BLN<6>_XI37/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI9/MM5 N_XI37/XI9/NET34_XI37/XI9/MM5_d N_XI37/XI9/NET33_XI37/XI9/MM5_g
+ N_VDD_XI37/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI9/MM4 N_XI37/XI9/NET33_XI37/XI9/MM4_d N_XI37/XI9/NET34_XI37/XI9/MM4_g
+ N_VDD_XI37/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI9/MM10 N_XI37/XI9/NET35_XI37/XI9/MM10_d N_XI37/XI9/NET36_XI37/XI9/MM10_g
+ N_VDD_XI37/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI9/MM11 N_XI37/XI9/NET36_XI37/XI9/MM11_d N_XI37/XI9/NET35_XI37/XI9/MM11_g
+ N_VDD_XI37/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI10/MM2 N_XI37/XI10/NET34_XI37/XI10/MM2_d
+ N_XI37/XI10/NET33_XI37/XI10/MM2_g N_VSS_XI37/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI10/MM3 N_XI37/XI10/NET33_XI37/XI10/MM3_d N_WL<70>_XI37/XI10/MM3_g
+ N_BLN<5>_XI37/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI10/MM0 N_XI37/XI10/NET34_XI37/XI10/MM0_d N_WL<70>_XI37/XI10/MM0_g
+ N_BL<5>_XI37/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI10/MM1 N_XI37/XI10/NET33_XI37/XI10/MM1_d
+ N_XI37/XI10/NET34_XI37/XI10/MM1_g N_VSS_XI37/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI10/MM9 N_XI37/XI10/NET36_XI37/XI10/MM9_d N_WL<71>_XI37/XI10/MM9_g
+ N_BL<5>_XI37/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI10/MM6 N_XI37/XI10/NET35_XI37/XI10/MM6_d
+ N_XI37/XI10/NET36_XI37/XI10/MM6_g N_VSS_XI37/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI10/MM7 N_XI37/XI10/NET36_XI37/XI10/MM7_d
+ N_XI37/XI10/NET35_XI37/XI10/MM7_g N_VSS_XI37/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI10/MM8 N_XI37/XI10/NET35_XI37/XI10/MM8_d N_WL<71>_XI37/XI10/MM8_g
+ N_BLN<5>_XI37/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI10/MM5 N_XI37/XI10/NET34_XI37/XI10/MM5_d
+ N_XI37/XI10/NET33_XI37/XI10/MM5_g N_VDD_XI37/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI10/MM4 N_XI37/XI10/NET33_XI37/XI10/MM4_d
+ N_XI37/XI10/NET34_XI37/XI10/MM4_g N_VDD_XI37/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI10/MM10 N_XI37/XI10/NET35_XI37/XI10/MM10_d
+ N_XI37/XI10/NET36_XI37/XI10/MM10_g N_VDD_XI37/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI10/MM11 N_XI37/XI10/NET36_XI37/XI10/MM11_d
+ N_XI37/XI10/NET35_XI37/XI10/MM11_g N_VDD_XI37/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI11/MM2 N_XI37/XI11/NET34_XI37/XI11/MM2_d
+ N_XI37/XI11/NET33_XI37/XI11/MM2_g N_VSS_XI37/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI11/MM3 N_XI37/XI11/NET33_XI37/XI11/MM3_d N_WL<70>_XI37/XI11/MM3_g
+ N_BLN<4>_XI37/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI11/MM0 N_XI37/XI11/NET34_XI37/XI11/MM0_d N_WL<70>_XI37/XI11/MM0_g
+ N_BL<4>_XI37/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI11/MM1 N_XI37/XI11/NET33_XI37/XI11/MM1_d
+ N_XI37/XI11/NET34_XI37/XI11/MM1_g N_VSS_XI37/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI11/MM9 N_XI37/XI11/NET36_XI37/XI11/MM9_d N_WL<71>_XI37/XI11/MM9_g
+ N_BL<4>_XI37/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI11/MM6 N_XI37/XI11/NET35_XI37/XI11/MM6_d
+ N_XI37/XI11/NET36_XI37/XI11/MM6_g N_VSS_XI37/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI11/MM7 N_XI37/XI11/NET36_XI37/XI11/MM7_d
+ N_XI37/XI11/NET35_XI37/XI11/MM7_g N_VSS_XI37/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI11/MM8 N_XI37/XI11/NET35_XI37/XI11/MM8_d N_WL<71>_XI37/XI11/MM8_g
+ N_BLN<4>_XI37/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI11/MM5 N_XI37/XI11/NET34_XI37/XI11/MM5_d
+ N_XI37/XI11/NET33_XI37/XI11/MM5_g N_VDD_XI37/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI11/MM4 N_XI37/XI11/NET33_XI37/XI11/MM4_d
+ N_XI37/XI11/NET34_XI37/XI11/MM4_g N_VDD_XI37/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI11/MM10 N_XI37/XI11/NET35_XI37/XI11/MM10_d
+ N_XI37/XI11/NET36_XI37/XI11/MM10_g N_VDD_XI37/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI11/MM11 N_XI37/XI11/NET36_XI37/XI11/MM11_d
+ N_XI37/XI11/NET35_XI37/XI11/MM11_g N_VDD_XI37/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI12/MM2 N_XI37/XI12/NET34_XI37/XI12/MM2_d
+ N_XI37/XI12/NET33_XI37/XI12/MM2_g N_VSS_XI37/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI12/MM3 N_XI37/XI12/NET33_XI37/XI12/MM3_d N_WL<70>_XI37/XI12/MM3_g
+ N_BLN<3>_XI37/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI12/MM0 N_XI37/XI12/NET34_XI37/XI12/MM0_d N_WL<70>_XI37/XI12/MM0_g
+ N_BL<3>_XI37/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI12/MM1 N_XI37/XI12/NET33_XI37/XI12/MM1_d
+ N_XI37/XI12/NET34_XI37/XI12/MM1_g N_VSS_XI37/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI12/MM9 N_XI37/XI12/NET36_XI37/XI12/MM9_d N_WL<71>_XI37/XI12/MM9_g
+ N_BL<3>_XI37/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI12/MM6 N_XI37/XI12/NET35_XI37/XI12/MM6_d
+ N_XI37/XI12/NET36_XI37/XI12/MM6_g N_VSS_XI37/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI12/MM7 N_XI37/XI12/NET36_XI37/XI12/MM7_d
+ N_XI37/XI12/NET35_XI37/XI12/MM7_g N_VSS_XI37/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI12/MM8 N_XI37/XI12/NET35_XI37/XI12/MM8_d N_WL<71>_XI37/XI12/MM8_g
+ N_BLN<3>_XI37/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI12/MM5 N_XI37/XI12/NET34_XI37/XI12/MM5_d
+ N_XI37/XI12/NET33_XI37/XI12/MM5_g N_VDD_XI37/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI12/MM4 N_XI37/XI12/NET33_XI37/XI12/MM4_d
+ N_XI37/XI12/NET34_XI37/XI12/MM4_g N_VDD_XI37/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI12/MM10 N_XI37/XI12/NET35_XI37/XI12/MM10_d
+ N_XI37/XI12/NET36_XI37/XI12/MM10_g N_VDD_XI37/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI12/MM11 N_XI37/XI12/NET36_XI37/XI12/MM11_d
+ N_XI37/XI12/NET35_XI37/XI12/MM11_g N_VDD_XI37/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI13/MM2 N_XI37/XI13/NET34_XI37/XI13/MM2_d
+ N_XI37/XI13/NET33_XI37/XI13/MM2_g N_VSS_XI37/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI13/MM3 N_XI37/XI13/NET33_XI37/XI13/MM3_d N_WL<70>_XI37/XI13/MM3_g
+ N_BLN<2>_XI37/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI13/MM0 N_XI37/XI13/NET34_XI37/XI13/MM0_d N_WL<70>_XI37/XI13/MM0_g
+ N_BL<2>_XI37/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI13/MM1 N_XI37/XI13/NET33_XI37/XI13/MM1_d
+ N_XI37/XI13/NET34_XI37/XI13/MM1_g N_VSS_XI37/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI13/MM9 N_XI37/XI13/NET36_XI37/XI13/MM9_d N_WL<71>_XI37/XI13/MM9_g
+ N_BL<2>_XI37/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI13/MM6 N_XI37/XI13/NET35_XI37/XI13/MM6_d
+ N_XI37/XI13/NET36_XI37/XI13/MM6_g N_VSS_XI37/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI13/MM7 N_XI37/XI13/NET36_XI37/XI13/MM7_d
+ N_XI37/XI13/NET35_XI37/XI13/MM7_g N_VSS_XI37/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI13/MM8 N_XI37/XI13/NET35_XI37/XI13/MM8_d N_WL<71>_XI37/XI13/MM8_g
+ N_BLN<2>_XI37/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI13/MM5 N_XI37/XI13/NET34_XI37/XI13/MM5_d
+ N_XI37/XI13/NET33_XI37/XI13/MM5_g N_VDD_XI37/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI13/MM4 N_XI37/XI13/NET33_XI37/XI13/MM4_d
+ N_XI37/XI13/NET34_XI37/XI13/MM4_g N_VDD_XI37/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI13/MM10 N_XI37/XI13/NET35_XI37/XI13/MM10_d
+ N_XI37/XI13/NET36_XI37/XI13/MM10_g N_VDD_XI37/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI13/MM11 N_XI37/XI13/NET36_XI37/XI13/MM11_d
+ N_XI37/XI13/NET35_XI37/XI13/MM11_g N_VDD_XI37/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI14/MM2 N_XI37/XI14/NET34_XI37/XI14/MM2_d
+ N_XI37/XI14/NET33_XI37/XI14/MM2_g N_VSS_XI37/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI14/MM3 N_XI37/XI14/NET33_XI37/XI14/MM3_d N_WL<70>_XI37/XI14/MM3_g
+ N_BLN<1>_XI37/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI14/MM0 N_XI37/XI14/NET34_XI37/XI14/MM0_d N_WL<70>_XI37/XI14/MM0_g
+ N_BL<1>_XI37/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI14/MM1 N_XI37/XI14/NET33_XI37/XI14/MM1_d
+ N_XI37/XI14/NET34_XI37/XI14/MM1_g N_VSS_XI37/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI14/MM9 N_XI37/XI14/NET36_XI37/XI14/MM9_d N_WL<71>_XI37/XI14/MM9_g
+ N_BL<1>_XI37/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI14/MM6 N_XI37/XI14/NET35_XI37/XI14/MM6_d
+ N_XI37/XI14/NET36_XI37/XI14/MM6_g N_VSS_XI37/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI14/MM7 N_XI37/XI14/NET36_XI37/XI14/MM7_d
+ N_XI37/XI14/NET35_XI37/XI14/MM7_g N_VSS_XI37/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI14/MM8 N_XI37/XI14/NET35_XI37/XI14/MM8_d N_WL<71>_XI37/XI14/MM8_g
+ N_BLN<1>_XI37/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI14/MM5 N_XI37/XI14/NET34_XI37/XI14/MM5_d
+ N_XI37/XI14/NET33_XI37/XI14/MM5_g N_VDD_XI37/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI14/MM4 N_XI37/XI14/NET33_XI37/XI14/MM4_d
+ N_XI37/XI14/NET34_XI37/XI14/MM4_g N_VDD_XI37/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI14/MM10 N_XI37/XI14/NET35_XI37/XI14/MM10_d
+ N_XI37/XI14/NET36_XI37/XI14/MM10_g N_VDD_XI37/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI14/MM11 N_XI37/XI14/NET36_XI37/XI14/MM11_d
+ N_XI37/XI14/NET35_XI37/XI14/MM11_g N_VDD_XI37/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI15/MM2 N_XI37/XI15/NET34_XI37/XI15/MM2_d
+ N_XI37/XI15/NET33_XI37/XI15/MM2_g N_VSS_XI37/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI15/MM3 N_XI37/XI15/NET33_XI37/XI15/MM3_d N_WL<70>_XI37/XI15/MM3_g
+ N_BLN<0>_XI37/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI15/MM0 N_XI37/XI15/NET34_XI37/XI15/MM0_d N_WL<70>_XI37/XI15/MM0_g
+ N_BL<0>_XI37/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI15/MM1 N_XI37/XI15/NET33_XI37/XI15/MM1_d
+ N_XI37/XI15/NET34_XI37/XI15/MM1_g N_VSS_XI37/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI15/MM9 N_XI37/XI15/NET36_XI37/XI15/MM9_d N_WL<71>_XI37/XI15/MM9_g
+ N_BL<0>_XI37/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI15/MM6 N_XI37/XI15/NET35_XI37/XI15/MM6_d
+ N_XI37/XI15/NET36_XI37/XI15/MM6_g N_VSS_XI37/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI15/MM7 N_XI37/XI15/NET36_XI37/XI15/MM7_d
+ N_XI37/XI15/NET35_XI37/XI15/MM7_g N_VSS_XI37/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI37/XI15/MM8 N_XI37/XI15/NET35_XI37/XI15/MM8_d N_WL<71>_XI37/XI15/MM8_g
+ N_BLN<0>_XI37/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI37/XI15/MM5 N_XI37/XI15/NET34_XI37/XI15/MM5_d
+ N_XI37/XI15/NET33_XI37/XI15/MM5_g N_VDD_XI37/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI15/MM4 N_XI37/XI15/NET33_XI37/XI15/MM4_d
+ N_XI37/XI15/NET34_XI37/XI15/MM4_g N_VDD_XI37/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI15/MM10 N_XI37/XI15/NET35_XI37/XI15/MM10_d
+ N_XI37/XI15/NET36_XI37/XI15/MM10_g N_VDD_XI37/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI37/XI15/MM11 N_XI37/XI15/NET36_XI37/XI15/MM11_d
+ N_XI37/XI15/NET35_XI37/XI15/MM11_g N_VDD_XI37/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI0/MM2 N_XI38/XI0/NET34_XI38/XI0/MM2_d N_XI38/XI0/NET33_XI38/XI0/MM2_g
+ N_VSS_XI38/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI0/MM3 N_XI38/XI0/NET33_XI38/XI0/MM3_d N_WL<72>_XI38/XI0/MM3_g
+ N_BLN<15>_XI38/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI0/MM0 N_XI38/XI0/NET34_XI38/XI0/MM0_d N_WL<72>_XI38/XI0/MM0_g
+ N_BL<15>_XI38/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI0/MM1 N_XI38/XI0/NET33_XI38/XI0/MM1_d N_XI38/XI0/NET34_XI38/XI0/MM1_g
+ N_VSS_XI38/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI0/MM9 N_XI38/XI0/NET36_XI38/XI0/MM9_d N_WL<73>_XI38/XI0/MM9_g
+ N_BL<15>_XI38/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI0/MM6 N_XI38/XI0/NET35_XI38/XI0/MM6_d N_XI38/XI0/NET36_XI38/XI0/MM6_g
+ N_VSS_XI38/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI0/MM7 N_XI38/XI0/NET36_XI38/XI0/MM7_d N_XI38/XI0/NET35_XI38/XI0/MM7_g
+ N_VSS_XI38/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI0/MM8 N_XI38/XI0/NET35_XI38/XI0/MM8_d N_WL<73>_XI38/XI0/MM8_g
+ N_BLN<15>_XI38/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI0/MM5 N_XI38/XI0/NET34_XI38/XI0/MM5_d N_XI38/XI0/NET33_XI38/XI0/MM5_g
+ N_VDD_XI38/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI0/MM4 N_XI38/XI0/NET33_XI38/XI0/MM4_d N_XI38/XI0/NET34_XI38/XI0/MM4_g
+ N_VDD_XI38/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI0/MM10 N_XI38/XI0/NET35_XI38/XI0/MM10_d N_XI38/XI0/NET36_XI38/XI0/MM10_g
+ N_VDD_XI38/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI0/MM11 N_XI38/XI0/NET36_XI38/XI0/MM11_d N_XI38/XI0/NET35_XI38/XI0/MM11_g
+ N_VDD_XI38/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI1/MM2 N_XI38/XI1/NET34_XI38/XI1/MM2_d N_XI38/XI1/NET33_XI38/XI1/MM2_g
+ N_VSS_XI38/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI1/MM3 N_XI38/XI1/NET33_XI38/XI1/MM3_d N_WL<72>_XI38/XI1/MM3_g
+ N_BLN<14>_XI38/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI1/MM0 N_XI38/XI1/NET34_XI38/XI1/MM0_d N_WL<72>_XI38/XI1/MM0_g
+ N_BL<14>_XI38/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI1/MM1 N_XI38/XI1/NET33_XI38/XI1/MM1_d N_XI38/XI1/NET34_XI38/XI1/MM1_g
+ N_VSS_XI38/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI1/MM9 N_XI38/XI1/NET36_XI38/XI1/MM9_d N_WL<73>_XI38/XI1/MM9_g
+ N_BL<14>_XI38/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI1/MM6 N_XI38/XI1/NET35_XI38/XI1/MM6_d N_XI38/XI1/NET36_XI38/XI1/MM6_g
+ N_VSS_XI38/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI1/MM7 N_XI38/XI1/NET36_XI38/XI1/MM7_d N_XI38/XI1/NET35_XI38/XI1/MM7_g
+ N_VSS_XI38/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI1/MM8 N_XI38/XI1/NET35_XI38/XI1/MM8_d N_WL<73>_XI38/XI1/MM8_g
+ N_BLN<14>_XI38/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI1/MM5 N_XI38/XI1/NET34_XI38/XI1/MM5_d N_XI38/XI1/NET33_XI38/XI1/MM5_g
+ N_VDD_XI38/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI1/MM4 N_XI38/XI1/NET33_XI38/XI1/MM4_d N_XI38/XI1/NET34_XI38/XI1/MM4_g
+ N_VDD_XI38/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI1/MM10 N_XI38/XI1/NET35_XI38/XI1/MM10_d N_XI38/XI1/NET36_XI38/XI1/MM10_g
+ N_VDD_XI38/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI1/MM11 N_XI38/XI1/NET36_XI38/XI1/MM11_d N_XI38/XI1/NET35_XI38/XI1/MM11_g
+ N_VDD_XI38/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI2/MM2 N_XI38/XI2/NET34_XI38/XI2/MM2_d N_XI38/XI2/NET33_XI38/XI2/MM2_g
+ N_VSS_XI38/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI2/MM3 N_XI38/XI2/NET33_XI38/XI2/MM3_d N_WL<72>_XI38/XI2/MM3_g
+ N_BLN<13>_XI38/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI2/MM0 N_XI38/XI2/NET34_XI38/XI2/MM0_d N_WL<72>_XI38/XI2/MM0_g
+ N_BL<13>_XI38/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI2/MM1 N_XI38/XI2/NET33_XI38/XI2/MM1_d N_XI38/XI2/NET34_XI38/XI2/MM1_g
+ N_VSS_XI38/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI2/MM9 N_XI38/XI2/NET36_XI38/XI2/MM9_d N_WL<73>_XI38/XI2/MM9_g
+ N_BL<13>_XI38/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI2/MM6 N_XI38/XI2/NET35_XI38/XI2/MM6_d N_XI38/XI2/NET36_XI38/XI2/MM6_g
+ N_VSS_XI38/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI2/MM7 N_XI38/XI2/NET36_XI38/XI2/MM7_d N_XI38/XI2/NET35_XI38/XI2/MM7_g
+ N_VSS_XI38/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI2/MM8 N_XI38/XI2/NET35_XI38/XI2/MM8_d N_WL<73>_XI38/XI2/MM8_g
+ N_BLN<13>_XI38/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI2/MM5 N_XI38/XI2/NET34_XI38/XI2/MM5_d N_XI38/XI2/NET33_XI38/XI2/MM5_g
+ N_VDD_XI38/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI2/MM4 N_XI38/XI2/NET33_XI38/XI2/MM4_d N_XI38/XI2/NET34_XI38/XI2/MM4_g
+ N_VDD_XI38/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI2/MM10 N_XI38/XI2/NET35_XI38/XI2/MM10_d N_XI38/XI2/NET36_XI38/XI2/MM10_g
+ N_VDD_XI38/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI2/MM11 N_XI38/XI2/NET36_XI38/XI2/MM11_d N_XI38/XI2/NET35_XI38/XI2/MM11_g
+ N_VDD_XI38/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI3/MM2 N_XI38/XI3/NET34_XI38/XI3/MM2_d N_XI38/XI3/NET33_XI38/XI3/MM2_g
+ N_VSS_XI38/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI3/MM3 N_XI38/XI3/NET33_XI38/XI3/MM3_d N_WL<72>_XI38/XI3/MM3_g
+ N_BLN<12>_XI38/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI3/MM0 N_XI38/XI3/NET34_XI38/XI3/MM0_d N_WL<72>_XI38/XI3/MM0_g
+ N_BL<12>_XI38/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI3/MM1 N_XI38/XI3/NET33_XI38/XI3/MM1_d N_XI38/XI3/NET34_XI38/XI3/MM1_g
+ N_VSS_XI38/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI3/MM9 N_XI38/XI3/NET36_XI38/XI3/MM9_d N_WL<73>_XI38/XI3/MM9_g
+ N_BL<12>_XI38/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI3/MM6 N_XI38/XI3/NET35_XI38/XI3/MM6_d N_XI38/XI3/NET36_XI38/XI3/MM6_g
+ N_VSS_XI38/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI3/MM7 N_XI38/XI3/NET36_XI38/XI3/MM7_d N_XI38/XI3/NET35_XI38/XI3/MM7_g
+ N_VSS_XI38/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI3/MM8 N_XI38/XI3/NET35_XI38/XI3/MM8_d N_WL<73>_XI38/XI3/MM8_g
+ N_BLN<12>_XI38/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI3/MM5 N_XI38/XI3/NET34_XI38/XI3/MM5_d N_XI38/XI3/NET33_XI38/XI3/MM5_g
+ N_VDD_XI38/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI3/MM4 N_XI38/XI3/NET33_XI38/XI3/MM4_d N_XI38/XI3/NET34_XI38/XI3/MM4_g
+ N_VDD_XI38/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI3/MM10 N_XI38/XI3/NET35_XI38/XI3/MM10_d N_XI38/XI3/NET36_XI38/XI3/MM10_g
+ N_VDD_XI38/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI3/MM11 N_XI38/XI3/NET36_XI38/XI3/MM11_d N_XI38/XI3/NET35_XI38/XI3/MM11_g
+ N_VDD_XI38/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI4/MM2 N_XI38/XI4/NET34_XI38/XI4/MM2_d N_XI38/XI4/NET33_XI38/XI4/MM2_g
+ N_VSS_XI38/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI4/MM3 N_XI38/XI4/NET33_XI38/XI4/MM3_d N_WL<72>_XI38/XI4/MM3_g
+ N_BLN<11>_XI38/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI4/MM0 N_XI38/XI4/NET34_XI38/XI4/MM0_d N_WL<72>_XI38/XI4/MM0_g
+ N_BL<11>_XI38/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI4/MM1 N_XI38/XI4/NET33_XI38/XI4/MM1_d N_XI38/XI4/NET34_XI38/XI4/MM1_g
+ N_VSS_XI38/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI4/MM9 N_XI38/XI4/NET36_XI38/XI4/MM9_d N_WL<73>_XI38/XI4/MM9_g
+ N_BL<11>_XI38/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI4/MM6 N_XI38/XI4/NET35_XI38/XI4/MM6_d N_XI38/XI4/NET36_XI38/XI4/MM6_g
+ N_VSS_XI38/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI4/MM7 N_XI38/XI4/NET36_XI38/XI4/MM7_d N_XI38/XI4/NET35_XI38/XI4/MM7_g
+ N_VSS_XI38/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI4/MM8 N_XI38/XI4/NET35_XI38/XI4/MM8_d N_WL<73>_XI38/XI4/MM8_g
+ N_BLN<11>_XI38/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI4/MM5 N_XI38/XI4/NET34_XI38/XI4/MM5_d N_XI38/XI4/NET33_XI38/XI4/MM5_g
+ N_VDD_XI38/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI4/MM4 N_XI38/XI4/NET33_XI38/XI4/MM4_d N_XI38/XI4/NET34_XI38/XI4/MM4_g
+ N_VDD_XI38/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI4/MM10 N_XI38/XI4/NET35_XI38/XI4/MM10_d N_XI38/XI4/NET36_XI38/XI4/MM10_g
+ N_VDD_XI38/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI4/MM11 N_XI38/XI4/NET36_XI38/XI4/MM11_d N_XI38/XI4/NET35_XI38/XI4/MM11_g
+ N_VDD_XI38/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI5/MM2 N_XI38/XI5/NET34_XI38/XI5/MM2_d N_XI38/XI5/NET33_XI38/XI5/MM2_g
+ N_VSS_XI38/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI5/MM3 N_XI38/XI5/NET33_XI38/XI5/MM3_d N_WL<72>_XI38/XI5/MM3_g
+ N_BLN<10>_XI38/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI5/MM0 N_XI38/XI5/NET34_XI38/XI5/MM0_d N_WL<72>_XI38/XI5/MM0_g
+ N_BL<10>_XI38/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI5/MM1 N_XI38/XI5/NET33_XI38/XI5/MM1_d N_XI38/XI5/NET34_XI38/XI5/MM1_g
+ N_VSS_XI38/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI5/MM9 N_XI38/XI5/NET36_XI38/XI5/MM9_d N_WL<73>_XI38/XI5/MM9_g
+ N_BL<10>_XI38/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI5/MM6 N_XI38/XI5/NET35_XI38/XI5/MM6_d N_XI38/XI5/NET36_XI38/XI5/MM6_g
+ N_VSS_XI38/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI5/MM7 N_XI38/XI5/NET36_XI38/XI5/MM7_d N_XI38/XI5/NET35_XI38/XI5/MM7_g
+ N_VSS_XI38/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI5/MM8 N_XI38/XI5/NET35_XI38/XI5/MM8_d N_WL<73>_XI38/XI5/MM8_g
+ N_BLN<10>_XI38/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI5/MM5 N_XI38/XI5/NET34_XI38/XI5/MM5_d N_XI38/XI5/NET33_XI38/XI5/MM5_g
+ N_VDD_XI38/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI5/MM4 N_XI38/XI5/NET33_XI38/XI5/MM4_d N_XI38/XI5/NET34_XI38/XI5/MM4_g
+ N_VDD_XI38/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI5/MM10 N_XI38/XI5/NET35_XI38/XI5/MM10_d N_XI38/XI5/NET36_XI38/XI5/MM10_g
+ N_VDD_XI38/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI5/MM11 N_XI38/XI5/NET36_XI38/XI5/MM11_d N_XI38/XI5/NET35_XI38/XI5/MM11_g
+ N_VDD_XI38/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI6/MM2 N_XI38/XI6/NET34_XI38/XI6/MM2_d N_XI38/XI6/NET33_XI38/XI6/MM2_g
+ N_VSS_XI38/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM3 N_XI38/XI6/NET33_XI38/XI6/MM3_d N_WL<72>_XI38/XI6/MM3_g
+ N_BLN<9>_XI38/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM0 N_XI38/XI6/NET34_XI38/XI6/MM0_d N_WL<72>_XI38/XI6/MM0_g
+ N_BL<9>_XI38/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM1 N_XI38/XI6/NET33_XI38/XI6/MM1_d N_XI38/XI6/NET34_XI38/XI6/MM1_g
+ N_VSS_XI38/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM9 N_XI38/XI6/NET36_XI38/XI6/MM9_d N_WL<73>_XI38/XI6/MM9_g
+ N_BL<9>_XI38/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM6 N_XI38/XI6/NET35_XI38/XI6/MM6_d N_XI38/XI6/NET36_XI38/XI6/MM6_g
+ N_VSS_XI38/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM7 N_XI38/XI6/NET36_XI38/XI6/MM7_d N_XI38/XI6/NET35_XI38/XI6/MM7_g
+ N_VSS_XI38/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM8 N_XI38/XI6/NET35_XI38/XI6/MM8_d N_WL<73>_XI38/XI6/MM8_g
+ N_BLN<9>_XI38/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI6/MM5 N_XI38/XI6/NET34_XI38/XI6/MM5_d N_XI38/XI6/NET33_XI38/XI6/MM5_g
+ N_VDD_XI38/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI6/MM4 N_XI38/XI6/NET33_XI38/XI6/MM4_d N_XI38/XI6/NET34_XI38/XI6/MM4_g
+ N_VDD_XI38/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI6/MM10 N_XI38/XI6/NET35_XI38/XI6/MM10_d N_XI38/XI6/NET36_XI38/XI6/MM10_g
+ N_VDD_XI38/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI6/MM11 N_XI38/XI6/NET36_XI38/XI6/MM11_d N_XI38/XI6/NET35_XI38/XI6/MM11_g
+ N_VDD_XI38/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI7/MM2 N_XI38/XI7/NET34_XI38/XI7/MM2_d N_XI38/XI7/NET33_XI38/XI7/MM2_g
+ N_VSS_XI38/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM3 N_XI38/XI7/NET33_XI38/XI7/MM3_d N_WL<72>_XI38/XI7/MM3_g
+ N_BLN<8>_XI38/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM0 N_XI38/XI7/NET34_XI38/XI7/MM0_d N_WL<72>_XI38/XI7/MM0_g
+ N_BL<8>_XI38/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM1 N_XI38/XI7/NET33_XI38/XI7/MM1_d N_XI38/XI7/NET34_XI38/XI7/MM1_g
+ N_VSS_XI38/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM9 N_XI38/XI7/NET36_XI38/XI7/MM9_d N_WL<73>_XI38/XI7/MM9_g
+ N_BL<8>_XI38/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM6 N_XI38/XI7/NET35_XI38/XI7/MM6_d N_XI38/XI7/NET36_XI38/XI7/MM6_g
+ N_VSS_XI38/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM7 N_XI38/XI7/NET36_XI38/XI7/MM7_d N_XI38/XI7/NET35_XI38/XI7/MM7_g
+ N_VSS_XI38/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM8 N_XI38/XI7/NET35_XI38/XI7/MM8_d N_WL<73>_XI38/XI7/MM8_g
+ N_BLN<8>_XI38/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI7/MM5 N_XI38/XI7/NET34_XI38/XI7/MM5_d N_XI38/XI7/NET33_XI38/XI7/MM5_g
+ N_VDD_XI38/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI7/MM4 N_XI38/XI7/NET33_XI38/XI7/MM4_d N_XI38/XI7/NET34_XI38/XI7/MM4_g
+ N_VDD_XI38/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI7/MM10 N_XI38/XI7/NET35_XI38/XI7/MM10_d N_XI38/XI7/NET36_XI38/XI7/MM10_g
+ N_VDD_XI38/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI7/MM11 N_XI38/XI7/NET36_XI38/XI7/MM11_d N_XI38/XI7/NET35_XI38/XI7/MM11_g
+ N_VDD_XI38/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI8/MM2 N_XI38/XI8/NET34_XI38/XI8/MM2_d N_XI38/XI8/NET33_XI38/XI8/MM2_g
+ N_VSS_XI38/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM3 N_XI38/XI8/NET33_XI38/XI8/MM3_d N_WL<72>_XI38/XI8/MM3_g
+ N_BLN<7>_XI38/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM0 N_XI38/XI8/NET34_XI38/XI8/MM0_d N_WL<72>_XI38/XI8/MM0_g
+ N_BL<7>_XI38/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM1 N_XI38/XI8/NET33_XI38/XI8/MM1_d N_XI38/XI8/NET34_XI38/XI8/MM1_g
+ N_VSS_XI38/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM9 N_XI38/XI8/NET36_XI38/XI8/MM9_d N_WL<73>_XI38/XI8/MM9_g
+ N_BL<7>_XI38/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM6 N_XI38/XI8/NET35_XI38/XI8/MM6_d N_XI38/XI8/NET36_XI38/XI8/MM6_g
+ N_VSS_XI38/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM7 N_XI38/XI8/NET36_XI38/XI8/MM7_d N_XI38/XI8/NET35_XI38/XI8/MM7_g
+ N_VSS_XI38/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM8 N_XI38/XI8/NET35_XI38/XI8/MM8_d N_WL<73>_XI38/XI8/MM8_g
+ N_BLN<7>_XI38/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI8/MM5 N_XI38/XI8/NET34_XI38/XI8/MM5_d N_XI38/XI8/NET33_XI38/XI8/MM5_g
+ N_VDD_XI38/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI8/MM4 N_XI38/XI8/NET33_XI38/XI8/MM4_d N_XI38/XI8/NET34_XI38/XI8/MM4_g
+ N_VDD_XI38/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI8/MM10 N_XI38/XI8/NET35_XI38/XI8/MM10_d N_XI38/XI8/NET36_XI38/XI8/MM10_g
+ N_VDD_XI38/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI8/MM11 N_XI38/XI8/NET36_XI38/XI8/MM11_d N_XI38/XI8/NET35_XI38/XI8/MM11_g
+ N_VDD_XI38/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI9/MM2 N_XI38/XI9/NET34_XI38/XI9/MM2_d N_XI38/XI9/NET33_XI38/XI9/MM2_g
+ N_VSS_XI38/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM3 N_XI38/XI9/NET33_XI38/XI9/MM3_d N_WL<72>_XI38/XI9/MM3_g
+ N_BLN<6>_XI38/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM0 N_XI38/XI9/NET34_XI38/XI9/MM0_d N_WL<72>_XI38/XI9/MM0_g
+ N_BL<6>_XI38/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM1 N_XI38/XI9/NET33_XI38/XI9/MM1_d N_XI38/XI9/NET34_XI38/XI9/MM1_g
+ N_VSS_XI38/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM9 N_XI38/XI9/NET36_XI38/XI9/MM9_d N_WL<73>_XI38/XI9/MM9_g
+ N_BL<6>_XI38/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM6 N_XI38/XI9/NET35_XI38/XI9/MM6_d N_XI38/XI9/NET36_XI38/XI9/MM6_g
+ N_VSS_XI38/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM7 N_XI38/XI9/NET36_XI38/XI9/MM7_d N_XI38/XI9/NET35_XI38/XI9/MM7_g
+ N_VSS_XI38/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM8 N_XI38/XI9/NET35_XI38/XI9/MM8_d N_WL<73>_XI38/XI9/MM8_g
+ N_BLN<6>_XI38/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI9/MM5 N_XI38/XI9/NET34_XI38/XI9/MM5_d N_XI38/XI9/NET33_XI38/XI9/MM5_g
+ N_VDD_XI38/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI9/MM4 N_XI38/XI9/NET33_XI38/XI9/MM4_d N_XI38/XI9/NET34_XI38/XI9/MM4_g
+ N_VDD_XI38/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI9/MM10 N_XI38/XI9/NET35_XI38/XI9/MM10_d N_XI38/XI9/NET36_XI38/XI9/MM10_g
+ N_VDD_XI38/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI9/MM11 N_XI38/XI9/NET36_XI38/XI9/MM11_d N_XI38/XI9/NET35_XI38/XI9/MM11_g
+ N_VDD_XI38/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI10/MM2 N_XI38/XI10/NET34_XI38/XI10/MM2_d
+ N_XI38/XI10/NET33_XI38/XI10/MM2_g N_VSS_XI38/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI10/MM3 N_XI38/XI10/NET33_XI38/XI10/MM3_d N_WL<72>_XI38/XI10/MM3_g
+ N_BLN<5>_XI38/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI10/MM0 N_XI38/XI10/NET34_XI38/XI10/MM0_d N_WL<72>_XI38/XI10/MM0_g
+ N_BL<5>_XI38/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI10/MM1 N_XI38/XI10/NET33_XI38/XI10/MM1_d
+ N_XI38/XI10/NET34_XI38/XI10/MM1_g N_VSS_XI38/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI10/MM9 N_XI38/XI10/NET36_XI38/XI10/MM9_d N_WL<73>_XI38/XI10/MM9_g
+ N_BL<5>_XI38/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI10/MM6 N_XI38/XI10/NET35_XI38/XI10/MM6_d
+ N_XI38/XI10/NET36_XI38/XI10/MM6_g N_VSS_XI38/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI10/MM7 N_XI38/XI10/NET36_XI38/XI10/MM7_d
+ N_XI38/XI10/NET35_XI38/XI10/MM7_g N_VSS_XI38/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI10/MM8 N_XI38/XI10/NET35_XI38/XI10/MM8_d N_WL<73>_XI38/XI10/MM8_g
+ N_BLN<5>_XI38/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI10/MM5 N_XI38/XI10/NET34_XI38/XI10/MM5_d
+ N_XI38/XI10/NET33_XI38/XI10/MM5_g N_VDD_XI38/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI10/MM4 N_XI38/XI10/NET33_XI38/XI10/MM4_d
+ N_XI38/XI10/NET34_XI38/XI10/MM4_g N_VDD_XI38/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI10/MM10 N_XI38/XI10/NET35_XI38/XI10/MM10_d
+ N_XI38/XI10/NET36_XI38/XI10/MM10_g N_VDD_XI38/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI10/MM11 N_XI38/XI10/NET36_XI38/XI10/MM11_d
+ N_XI38/XI10/NET35_XI38/XI10/MM11_g N_VDD_XI38/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI11/MM2 N_XI38/XI11/NET34_XI38/XI11/MM2_d
+ N_XI38/XI11/NET33_XI38/XI11/MM2_g N_VSS_XI38/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI11/MM3 N_XI38/XI11/NET33_XI38/XI11/MM3_d N_WL<72>_XI38/XI11/MM3_g
+ N_BLN<4>_XI38/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI11/MM0 N_XI38/XI11/NET34_XI38/XI11/MM0_d N_WL<72>_XI38/XI11/MM0_g
+ N_BL<4>_XI38/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI11/MM1 N_XI38/XI11/NET33_XI38/XI11/MM1_d
+ N_XI38/XI11/NET34_XI38/XI11/MM1_g N_VSS_XI38/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI11/MM9 N_XI38/XI11/NET36_XI38/XI11/MM9_d N_WL<73>_XI38/XI11/MM9_g
+ N_BL<4>_XI38/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI11/MM6 N_XI38/XI11/NET35_XI38/XI11/MM6_d
+ N_XI38/XI11/NET36_XI38/XI11/MM6_g N_VSS_XI38/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI11/MM7 N_XI38/XI11/NET36_XI38/XI11/MM7_d
+ N_XI38/XI11/NET35_XI38/XI11/MM7_g N_VSS_XI38/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI11/MM8 N_XI38/XI11/NET35_XI38/XI11/MM8_d N_WL<73>_XI38/XI11/MM8_g
+ N_BLN<4>_XI38/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI11/MM5 N_XI38/XI11/NET34_XI38/XI11/MM5_d
+ N_XI38/XI11/NET33_XI38/XI11/MM5_g N_VDD_XI38/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI11/MM4 N_XI38/XI11/NET33_XI38/XI11/MM4_d
+ N_XI38/XI11/NET34_XI38/XI11/MM4_g N_VDD_XI38/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI11/MM10 N_XI38/XI11/NET35_XI38/XI11/MM10_d
+ N_XI38/XI11/NET36_XI38/XI11/MM10_g N_VDD_XI38/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI11/MM11 N_XI38/XI11/NET36_XI38/XI11/MM11_d
+ N_XI38/XI11/NET35_XI38/XI11/MM11_g N_VDD_XI38/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI12/MM2 N_XI38/XI12/NET34_XI38/XI12/MM2_d
+ N_XI38/XI12/NET33_XI38/XI12/MM2_g N_VSS_XI38/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI12/MM3 N_XI38/XI12/NET33_XI38/XI12/MM3_d N_WL<72>_XI38/XI12/MM3_g
+ N_BLN<3>_XI38/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI12/MM0 N_XI38/XI12/NET34_XI38/XI12/MM0_d N_WL<72>_XI38/XI12/MM0_g
+ N_BL<3>_XI38/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI12/MM1 N_XI38/XI12/NET33_XI38/XI12/MM1_d
+ N_XI38/XI12/NET34_XI38/XI12/MM1_g N_VSS_XI38/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI12/MM9 N_XI38/XI12/NET36_XI38/XI12/MM9_d N_WL<73>_XI38/XI12/MM9_g
+ N_BL<3>_XI38/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI12/MM6 N_XI38/XI12/NET35_XI38/XI12/MM6_d
+ N_XI38/XI12/NET36_XI38/XI12/MM6_g N_VSS_XI38/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI12/MM7 N_XI38/XI12/NET36_XI38/XI12/MM7_d
+ N_XI38/XI12/NET35_XI38/XI12/MM7_g N_VSS_XI38/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI12/MM8 N_XI38/XI12/NET35_XI38/XI12/MM8_d N_WL<73>_XI38/XI12/MM8_g
+ N_BLN<3>_XI38/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI12/MM5 N_XI38/XI12/NET34_XI38/XI12/MM5_d
+ N_XI38/XI12/NET33_XI38/XI12/MM5_g N_VDD_XI38/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI12/MM4 N_XI38/XI12/NET33_XI38/XI12/MM4_d
+ N_XI38/XI12/NET34_XI38/XI12/MM4_g N_VDD_XI38/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI12/MM10 N_XI38/XI12/NET35_XI38/XI12/MM10_d
+ N_XI38/XI12/NET36_XI38/XI12/MM10_g N_VDD_XI38/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI12/MM11 N_XI38/XI12/NET36_XI38/XI12/MM11_d
+ N_XI38/XI12/NET35_XI38/XI12/MM11_g N_VDD_XI38/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI13/MM2 N_XI38/XI13/NET34_XI38/XI13/MM2_d
+ N_XI38/XI13/NET33_XI38/XI13/MM2_g N_VSS_XI38/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI13/MM3 N_XI38/XI13/NET33_XI38/XI13/MM3_d N_WL<72>_XI38/XI13/MM3_g
+ N_BLN<2>_XI38/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI13/MM0 N_XI38/XI13/NET34_XI38/XI13/MM0_d N_WL<72>_XI38/XI13/MM0_g
+ N_BL<2>_XI38/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI13/MM1 N_XI38/XI13/NET33_XI38/XI13/MM1_d
+ N_XI38/XI13/NET34_XI38/XI13/MM1_g N_VSS_XI38/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI13/MM9 N_XI38/XI13/NET36_XI38/XI13/MM9_d N_WL<73>_XI38/XI13/MM9_g
+ N_BL<2>_XI38/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI13/MM6 N_XI38/XI13/NET35_XI38/XI13/MM6_d
+ N_XI38/XI13/NET36_XI38/XI13/MM6_g N_VSS_XI38/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI13/MM7 N_XI38/XI13/NET36_XI38/XI13/MM7_d
+ N_XI38/XI13/NET35_XI38/XI13/MM7_g N_VSS_XI38/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI13/MM8 N_XI38/XI13/NET35_XI38/XI13/MM8_d N_WL<73>_XI38/XI13/MM8_g
+ N_BLN<2>_XI38/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI13/MM5 N_XI38/XI13/NET34_XI38/XI13/MM5_d
+ N_XI38/XI13/NET33_XI38/XI13/MM5_g N_VDD_XI38/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI13/MM4 N_XI38/XI13/NET33_XI38/XI13/MM4_d
+ N_XI38/XI13/NET34_XI38/XI13/MM4_g N_VDD_XI38/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI13/MM10 N_XI38/XI13/NET35_XI38/XI13/MM10_d
+ N_XI38/XI13/NET36_XI38/XI13/MM10_g N_VDD_XI38/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI13/MM11 N_XI38/XI13/NET36_XI38/XI13/MM11_d
+ N_XI38/XI13/NET35_XI38/XI13/MM11_g N_VDD_XI38/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI14/MM2 N_XI38/XI14/NET34_XI38/XI14/MM2_d
+ N_XI38/XI14/NET33_XI38/XI14/MM2_g N_VSS_XI38/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI14/MM3 N_XI38/XI14/NET33_XI38/XI14/MM3_d N_WL<72>_XI38/XI14/MM3_g
+ N_BLN<1>_XI38/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI14/MM0 N_XI38/XI14/NET34_XI38/XI14/MM0_d N_WL<72>_XI38/XI14/MM0_g
+ N_BL<1>_XI38/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI14/MM1 N_XI38/XI14/NET33_XI38/XI14/MM1_d
+ N_XI38/XI14/NET34_XI38/XI14/MM1_g N_VSS_XI38/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI14/MM9 N_XI38/XI14/NET36_XI38/XI14/MM9_d N_WL<73>_XI38/XI14/MM9_g
+ N_BL<1>_XI38/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI14/MM6 N_XI38/XI14/NET35_XI38/XI14/MM6_d
+ N_XI38/XI14/NET36_XI38/XI14/MM6_g N_VSS_XI38/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI14/MM7 N_XI38/XI14/NET36_XI38/XI14/MM7_d
+ N_XI38/XI14/NET35_XI38/XI14/MM7_g N_VSS_XI38/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI14/MM8 N_XI38/XI14/NET35_XI38/XI14/MM8_d N_WL<73>_XI38/XI14/MM8_g
+ N_BLN<1>_XI38/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI14/MM5 N_XI38/XI14/NET34_XI38/XI14/MM5_d
+ N_XI38/XI14/NET33_XI38/XI14/MM5_g N_VDD_XI38/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI14/MM4 N_XI38/XI14/NET33_XI38/XI14/MM4_d
+ N_XI38/XI14/NET34_XI38/XI14/MM4_g N_VDD_XI38/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI14/MM10 N_XI38/XI14/NET35_XI38/XI14/MM10_d
+ N_XI38/XI14/NET36_XI38/XI14/MM10_g N_VDD_XI38/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI14/MM11 N_XI38/XI14/NET36_XI38/XI14/MM11_d
+ N_XI38/XI14/NET35_XI38/XI14/MM11_g N_VDD_XI38/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI15/MM2 N_XI38/XI15/NET34_XI38/XI15/MM2_d
+ N_XI38/XI15/NET33_XI38/XI15/MM2_g N_VSS_XI38/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI15/MM3 N_XI38/XI15/NET33_XI38/XI15/MM3_d N_WL<72>_XI38/XI15/MM3_g
+ N_BLN<0>_XI38/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI15/MM0 N_XI38/XI15/NET34_XI38/XI15/MM0_d N_WL<72>_XI38/XI15/MM0_g
+ N_BL<0>_XI38/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI15/MM1 N_XI38/XI15/NET33_XI38/XI15/MM1_d
+ N_XI38/XI15/NET34_XI38/XI15/MM1_g N_VSS_XI38/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI15/MM9 N_XI38/XI15/NET36_XI38/XI15/MM9_d N_WL<73>_XI38/XI15/MM9_g
+ N_BL<0>_XI38/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI15/MM6 N_XI38/XI15/NET35_XI38/XI15/MM6_d
+ N_XI38/XI15/NET36_XI38/XI15/MM6_g N_VSS_XI38/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI15/MM7 N_XI38/XI15/NET36_XI38/XI15/MM7_d
+ N_XI38/XI15/NET35_XI38/XI15/MM7_g N_VSS_XI38/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI38/XI15/MM8 N_XI38/XI15/NET35_XI38/XI15/MM8_d N_WL<73>_XI38/XI15/MM8_g
+ N_BLN<0>_XI38/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI38/XI15/MM5 N_XI38/XI15/NET34_XI38/XI15/MM5_d
+ N_XI38/XI15/NET33_XI38/XI15/MM5_g N_VDD_XI38/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI15/MM4 N_XI38/XI15/NET33_XI38/XI15/MM4_d
+ N_XI38/XI15/NET34_XI38/XI15/MM4_g N_VDD_XI38/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI15/MM10 N_XI38/XI15/NET35_XI38/XI15/MM10_d
+ N_XI38/XI15/NET36_XI38/XI15/MM10_g N_VDD_XI38/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI38/XI15/MM11 N_XI38/XI15/NET36_XI38/XI15/MM11_d
+ N_XI38/XI15/NET35_XI38/XI15/MM11_g N_VDD_XI38/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI0/MM2 N_XI39/XI0/NET34_XI39/XI0/MM2_d N_XI39/XI0/NET33_XI39/XI0/MM2_g
+ N_VSS_XI39/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI0/MM3 N_XI39/XI0/NET33_XI39/XI0/MM3_d N_WL<74>_XI39/XI0/MM3_g
+ N_BLN<15>_XI39/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI0/MM0 N_XI39/XI0/NET34_XI39/XI0/MM0_d N_WL<74>_XI39/XI0/MM0_g
+ N_BL<15>_XI39/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI0/MM1 N_XI39/XI0/NET33_XI39/XI0/MM1_d N_XI39/XI0/NET34_XI39/XI0/MM1_g
+ N_VSS_XI39/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI0/MM9 N_XI39/XI0/NET36_XI39/XI0/MM9_d N_WL<75>_XI39/XI0/MM9_g
+ N_BL<15>_XI39/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI0/MM6 N_XI39/XI0/NET35_XI39/XI0/MM6_d N_XI39/XI0/NET36_XI39/XI0/MM6_g
+ N_VSS_XI39/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI0/MM7 N_XI39/XI0/NET36_XI39/XI0/MM7_d N_XI39/XI0/NET35_XI39/XI0/MM7_g
+ N_VSS_XI39/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI0/MM8 N_XI39/XI0/NET35_XI39/XI0/MM8_d N_WL<75>_XI39/XI0/MM8_g
+ N_BLN<15>_XI39/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI0/MM5 N_XI39/XI0/NET34_XI39/XI0/MM5_d N_XI39/XI0/NET33_XI39/XI0/MM5_g
+ N_VDD_XI39/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI0/MM4 N_XI39/XI0/NET33_XI39/XI0/MM4_d N_XI39/XI0/NET34_XI39/XI0/MM4_g
+ N_VDD_XI39/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI0/MM10 N_XI39/XI0/NET35_XI39/XI0/MM10_d N_XI39/XI0/NET36_XI39/XI0/MM10_g
+ N_VDD_XI39/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI0/MM11 N_XI39/XI0/NET36_XI39/XI0/MM11_d N_XI39/XI0/NET35_XI39/XI0/MM11_g
+ N_VDD_XI39/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI1/MM2 N_XI39/XI1/NET34_XI39/XI1/MM2_d N_XI39/XI1/NET33_XI39/XI1/MM2_g
+ N_VSS_XI39/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI1/MM3 N_XI39/XI1/NET33_XI39/XI1/MM3_d N_WL<74>_XI39/XI1/MM3_g
+ N_BLN<14>_XI39/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI1/MM0 N_XI39/XI1/NET34_XI39/XI1/MM0_d N_WL<74>_XI39/XI1/MM0_g
+ N_BL<14>_XI39/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI1/MM1 N_XI39/XI1/NET33_XI39/XI1/MM1_d N_XI39/XI1/NET34_XI39/XI1/MM1_g
+ N_VSS_XI39/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI1/MM9 N_XI39/XI1/NET36_XI39/XI1/MM9_d N_WL<75>_XI39/XI1/MM9_g
+ N_BL<14>_XI39/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI1/MM6 N_XI39/XI1/NET35_XI39/XI1/MM6_d N_XI39/XI1/NET36_XI39/XI1/MM6_g
+ N_VSS_XI39/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI1/MM7 N_XI39/XI1/NET36_XI39/XI1/MM7_d N_XI39/XI1/NET35_XI39/XI1/MM7_g
+ N_VSS_XI39/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI1/MM8 N_XI39/XI1/NET35_XI39/XI1/MM8_d N_WL<75>_XI39/XI1/MM8_g
+ N_BLN<14>_XI39/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI1/MM5 N_XI39/XI1/NET34_XI39/XI1/MM5_d N_XI39/XI1/NET33_XI39/XI1/MM5_g
+ N_VDD_XI39/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI1/MM4 N_XI39/XI1/NET33_XI39/XI1/MM4_d N_XI39/XI1/NET34_XI39/XI1/MM4_g
+ N_VDD_XI39/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI1/MM10 N_XI39/XI1/NET35_XI39/XI1/MM10_d N_XI39/XI1/NET36_XI39/XI1/MM10_g
+ N_VDD_XI39/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI1/MM11 N_XI39/XI1/NET36_XI39/XI1/MM11_d N_XI39/XI1/NET35_XI39/XI1/MM11_g
+ N_VDD_XI39/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI2/MM2 N_XI39/XI2/NET34_XI39/XI2/MM2_d N_XI39/XI2/NET33_XI39/XI2/MM2_g
+ N_VSS_XI39/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI2/MM3 N_XI39/XI2/NET33_XI39/XI2/MM3_d N_WL<74>_XI39/XI2/MM3_g
+ N_BLN<13>_XI39/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI2/MM0 N_XI39/XI2/NET34_XI39/XI2/MM0_d N_WL<74>_XI39/XI2/MM0_g
+ N_BL<13>_XI39/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI2/MM1 N_XI39/XI2/NET33_XI39/XI2/MM1_d N_XI39/XI2/NET34_XI39/XI2/MM1_g
+ N_VSS_XI39/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI2/MM9 N_XI39/XI2/NET36_XI39/XI2/MM9_d N_WL<75>_XI39/XI2/MM9_g
+ N_BL<13>_XI39/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI2/MM6 N_XI39/XI2/NET35_XI39/XI2/MM6_d N_XI39/XI2/NET36_XI39/XI2/MM6_g
+ N_VSS_XI39/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI2/MM7 N_XI39/XI2/NET36_XI39/XI2/MM7_d N_XI39/XI2/NET35_XI39/XI2/MM7_g
+ N_VSS_XI39/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI2/MM8 N_XI39/XI2/NET35_XI39/XI2/MM8_d N_WL<75>_XI39/XI2/MM8_g
+ N_BLN<13>_XI39/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI2/MM5 N_XI39/XI2/NET34_XI39/XI2/MM5_d N_XI39/XI2/NET33_XI39/XI2/MM5_g
+ N_VDD_XI39/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI2/MM4 N_XI39/XI2/NET33_XI39/XI2/MM4_d N_XI39/XI2/NET34_XI39/XI2/MM4_g
+ N_VDD_XI39/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI2/MM10 N_XI39/XI2/NET35_XI39/XI2/MM10_d N_XI39/XI2/NET36_XI39/XI2/MM10_g
+ N_VDD_XI39/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI2/MM11 N_XI39/XI2/NET36_XI39/XI2/MM11_d N_XI39/XI2/NET35_XI39/XI2/MM11_g
+ N_VDD_XI39/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI3/MM2 N_XI39/XI3/NET34_XI39/XI3/MM2_d N_XI39/XI3/NET33_XI39/XI3/MM2_g
+ N_VSS_XI39/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI3/MM3 N_XI39/XI3/NET33_XI39/XI3/MM3_d N_WL<74>_XI39/XI3/MM3_g
+ N_BLN<12>_XI39/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI3/MM0 N_XI39/XI3/NET34_XI39/XI3/MM0_d N_WL<74>_XI39/XI3/MM0_g
+ N_BL<12>_XI39/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI3/MM1 N_XI39/XI3/NET33_XI39/XI3/MM1_d N_XI39/XI3/NET34_XI39/XI3/MM1_g
+ N_VSS_XI39/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI3/MM9 N_XI39/XI3/NET36_XI39/XI3/MM9_d N_WL<75>_XI39/XI3/MM9_g
+ N_BL<12>_XI39/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI3/MM6 N_XI39/XI3/NET35_XI39/XI3/MM6_d N_XI39/XI3/NET36_XI39/XI3/MM6_g
+ N_VSS_XI39/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI3/MM7 N_XI39/XI3/NET36_XI39/XI3/MM7_d N_XI39/XI3/NET35_XI39/XI3/MM7_g
+ N_VSS_XI39/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI3/MM8 N_XI39/XI3/NET35_XI39/XI3/MM8_d N_WL<75>_XI39/XI3/MM8_g
+ N_BLN<12>_XI39/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI3/MM5 N_XI39/XI3/NET34_XI39/XI3/MM5_d N_XI39/XI3/NET33_XI39/XI3/MM5_g
+ N_VDD_XI39/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI3/MM4 N_XI39/XI3/NET33_XI39/XI3/MM4_d N_XI39/XI3/NET34_XI39/XI3/MM4_g
+ N_VDD_XI39/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI3/MM10 N_XI39/XI3/NET35_XI39/XI3/MM10_d N_XI39/XI3/NET36_XI39/XI3/MM10_g
+ N_VDD_XI39/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI3/MM11 N_XI39/XI3/NET36_XI39/XI3/MM11_d N_XI39/XI3/NET35_XI39/XI3/MM11_g
+ N_VDD_XI39/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI4/MM2 N_XI39/XI4/NET34_XI39/XI4/MM2_d N_XI39/XI4/NET33_XI39/XI4/MM2_g
+ N_VSS_XI39/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI4/MM3 N_XI39/XI4/NET33_XI39/XI4/MM3_d N_WL<74>_XI39/XI4/MM3_g
+ N_BLN<11>_XI39/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI4/MM0 N_XI39/XI4/NET34_XI39/XI4/MM0_d N_WL<74>_XI39/XI4/MM0_g
+ N_BL<11>_XI39/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI4/MM1 N_XI39/XI4/NET33_XI39/XI4/MM1_d N_XI39/XI4/NET34_XI39/XI4/MM1_g
+ N_VSS_XI39/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI4/MM9 N_XI39/XI4/NET36_XI39/XI4/MM9_d N_WL<75>_XI39/XI4/MM9_g
+ N_BL<11>_XI39/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI4/MM6 N_XI39/XI4/NET35_XI39/XI4/MM6_d N_XI39/XI4/NET36_XI39/XI4/MM6_g
+ N_VSS_XI39/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI4/MM7 N_XI39/XI4/NET36_XI39/XI4/MM7_d N_XI39/XI4/NET35_XI39/XI4/MM7_g
+ N_VSS_XI39/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI4/MM8 N_XI39/XI4/NET35_XI39/XI4/MM8_d N_WL<75>_XI39/XI4/MM8_g
+ N_BLN<11>_XI39/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI4/MM5 N_XI39/XI4/NET34_XI39/XI4/MM5_d N_XI39/XI4/NET33_XI39/XI4/MM5_g
+ N_VDD_XI39/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI4/MM4 N_XI39/XI4/NET33_XI39/XI4/MM4_d N_XI39/XI4/NET34_XI39/XI4/MM4_g
+ N_VDD_XI39/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI4/MM10 N_XI39/XI4/NET35_XI39/XI4/MM10_d N_XI39/XI4/NET36_XI39/XI4/MM10_g
+ N_VDD_XI39/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI4/MM11 N_XI39/XI4/NET36_XI39/XI4/MM11_d N_XI39/XI4/NET35_XI39/XI4/MM11_g
+ N_VDD_XI39/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI5/MM2 N_XI39/XI5/NET34_XI39/XI5/MM2_d N_XI39/XI5/NET33_XI39/XI5/MM2_g
+ N_VSS_XI39/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI5/MM3 N_XI39/XI5/NET33_XI39/XI5/MM3_d N_WL<74>_XI39/XI5/MM3_g
+ N_BLN<10>_XI39/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI5/MM0 N_XI39/XI5/NET34_XI39/XI5/MM0_d N_WL<74>_XI39/XI5/MM0_g
+ N_BL<10>_XI39/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI5/MM1 N_XI39/XI5/NET33_XI39/XI5/MM1_d N_XI39/XI5/NET34_XI39/XI5/MM1_g
+ N_VSS_XI39/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI5/MM9 N_XI39/XI5/NET36_XI39/XI5/MM9_d N_WL<75>_XI39/XI5/MM9_g
+ N_BL<10>_XI39/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI5/MM6 N_XI39/XI5/NET35_XI39/XI5/MM6_d N_XI39/XI5/NET36_XI39/XI5/MM6_g
+ N_VSS_XI39/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI5/MM7 N_XI39/XI5/NET36_XI39/XI5/MM7_d N_XI39/XI5/NET35_XI39/XI5/MM7_g
+ N_VSS_XI39/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI5/MM8 N_XI39/XI5/NET35_XI39/XI5/MM8_d N_WL<75>_XI39/XI5/MM8_g
+ N_BLN<10>_XI39/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI5/MM5 N_XI39/XI5/NET34_XI39/XI5/MM5_d N_XI39/XI5/NET33_XI39/XI5/MM5_g
+ N_VDD_XI39/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI5/MM4 N_XI39/XI5/NET33_XI39/XI5/MM4_d N_XI39/XI5/NET34_XI39/XI5/MM4_g
+ N_VDD_XI39/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI5/MM10 N_XI39/XI5/NET35_XI39/XI5/MM10_d N_XI39/XI5/NET36_XI39/XI5/MM10_g
+ N_VDD_XI39/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI5/MM11 N_XI39/XI5/NET36_XI39/XI5/MM11_d N_XI39/XI5/NET35_XI39/XI5/MM11_g
+ N_VDD_XI39/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI6/MM2 N_XI39/XI6/NET34_XI39/XI6/MM2_d N_XI39/XI6/NET33_XI39/XI6/MM2_g
+ N_VSS_XI39/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM3 N_XI39/XI6/NET33_XI39/XI6/MM3_d N_WL<74>_XI39/XI6/MM3_g
+ N_BLN<9>_XI39/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM0 N_XI39/XI6/NET34_XI39/XI6/MM0_d N_WL<74>_XI39/XI6/MM0_g
+ N_BL<9>_XI39/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM1 N_XI39/XI6/NET33_XI39/XI6/MM1_d N_XI39/XI6/NET34_XI39/XI6/MM1_g
+ N_VSS_XI39/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM9 N_XI39/XI6/NET36_XI39/XI6/MM9_d N_WL<75>_XI39/XI6/MM9_g
+ N_BL<9>_XI39/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM6 N_XI39/XI6/NET35_XI39/XI6/MM6_d N_XI39/XI6/NET36_XI39/XI6/MM6_g
+ N_VSS_XI39/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM7 N_XI39/XI6/NET36_XI39/XI6/MM7_d N_XI39/XI6/NET35_XI39/XI6/MM7_g
+ N_VSS_XI39/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM8 N_XI39/XI6/NET35_XI39/XI6/MM8_d N_WL<75>_XI39/XI6/MM8_g
+ N_BLN<9>_XI39/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI6/MM5 N_XI39/XI6/NET34_XI39/XI6/MM5_d N_XI39/XI6/NET33_XI39/XI6/MM5_g
+ N_VDD_XI39/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI6/MM4 N_XI39/XI6/NET33_XI39/XI6/MM4_d N_XI39/XI6/NET34_XI39/XI6/MM4_g
+ N_VDD_XI39/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI6/MM10 N_XI39/XI6/NET35_XI39/XI6/MM10_d N_XI39/XI6/NET36_XI39/XI6/MM10_g
+ N_VDD_XI39/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI6/MM11 N_XI39/XI6/NET36_XI39/XI6/MM11_d N_XI39/XI6/NET35_XI39/XI6/MM11_g
+ N_VDD_XI39/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI7/MM2 N_XI39/XI7/NET34_XI39/XI7/MM2_d N_XI39/XI7/NET33_XI39/XI7/MM2_g
+ N_VSS_XI39/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM3 N_XI39/XI7/NET33_XI39/XI7/MM3_d N_WL<74>_XI39/XI7/MM3_g
+ N_BLN<8>_XI39/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM0 N_XI39/XI7/NET34_XI39/XI7/MM0_d N_WL<74>_XI39/XI7/MM0_g
+ N_BL<8>_XI39/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM1 N_XI39/XI7/NET33_XI39/XI7/MM1_d N_XI39/XI7/NET34_XI39/XI7/MM1_g
+ N_VSS_XI39/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM9 N_XI39/XI7/NET36_XI39/XI7/MM9_d N_WL<75>_XI39/XI7/MM9_g
+ N_BL<8>_XI39/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM6 N_XI39/XI7/NET35_XI39/XI7/MM6_d N_XI39/XI7/NET36_XI39/XI7/MM6_g
+ N_VSS_XI39/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM7 N_XI39/XI7/NET36_XI39/XI7/MM7_d N_XI39/XI7/NET35_XI39/XI7/MM7_g
+ N_VSS_XI39/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM8 N_XI39/XI7/NET35_XI39/XI7/MM8_d N_WL<75>_XI39/XI7/MM8_g
+ N_BLN<8>_XI39/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI7/MM5 N_XI39/XI7/NET34_XI39/XI7/MM5_d N_XI39/XI7/NET33_XI39/XI7/MM5_g
+ N_VDD_XI39/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI7/MM4 N_XI39/XI7/NET33_XI39/XI7/MM4_d N_XI39/XI7/NET34_XI39/XI7/MM4_g
+ N_VDD_XI39/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI7/MM10 N_XI39/XI7/NET35_XI39/XI7/MM10_d N_XI39/XI7/NET36_XI39/XI7/MM10_g
+ N_VDD_XI39/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI7/MM11 N_XI39/XI7/NET36_XI39/XI7/MM11_d N_XI39/XI7/NET35_XI39/XI7/MM11_g
+ N_VDD_XI39/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI8/MM2 N_XI39/XI8/NET34_XI39/XI8/MM2_d N_XI39/XI8/NET33_XI39/XI8/MM2_g
+ N_VSS_XI39/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM3 N_XI39/XI8/NET33_XI39/XI8/MM3_d N_WL<74>_XI39/XI8/MM3_g
+ N_BLN<7>_XI39/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM0 N_XI39/XI8/NET34_XI39/XI8/MM0_d N_WL<74>_XI39/XI8/MM0_g
+ N_BL<7>_XI39/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM1 N_XI39/XI8/NET33_XI39/XI8/MM1_d N_XI39/XI8/NET34_XI39/XI8/MM1_g
+ N_VSS_XI39/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM9 N_XI39/XI8/NET36_XI39/XI8/MM9_d N_WL<75>_XI39/XI8/MM9_g
+ N_BL<7>_XI39/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM6 N_XI39/XI8/NET35_XI39/XI8/MM6_d N_XI39/XI8/NET36_XI39/XI8/MM6_g
+ N_VSS_XI39/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM7 N_XI39/XI8/NET36_XI39/XI8/MM7_d N_XI39/XI8/NET35_XI39/XI8/MM7_g
+ N_VSS_XI39/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM8 N_XI39/XI8/NET35_XI39/XI8/MM8_d N_WL<75>_XI39/XI8/MM8_g
+ N_BLN<7>_XI39/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI8/MM5 N_XI39/XI8/NET34_XI39/XI8/MM5_d N_XI39/XI8/NET33_XI39/XI8/MM5_g
+ N_VDD_XI39/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI8/MM4 N_XI39/XI8/NET33_XI39/XI8/MM4_d N_XI39/XI8/NET34_XI39/XI8/MM4_g
+ N_VDD_XI39/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI8/MM10 N_XI39/XI8/NET35_XI39/XI8/MM10_d N_XI39/XI8/NET36_XI39/XI8/MM10_g
+ N_VDD_XI39/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI8/MM11 N_XI39/XI8/NET36_XI39/XI8/MM11_d N_XI39/XI8/NET35_XI39/XI8/MM11_g
+ N_VDD_XI39/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI9/MM2 N_XI39/XI9/NET34_XI39/XI9/MM2_d N_XI39/XI9/NET33_XI39/XI9/MM2_g
+ N_VSS_XI39/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM3 N_XI39/XI9/NET33_XI39/XI9/MM3_d N_WL<74>_XI39/XI9/MM3_g
+ N_BLN<6>_XI39/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM0 N_XI39/XI9/NET34_XI39/XI9/MM0_d N_WL<74>_XI39/XI9/MM0_g
+ N_BL<6>_XI39/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM1 N_XI39/XI9/NET33_XI39/XI9/MM1_d N_XI39/XI9/NET34_XI39/XI9/MM1_g
+ N_VSS_XI39/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM9 N_XI39/XI9/NET36_XI39/XI9/MM9_d N_WL<75>_XI39/XI9/MM9_g
+ N_BL<6>_XI39/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM6 N_XI39/XI9/NET35_XI39/XI9/MM6_d N_XI39/XI9/NET36_XI39/XI9/MM6_g
+ N_VSS_XI39/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM7 N_XI39/XI9/NET36_XI39/XI9/MM7_d N_XI39/XI9/NET35_XI39/XI9/MM7_g
+ N_VSS_XI39/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM8 N_XI39/XI9/NET35_XI39/XI9/MM8_d N_WL<75>_XI39/XI9/MM8_g
+ N_BLN<6>_XI39/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI9/MM5 N_XI39/XI9/NET34_XI39/XI9/MM5_d N_XI39/XI9/NET33_XI39/XI9/MM5_g
+ N_VDD_XI39/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI9/MM4 N_XI39/XI9/NET33_XI39/XI9/MM4_d N_XI39/XI9/NET34_XI39/XI9/MM4_g
+ N_VDD_XI39/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI9/MM10 N_XI39/XI9/NET35_XI39/XI9/MM10_d N_XI39/XI9/NET36_XI39/XI9/MM10_g
+ N_VDD_XI39/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI9/MM11 N_XI39/XI9/NET36_XI39/XI9/MM11_d N_XI39/XI9/NET35_XI39/XI9/MM11_g
+ N_VDD_XI39/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI10/MM2 N_XI39/XI10/NET34_XI39/XI10/MM2_d
+ N_XI39/XI10/NET33_XI39/XI10/MM2_g N_VSS_XI39/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI10/MM3 N_XI39/XI10/NET33_XI39/XI10/MM3_d N_WL<74>_XI39/XI10/MM3_g
+ N_BLN<5>_XI39/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI10/MM0 N_XI39/XI10/NET34_XI39/XI10/MM0_d N_WL<74>_XI39/XI10/MM0_g
+ N_BL<5>_XI39/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI10/MM1 N_XI39/XI10/NET33_XI39/XI10/MM1_d
+ N_XI39/XI10/NET34_XI39/XI10/MM1_g N_VSS_XI39/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI10/MM9 N_XI39/XI10/NET36_XI39/XI10/MM9_d N_WL<75>_XI39/XI10/MM9_g
+ N_BL<5>_XI39/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI10/MM6 N_XI39/XI10/NET35_XI39/XI10/MM6_d
+ N_XI39/XI10/NET36_XI39/XI10/MM6_g N_VSS_XI39/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI10/MM7 N_XI39/XI10/NET36_XI39/XI10/MM7_d
+ N_XI39/XI10/NET35_XI39/XI10/MM7_g N_VSS_XI39/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI10/MM8 N_XI39/XI10/NET35_XI39/XI10/MM8_d N_WL<75>_XI39/XI10/MM8_g
+ N_BLN<5>_XI39/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI10/MM5 N_XI39/XI10/NET34_XI39/XI10/MM5_d
+ N_XI39/XI10/NET33_XI39/XI10/MM5_g N_VDD_XI39/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI10/MM4 N_XI39/XI10/NET33_XI39/XI10/MM4_d
+ N_XI39/XI10/NET34_XI39/XI10/MM4_g N_VDD_XI39/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI10/MM10 N_XI39/XI10/NET35_XI39/XI10/MM10_d
+ N_XI39/XI10/NET36_XI39/XI10/MM10_g N_VDD_XI39/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI10/MM11 N_XI39/XI10/NET36_XI39/XI10/MM11_d
+ N_XI39/XI10/NET35_XI39/XI10/MM11_g N_VDD_XI39/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI11/MM2 N_XI39/XI11/NET34_XI39/XI11/MM2_d
+ N_XI39/XI11/NET33_XI39/XI11/MM2_g N_VSS_XI39/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI11/MM3 N_XI39/XI11/NET33_XI39/XI11/MM3_d N_WL<74>_XI39/XI11/MM3_g
+ N_BLN<4>_XI39/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI11/MM0 N_XI39/XI11/NET34_XI39/XI11/MM0_d N_WL<74>_XI39/XI11/MM0_g
+ N_BL<4>_XI39/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI11/MM1 N_XI39/XI11/NET33_XI39/XI11/MM1_d
+ N_XI39/XI11/NET34_XI39/XI11/MM1_g N_VSS_XI39/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI11/MM9 N_XI39/XI11/NET36_XI39/XI11/MM9_d N_WL<75>_XI39/XI11/MM9_g
+ N_BL<4>_XI39/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI11/MM6 N_XI39/XI11/NET35_XI39/XI11/MM6_d
+ N_XI39/XI11/NET36_XI39/XI11/MM6_g N_VSS_XI39/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI11/MM7 N_XI39/XI11/NET36_XI39/XI11/MM7_d
+ N_XI39/XI11/NET35_XI39/XI11/MM7_g N_VSS_XI39/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI11/MM8 N_XI39/XI11/NET35_XI39/XI11/MM8_d N_WL<75>_XI39/XI11/MM8_g
+ N_BLN<4>_XI39/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI11/MM5 N_XI39/XI11/NET34_XI39/XI11/MM5_d
+ N_XI39/XI11/NET33_XI39/XI11/MM5_g N_VDD_XI39/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI11/MM4 N_XI39/XI11/NET33_XI39/XI11/MM4_d
+ N_XI39/XI11/NET34_XI39/XI11/MM4_g N_VDD_XI39/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI11/MM10 N_XI39/XI11/NET35_XI39/XI11/MM10_d
+ N_XI39/XI11/NET36_XI39/XI11/MM10_g N_VDD_XI39/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI11/MM11 N_XI39/XI11/NET36_XI39/XI11/MM11_d
+ N_XI39/XI11/NET35_XI39/XI11/MM11_g N_VDD_XI39/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI12/MM2 N_XI39/XI12/NET34_XI39/XI12/MM2_d
+ N_XI39/XI12/NET33_XI39/XI12/MM2_g N_VSS_XI39/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI12/MM3 N_XI39/XI12/NET33_XI39/XI12/MM3_d N_WL<74>_XI39/XI12/MM3_g
+ N_BLN<3>_XI39/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI12/MM0 N_XI39/XI12/NET34_XI39/XI12/MM0_d N_WL<74>_XI39/XI12/MM0_g
+ N_BL<3>_XI39/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI12/MM1 N_XI39/XI12/NET33_XI39/XI12/MM1_d
+ N_XI39/XI12/NET34_XI39/XI12/MM1_g N_VSS_XI39/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI12/MM9 N_XI39/XI12/NET36_XI39/XI12/MM9_d N_WL<75>_XI39/XI12/MM9_g
+ N_BL<3>_XI39/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI12/MM6 N_XI39/XI12/NET35_XI39/XI12/MM6_d
+ N_XI39/XI12/NET36_XI39/XI12/MM6_g N_VSS_XI39/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI12/MM7 N_XI39/XI12/NET36_XI39/XI12/MM7_d
+ N_XI39/XI12/NET35_XI39/XI12/MM7_g N_VSS_XI39/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI12/MM8 N_XI39/XI12/NET35_XI39/XI12/MM8_d N_WL<75>_XI39/XI12/MM8_g
+ N_BLN<3>_XI39/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI12/MM5 N_XI39/XI12/NET34_XI39/XI12/MM5_d
+ N_XI39/XI12/NET33_XI39/XI12/MM5_g N_VDD_XI39/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI12/MM4 N_XI39/XI12/NET33_XI39/XI12/MM4_d
+ N_XI39/XI12/NET34_XI39/XI12/MM4_g N_VDD_XI39/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI12/MM10 N_XI39/XI12/NET35_XI39/XI12/MM10_d
+ N_XI39/XI12/NET36_XI39/XI12/MM10_g N_VDD_XI39/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI12/MM11 N_XI39/XI12/NET36_XI39/XI12/MM11_d
+ N_XI39/XI12/NET35_XI39/XI12/MM11_g N_VDD_XI39/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI13/MM2 N_XI39/XI13/NET34_XI39/XI13/MM2_d
+ N_XI39/XI13/NET33_XI39/XI13/MM2_g N_VSS_XI39/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI13/MM3 N_XI39/XI13/NET33_XI39/XI13/MM3_d N_WL<74>_XI39/XI13/MM3_g
+ N_BLN<2>_XI39/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI13/MM0 N_XI39/XI13/NET34_XI39/XI13/MM0_d N_WL<74>_XI39/XI13/MM0_g
+ N_BL<2>_XI39/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI13/MM1 N_XI39/XI13/NET33_XI39/XI13/MM1_d
+ N_XI39/XI13/NET34_XI39/XI13/MM1_g N_VSS_XI39/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI13/MM9 N_XI39/XI13/NET36_XI39/XI13/MM9_d N_WL<75>_XI39/XI13/MM9_g
+ N_BL<2>_XI39/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI13/MM6 N_XI39/XI13/NET35_XI39/XI13/MM6_d
+ N_XI39/XI13/NET36_XI39/XI13/MM6_g N_VSS_XI39/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI13/MM7 N_XI39/XI13/NET36_XI39/XI13/MM7_d
+ N_XI39/XI13/NET35_XI39/XI13/MM7_g N_VSS_XI39/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI13/MM8 N_XI39/XI13/NET35_XI39/XI13/MM8_d N_WL<75>_XI39/XI13/MM8_g
+ N_BLN<2>_XI39/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI13/MM5 N_XI39/XI13/NET34_XI39/XI13/MM5_d
+ N_XI39/XI13/NET33_XI39/XI13/MM5_g N_VDD_XI39/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI13/MM4 N_XI39/XI13/NET33_XI39/XI13/MM4_d
+ N_XI39/XI13/NET34_XI39/XI13/MM4_g N_VDD_XI39/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI13/MM10 N_XI39/XI13/NET35_XI39/XI13/MM10_d
+ N_XI39/XI13/NET36_XI39/XI13/MM10_g N_VDD_XI39/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI13/MM11 N_XI39/XI13/NET36_XI39/XI13/MM11_d
+ N_XI39/XI13/NET35_XI39/XI13/MM11_g N_VDD_XI39/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI14/MM2 N_XI39/XI14/NET34_XI39/XI14/MM2_d
+ N_XI39/XI14/NET33_XI39/XI14/MM2_g N_VSS_XI39/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI14/MM3 N_XI39/XI14/NET33_XI39/XI14/MM3_d N_WL<74>_XI39/XI14/MM3_g
+ N_BLN<1>_XI39/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI14/MM0 N_XI39/XI14/NET34_XI39/XI14/MM0_d N_WL<74>_XI39/XI14/MM0_g
+ N_BL<1>_XI39/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI14/MM1 N_XI39/XI14/NET33_XI39/XI14/MM1_d
+ N_XI39/XI14/NET34_XI39/XI14/MM1_g N_VSS_XI39/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI14/MM9 N_XI39/XI14/NET36_XI39/XI14/MM9_d N_WL<75>_XI39/XI14/MM9_g
+ N_BL<1>_XI39/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI14/MM6 N_XI39/XI14/NET35_XI39/XI14/MM6_d
+ N_XI39/XI14/NET36_XI39/XI14/MM6_g N_VSS_XI39/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI14/MM7 N_XI39/XI14/NET36_XI39/XI14/MM7_d
+ N_XI39/XI14/NET35_XI39/XI14/MM7_g N_VSS_XI39/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI14/MM8 N_XI39/XI14/NET35_XI39/XI14/MM8_d N_WL<75>_XI39/XI14/MM8_g
+ N_BLN<1>_XI39/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI14/MM5 N_XI39/XI14/NET34_XI39/XI14/MM5_d
+ N_XI39/XI14/NET33_XI39/XI14/MM5_g N_VDD_XI39/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI14/MM4 N_XI39/XI14/NET33_XI39/XI14/MM4_d
+ N_XI39/XI14/NET34_XI39/XI14/MM4_g N_VDD_XI39/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI14/MM10 N_XI39/XI14/NET35_XI39/XI14/MM10_d
+ N_XI39/XI14/NET36_XI39/XI14/MM10_g N_VDD_XI39/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI14/MM11 N_XI39/XI14/NET36_XI39/XI14/MM11_d
+ N_XI39/XI14/NET35_XI39/XI14/MM11_g N_VDD_XI39/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI15/MM2 N_XI39/XI15/NET34_XI39/XI15/MM2_d
+ N_XI39/XI15/NET33_XI39/XI15/MM2_g N_VSS_XI39/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI15/MM3 N_XI39/XI15/NET33_XI39/XI15/MM3_d N_WL<74>_XI39/XI15/MM3_g
+ N_BLN<0>_XI39/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI15/MM0 N_XI39/XI15/NET34_XI39/XI15/MM0_d N_WL<74>_XI39/XI15/MM0_g
+ N_BL<0>_XI39/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI15/MM1 N_XI39/XI15/NET33_XI39/XI15/MM1_d
+ N_XI39/XI15/NET34_XI39/XI15/MM1_g N_VSS_XI39/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI15/MM9 N_XI39/XI15/NET36_XI39/XI15/MM9_d N_WL<75>_XI39/XI15/MM9_g
+ N_BL<0>_XI39/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI15/MM6 N_XI39/XI15/NET35_XI39/XI15/MM6_d
+ N_XI39/XI15/NET36_XI39/XI15/MM6_g N_VSS_XI39/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI15/MM7 N_XI39/XI15/NET36_XI39/XI15/MM7_d
+ N_XI39/XI15/NET35_XI39/XI15/MM7_g N_VSS_XI39/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI39/XI15/MM8 N_XI39/XI15/NET35_XI39/XI15/MM8_d N_WL<75>_XI39/XI15/MM8_g
+ N_BLN<0>_XI39/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI39/XI15/MM5 N_XI39/XI15/NET34_XI39/XI15/MM5_d
+ N_XI39/XI15/NET33_XI39/XI15/MM5_g N_VDD_XI39/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI15/MM4 N_XI39/XI15/NET33_XI39/XI15/MM4_d
+ N_XI39/XI15/NET34_XI39/XI15/MM4_g N_VDD_XI39/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI15/MM10 N_XI39/XI15/NET35_XI39/XI15/MM10_d
+ N_XI39/XI15/NET36_XI39/XI15/MM10_g N_VDD_XI39/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI39/XI15/MM11 N_XI39/XI15/NET36_XI39/XI15/MM11_d
+ N_XI39/XI15/NET35_XI39/XI15/MM11_g N_VDD_XI39/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI0/MM2 N_XI40/XI0/NET34_XI40/XI0/MM2_d N_XI40/XI0/NET33_XI40/XI0/MM2_g
+ N_VSS_XI40/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI0/MM3 N_XI40/XI0/NET33_XI40/XI0/MM3_d N_WL<76>_XI40/XI0/MM3_g
+ N_BLN<15>_XI40/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI0/MM0 N_XI40/XI0/NET34_XI40/XI0/MM0_d N_WL<76>_XI40/XI0/MM0_g
+ N_BL<15>_XI40/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI0/MM1 N_XI40/XI0/NET33_XI40/XI0/MM1_d N_XI40/XI0/NET34_XI40/XI0/MM1_g
+ N_VSS_XI40/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI0/MM9 N_XI40/XI0/NET36_XI40/XI0/MM9_d N_WL<77>_XI40/XI0/MM9_g
+ N_BL<15>_XI40/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI0/MM6 N_XI40/XI0/NET35_XI40/XI0/MM6_d N_XI40/XI0/NET36_XI40/XI0/MM6_g
+ N_VSS_XI40/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI0/MM7 N_XI40/XI0/NET36_XI40/XI0/MM7_d N_XI40/XI0/NET35_XI40/XI0/MM7_g
+ N_VSS_XI40/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI0/MM8 N_XI40/XI0/NET35_XI40/XI0/MM8_d N_WL<77>_XI40/XI0/MM8_g
+ N_BLN<15>_XI40/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI0/MM5 N_XI40/XI0/NET34_XI40/XI0/MM5_d N_XI40/XI0/NET33_XI40/XI0/MM5_g
+ N_VDD_XI40/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI0/MM4 N_XI40/XI0/NET33_XI40/XI0/MM4_d N_XI40/XI0/NET34_XI40/XI0/MM4_g
+ N_VDD_XI40/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI0/MM10 N_XI40/XI0/NET35_XI40/XI0/MM10_d N_XI40/XI0/NET36_XI40/XI0/MM10_g
+ N_VDD_XI40/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI0/MM11 N_XI40/XI0/NET36_XI40/XI0/MM11_d N_XI40/XI0/NET35_XI40/XI0/MM11_g
+ N_VDD_XI40/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI1/MM2 N_XI40/XI1/NET34_XI40/XI1/MM2_d N_XI40/XI1/NET33_XI40/XI1/MM2_g
+ N_VSS_XI40/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI1/MM3 N_XI40/XI1/NET33_XI40/XI1/MM3_d N_WL<76>_XI40/XI1/MM3_g
+ N_BLN<14>_XI40/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI1/MM0 N_XI40/XI1/NET34_XI40/XI1/MM0_d N_WL<76>_XI40/XI1/MM0_g
+ N_BL<14>_XI40/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI1/MM1 N_XI40/XI1/NET33_XI40/XI1/MM1_d N_XI40/XI1/NET34_XI40/XI1/MM1_g
+ N_VSS_XI40/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI1/MM9 N_XI40/XI1/NET36_XI40/XI1/MM9_d N_WL<77>_XI40/XI1/MM9_g
+ N_BL<14>_XI40/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI1/MM6 N_XI40/XI1/NET35_XI40/XI1/MM6_d N_XI40/XI1/NET36_XI40/XI1/MM6_g
+ N_VSS_XI40/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI1/MM7 N_XI40/XI1/NET36_XI40/XI1/MM7_d N_XI40/XI1/NET35_XI40/XI1/MM7_g
+ N_VSS_XI40/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI1/MM8 N_XI40/XI1/NET35_XI40/XI1/MM8_d N_WL<77>_XI40/XI1/MM8_g
+ N_BLN<14>_XI40/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI1/MM5 N_XI40/XI1/NET34_XI40/XI1/MM5_d N_XI40/XI1/NET33_XI40/XI1/MM5_g
+ N_VDD_XI40/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI1/MM4 N_XI40/XI1/NET33_XI40/XI1/MM4_d N_XI40/XI1/NET34_XI40/XI1/MM4_g
+ N_VDD_XI40/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI1/MM10 N_XI40/XI1/NET35_XI40/XI1/MM10_d N_XI40/XI1/NET36_XI40/XI1/MM10_g
+ N_VDD_XI40/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI1/MM11 N_XI40/XI1/NET36_XI40/XI1/MM11_d N_XI40/XI1/NET35_XI40/XI1/MM11_g
+ N_VDD_XI40/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI2/MM2 N_XI40/XI2/NET34_XI40/XI2/MM2_d N_XI40/XI2/NET33_XI40/XI2/MM2_g
+ N_VSS_XI40/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI2/MM3 N_XI40/XI2/NET33_XI40/XI2/MM3_d N_WL<76>_XI40/XI2/MM3_g
+ N_BLN<13>_XI40/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI2/MM0 N_XI40/XI2/NET34_XI40/XI2/MM0_d N_WL<76>_XI40/XI2/MM0_g
+ N_BL<13>_XI40/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI2/MM1 N_XI40/XI2/NET33_XI40/XI2/MM1_d N_XI40/XI2/NET34_XI40/XI2/MM1_g
+ N_VSS_XI40/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI2/MM9 N_XI40/XI2/NET36_XI40/XI2/MM9_d N_WL<77>_XI40/XI2/MM9_g
+ N_BL<13>_XI40/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI2/MM6 N_XI40/XI2/NET35_XI40/XI2/MM6_d N_XI40/XI2/NET36_XI40/XI2/MM6_g
+ N_VSS_XI40/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI2/MM7 N_XI40/XI2/NET36_XI40/XI2/MM7_d N_XI40/XI2/NET35_XI40/XI2/MM7_g
+ N_VSS_XI40/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI2/MM8 N_XI40/XI2/NET35_XI40/XI2/MM8_d N_WL<77>_XI40/XI2/MM8_g
+ N_BLN<13>_XI40/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI2/MM5 N_XI40/XI2/NET34_XI40/XI2/MM5_d N_XI40/XI2/NET33_XI40/XI2/MM5_g
+ N_VDD_XI40/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI2/MM4 N_XI40/XI2/NET33_XI40/XI2/MM4_d N_XI40/XI2/NET34_XI40/XI2/MM4_g
+ N_VDD_XI40/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI2/MM10 N_XI40/XI2/NET35_XI40/XI2/MM10_d N_XI40/XI2/NET36_XI40/XI2/MM10_g
+ N_VDD_XI40/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI2/MM11 N_XI40/XI2/NET36_XI40/XI2/MM11_d N_XI40/XI2/NET35_XI40/XI2/MM11_g
+ N_VDD_XI40/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI3/MM2 N_XI40/XI3/NET34_XI40/XI3/MM2_d N_XI40/XI3/NET33_XI40/XI3/MM2_g
+ N_VSS_XI40/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI3/MM3 N_XI40/XI3/NET33_XI40/XI3/MM3_d N_WL<76>_XI40/XI3/MM3_g
+ N_BLN<12>_XI40/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI3/MM0 N_XI40/XI3/NET34_XI40/XI3/MM0_d N_WL<76>_XI40/XI3/MM0_g
+ N_BL<12>_XI40/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI3/MM1 N_XI40/XI3/NET33_XI40/XI3/MM1_d N_XI40/XI3/NET34_XI40/XI3/MM1_g
+ N_VSS_XI40/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI3/MM9 N_XI40/XI3/NET36_XI40/XI3/MM9_d N_WL<77>_XI40/XI3/MM9_g
+ N_BL<12>_XI40/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI3/MM6 N_XI40/XI3/NET35_XI40/XI3/MM6_d N_XI40/XI3/NET36_XI40/XI3/MM6_g
+ N_VSS_XI40/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI3/MM7 N_XI40/XI3/NET36_XI40/XI3/MM7_d N_XI40/XI3/NET35_XI40/XI3/MM7_g
+ N_VSS_XI40/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI3/MM8 N_XI40/XI3/NET35_XI40/XI3/MM8_d N_WL<77>_XI40/XI3/MM8_g
+ N_BLN<12>_XI40/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI3/MM5 N_XI40/XI3/NET34_XI40/XI3/MM5_d N_XI40/XI3/NET33_XI40/XI3/MM5_g
+ N_VDD_XI40/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI3/MM4 N_XI40/XI3/NET33_XI40/XI3/MM4_d N_XI40/XI3/NET34_XI40/XI3/MM4_g
+ N_VDD_XI40/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI3/MM10 N_XI40/XI3/NET35_XI40/XI3/MM10_d N_XI40/XI3/NET36_XI40/XI3/MM10_g
+ N_VDD_XI40/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI3/MM11 N_XI40/XI3/NET36_XI40/XI3/MM11_d N_XI40/XI3/NET35_XI40/XI3/MM11_g
+ N_VDD_XI40/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI4/MM2 N_XI40/XI4/NET34_XI40/XI4/MM2_d N_XI40/XI4/NET33_XI40/XI4/MM2_g
+ N_VSS_XI40/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI4/MM3 N_XI40/XI4/NET33_XI40/XI4/MM3_d N_WL<76>_XI40/XI4/MM3_g
+ N_BLN<11>_XI40/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI4/MM0 N_XI40/XI4/NET34_XI40/XI4/MM0_d N_WL<76>_XI40/XI4/MM0_g
+ N_BL<11>_XI40/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI4/MM1 N_XI40/XI4/NET33_XI40/XI4/MM1_d N_XI40/XI4/NET34_XI40/XI4/MM1_g
+ N_VSS_XI40/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI4/MM9 N_XI40/XI4/NET36_XI40/XI4/MM9_d N_WL<77>_XI40/XI4/MM9_g
+ N_BL<11>_XI40/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI4/MM6 N_XI40/XI4/NET35_XI40/XI4/MM6_d N_XI40/XI4/NET36_XI40/XI4/MM6_g
+ N_VSS_XI40/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI4/MM7 N_XI40/XI4/NET36_XI40/XI4/MM7_d N_XI40/XI4/NET35_XI40/XI4/MM7_g
+ N_VSS_XI40/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI4/MM8 N_XI40/XI4/NET35_XI40/XI4/MM8_d N_WL<77>_XI40/XI4/MM8_g
+ N_BLN<11>_XI40/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI4/MM5 N_XI40/XI4/NET34_XI40/XI4/MM5_d N_XI40/XI4/NET33_XI40/XI4/MM5_g
+ N_VDD_XI40/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI4/MM4 N_XI40/XI4/NET33_XI40/XI4/MM4_d N_XI40/XI4/NET34_XI40/XI4/MM4_g
+ N_VDD_XI40/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI4/MM10 N_XI40/XI4/NET35_XI40/XI4/MM10_d N_XI40/XI4/NET36_XI40/XI4/MM10_g
+ N_VDD_XI40/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI4/MM11 N_XI40/XI4/NET36_XI40/XI4/MM11_d N_XI40/XI4/NET35_XI40/XI4/MM11_g
+ N_VDD_XI40/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI5/MM2 N_XI40/XI5/NET34_XI40/XI5/MM2_d N_XI40/XI5/NET33_XI40/XI5/MM2_g
+ N_VSS_XI40/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI5/MM3 N_XI40/XI5/NET33_XI40/XI5/MM3_d N_WL<76>_XI40/XI5/MM3_g
+ N_BLN<10>_XI40/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI5/MM0 N_XI40/XI5/NET34_XI40/XI5/MM0_d N_WL<76>_XI40/XI5/MM0_g
+ N_BL<10>_XI40/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI5/MM1 N_XI40/XI5/NET33_XI40/XI5/MM1_d N_XI40/XI5/NET34_XI40/XI5/MM1_g
+ N_VSS_XI40/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI5/MM9 N_XI40/XI5/NET36_XI40/XI5/MM9_d N_WL<77>_XI40/XI5/MM9_g
+ N_BL<10>_XI40/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI5/MM6 N_XI40/XI5/NET35_XI40/XI5/MM6_d N_XI40/XI5/NET36_XI40/XI5/MM6_g
+ N_VSS_XI40/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI5/MM7 N_XI40/XI5/NET36_XI40/XI5/MM7_d N_XI40/XI5/NET35_XI40/XI5/MM7_g
+ N_VSS_XI40/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI5/MM8 N_XI40/XI5/NET35_XI40/XI5/MM8_d N_WL<77>_XI40/XI5/MM8_g
+ N_BLN<10>_XI40/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI5/MM5 N_XI40/XI5/NET34_XI40/XI5/MM5_d N_XI40/XI5/NET33_XI40/XI5/MM5_g
+ N_VDD_XI40/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI5/MM4 N_XI40/XI5/NET33_XI40/XI5/MM4_d N_XI40/XI5/NET34_XI40/XI5/MM4_g
+ N_VDD_XI40/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI5/MM10 N_XI40/XI5/NET35_XI40/XI5/MM10_d N_XI40/XI5/NET36_XI40/XI5/MM10_g
+ N_VDD_XI40/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI5/MM11 N_XI40/XI5/NET36_XI40/XI5/MM11_d N_XI40/XI5/NET35_XI40/XI5/MM11_g
+ N_VDD_XI40/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI6/MM2 N_XI40/XI6/NET34_XI40/XI6/MM2_d N_XI40/XI6/NET33_XI40/XI6/MM2_g
+ N_VSS_XI40/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM3 N_XI40/XI6/NET33_XI40/XI6/MM3_d N_WL<76>_XI40/XI6/MM3_g
+ N_BLN<9>_XI40/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM0 N_XI40/XI6/NET34_XI40/XI6/MM0_d N_WL<76>_XI40/XI6/MM0_g
+ N_BL<9>_XI40/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM1 N_XI40/XI6/NET33_XI40/XI6/MM1_d N_XI40/XI6/NET34_XI40/XI6/MM1_g
+ N_VSS_XI40/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM9 N_XI40/XI6/NET36_XI40/XI6/MM9_d N_WL<77>_XI40/XI6/MM9_g
+ N_BL<9>_XI40/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM6 N_XI40/XI6/NET35_XI40/XI6/MM6_d N_XI40/XI6/NET36_XI40/XI6/MM6_g
+ N_VSS_XI40/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM7 N_XI40/XI6/NET36_XI40/XI6/MM7_d N_XI40/XI6/NET35_XI40/XI6/MM7_g
+ N_VSS_XI40/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM8 N_XI40/XI6/NET35_XI40/XI6/MM8_d N_WL<77>_XI40/XI6/MM8_g
+ N_BLN<9>_XI40/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI6/MM5 N_XI40/XI6/NET34_XI40/XI6/MM5_d N_XI40/XI6/NET33_XI40/XI6/MM5_g
+ N_VDD_XI40/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI6/MM4 N_XI40/XI6/NET33_XI40/XI6/MM4_d N_XI40/XI6/NET34_XI40/XI6/MM4_g
+ N_VDD_XI40/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI6/MM10 N_XI40/XI6/NET35_XI40/XI6/MM10_d N_XI40/XI6/NET36_XI40/XI6/MM10_g
+ N_VDD_XI40/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI6/MM11 N_XI40/XI6/NET36_XI40/XI6/MM11_d N_XI40/XI6/NET35_XI40/XI6/MM11_g
+ N_VDD_XI40/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI7/MM2 N_XI40/XI7/NET34_XI40/XI7/MM2_d N_XI40/XI7/NET33_XI40/XI7/MM2_g
+ N_VSS_XI40/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM3 N_XI40/XI7/NET33_XI40/XI7/MM3_d N_WL<76>_XI40/XI7/MM3_g
+ N_BLN<8>_XI40/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM0 N_XI40/XI7/NET34_XI40/XI7/MM0_d N_WL<76>_XI40/XI7/MM0_g
+ N_BL<8>_XI40/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM1 N_XI40/XI7/NET33_XI40/XI7/MM1_d N_XI40/XI7/NET34_XI40/XI7/MM1_g
+ N_VSS_XI40/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM9 N_XI40/XI7/NET36_XI40/XI7/MM9_d N_WL<77>_XI40/XI7/MM9_g
+ N_BL<8>_XI40/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM6 N_XI40/XI7/NET35_XI40/XI7/MM6_d N_XI40/XI7/NET36_XI40/XI7/MM6_g
+ N_VSS_XI40/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM7 N_XI40/XI7/NET36_XI40/XI7/MM7_d N_XI40/XI7/NET35_XI40/XI7/MM7_g
+ N_VSS_XI40/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM8 N_XI40/XI7/NET35_XI40/XI7/MM8_d N_WL<77>_XI40/XI7/MM8_g
+ N_BLN<8>_XI40/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI7/MM5 N_XI40/XI7/NET34_XI40/XI7/MM5_d N_XI40/XI7/NET33_XI40/XI7/MM5_g
+ N_VDD_XI40/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI7/MM4 N_XI40/XI7/NET33_XI40/XI7/MM4_d N_XI40/XI7/NET34_XI40/XI7/MM4_g
+ N_VDD_XI40/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI7/MM10 N_XI40/XI7/NET35_XI40/XI7/MM10_d N_XI40/XI7/NET36_XI40/XI7/MM10_g
+ N_VDD_XI40/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI7/MM11 N_XI40/XI7/NET36_XI40/XI7/MM11_d N_XI40/XI7/NET35_XI40/XI7/MM11_g
+ N_VDD_XI40/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI8/MM2 N_XI40/XI8/NET34_XI40/XI8/MM2_d N_XI40/XI8/NET33_XI40/XI8/MM2_g
+ N_VSS_XI40/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM3 N_XI40/XI8/NET33_XI40/XI8/MM3_d N_WL<76>_XI40/XI8/MM3_g
+ N_BLN<7>_XI40/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM0 N_XI40/XI8/NET34_XI40/XI8/MM0_d N_WL<76>_XI40/XI8/MM0_g
+ N_BL<7>_XI40/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM1 N_XI40/XI8/NET33_XI40/XI8/MM1_d N_XI40/XI8/NET34_XI40/XI8/MM1_g
+ N_VSS_XI40/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM9 N_XI40/XI8/NET36_XI40/XI8/MM9_d N_WL<77>_XI40/XI8/MM9_g
+ N_BL<7>_XI40/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM6 N_XI40/XI8/NET35_XI40/XI8/MM6_d N_XI40/XI8/NET36_XI40/XI8/MM6_g
+ N_VSS_XI40/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM7 N_XI40/XI8/NET36_XI40/XI8/MM7_d N_XI40/XI8/NET35_XI40/XI8/MM7_g
+ N_VSS_XI40/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM8 N_XI40/XI8/NET35_XI40/XI8/MM8_d N_WL<77>_XI40/XI8/MM8_g
+ N_BLN<7>_XI40/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI8/MM5 N_XI40/XI8/NET34_XI40/XI8/MM5_d N_XI40/XI8/NET33_XI40/XI8/MM5_g
+ N_VDD_XI40/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI8/MM4 N_XI40/XI8/NET33_XI40/XI8/MM4_d N_XI40/XI8/NET34_XI40/XI8/MM4_g
+ N_VDD_XI40/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI8/MM10 N_XI40/XI8/NET35_XI40/XI8/MM10_d N_XI40/XI8/NET36_XI40/XI8/MM10_g
+ N_VDD_XI40/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI8/MM11 N_XI40/XI8/NET36_XI40/XI8/MM11_d N_XI40/XI8/NET35_XI40/XI8/MM11_g
+ N_VDD_XI40/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI9/MM2 N_XI40/XI9/NET34_XI40/XI9/MM2_d N_XI40/XI9/NET33_XI40/XI9/MM2_g
+ N_VSS_XI40/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM3 N_XI40/XI9/NET33_XI40/XI9/MM3_d N_WL<76>_XI40/XI9/MM3_g
+ N_BLN<6>_XI40/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM0 N_XI40/XI9/NET34_XI40/XI9/MM0_d N_WL<76>_XI40/XI9/MM0_g
+ N_BL<6>_XI40/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM1 N_XI40/XI9/NET33_XI40/XI9/MM1_d N_XI40/XI9/NET34_XI40/XI9/MM1_g
+ N_VSS_XI40/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM9 N_XI40/XI9/NET36_XI40/XI9/MM9_d N_WL<77>_XI40/XI9/MM9_g
+ N_BL<6>_XI40/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM6 N_XI40/XI9/NET35_XI40/XI9/MM6_d N_XI40/XI9/NET36_XI40/XI9/MM6_g
+ N_VSS_XI40/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM7 N_XI40/XI9/NET36_XI40/XI9/MM7_d N_XI40/XI9/NET35_XI40/XI9/MM7_g
+ N_VSS_XI40/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM8 N_XI40/XI9/NET35_XI40/XI9/MM8_d N_WL<77>_XI40/XI9/MM8_g
+ N_BLN<6>_XI40/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI9/MM5 N_XI40/XI9/NET34_XI40/XI9/MM5_d N_XI40/XI9/NET33_XI40/XI9/MM5_g
+ N_VDD_XI40/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI9/MM4 N_XI40/XI9/NET33_XI40/XI9/MM4_d N_XI40/XI9/NET34_XI40/XI9/MM4_g
+ N_VDD_XI40/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI9/MM10 N_XI40/XI9/NET35_XI40/XI9/MM10_d N_XI40/XI9/NET36_XI40/XI9/MM10_g
+ N_VDD_XI40/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI9/MM11 N_XI40/XI9/NET36_XI40/XI9/MM11_d N_XI40/XI9/NET35_XI40/XI9/MM11_g
+ N_VDD_XI40/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI10/MM2 N_XI40/XI10/NET34_XI40/XI10/MM2_d
+ N_XI40/XI10/NET33_XI40/XI10/MM2_g N_VSS_XI40/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI10/MM3 N_XI40/XI10/NET33_XI40/XI10/MM3_d N_WL<76>_XI40/XI10/MM3_g
+ N_BLN<5>_XI40/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI10/MM0 N_XI40/XI10/NET34_XI40/XI10/MM0_d N_WL<76>_XI40/XI10/MM0_g
+ N_BL<5>_XI40/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI10/MM1 N_XI40/XI10/NET33_XI40/XI10/MM1_d
+ N_XI40/XI10/NET34_XI40/XI10/MM1_g N_VSS_XI40/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI10/MM9 N_XI40/XI10/NET36_XI40/XI10/MM9_d N_WL<77>_XI40/XI10/MM9_g
+ N_BL<5>_XI40/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI10/MM6 N_XI40/XI10/NET35_XI40/XI10/MM6_d
+ N_XI40/XI10/NET36_XI40/XI10/MM6_g N_VSS_XI40/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI10/MM7 N_XI40/XI10/NET36_XI40/XI10/MM7_d
+ N_XI40/XI10/NET35_XI40/XI10/MM7_g N_VSS_XI40/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI10/MM8 N_XI40/XI10/NET35_XI40/XI10/MM8_d N_WL<77>_XI40/XI10/MM8_g
+ N_BLN<5>_XI40/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI10/MM5 N_XI40/XI10/NET34_XI40/XI10/MM5_d
+ N_XI40/XI10/NET33_XI40/XI10/MM5_g N_VDD_XI40/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI10/MM4 N_XI40/XI10/NET33_XI40/XI10/MM4_d
+ N_XI40/XI10/NET34_XI40/XI10/MM4_g N_VDD_XI40/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI10/MM10 N_XI40/XI10/NET35_XI40/XI10/MM10_d
+ N_XI40/XI10/NET36_XI40/XI10/MM10_g N_VDD_XI40/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI10/MM11 N_XI40/XI10/NET36_XI40/XI10/MM11_d
+ N_XI40/XI10/NET35_XI40/XI10/MM11_g N_VDD_XI40/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI11/MM2 N_XI40/XI11/NET34_XI40/XI11/MM2_d
+ N_XI40/XI11/NET33_XI40/XI11/MM2_g N_VSS_XI40/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI11/MM3 N_XI40/XI11/NET33_XI40/XI11/MM3_d N_WL<76>_XI40/XI11/MM3_g
+ N_BLN<4>_XI40/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI11/MM0 N_XI40/XI11/NET34_XI40/XI11/MM0_d N_WL<76>_XI40/XI11/MM0_g
+ N_BL<4>_XI40/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI11/MM1 N_XI40/XI11/NET33_XI40/XI11/MM1_d
+ N_XI40/XI11/NET34_XI40/XI11/MM1_g N_VSS_XI40/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI11/MM9 N_XI40/XI11/NET36_XI40/XI11/MM9_d N_WL<77>_XI40/XI11/MM9_g
+ N_BL<4>_XI40/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI11/MM6 N_XI40/XI11/NET35_XI40/XI11/MM6_d
+ N_XI40/XI11/NET36_XI40/XI11/MM6_g N_VSS_XI40/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI11/MM7 N_XI40/XI11/NET36_XI40/XI11/MM7_d
+ N_XI40/XI11/NET35_XI40/XI11/MM7_g N_VSS_XI40/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI11/MM8 N_XI40/XI11/NET35_XI40/XI11/MM8_d N_WL<77>_XI40/XI11/MM8_g
+ N_BLN<4>_XI40/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI11/MM5 N_XI40/XI11/NET34_XI40/XI11/MM5_d
+ N_XI40/XI11/NET33_XI40/XI11/MM5_g N_VDD_XI40/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI11/MM4 N_XI40/XI11/NET33_XI40/XI11/MM4_d
+ N_XI40/XI11/NET34_XI40/XI11/MM4_g N_VDD_XI40/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI11/MM10 N_XI40/XI11/NET35_XI40/XI11/MM10_d
+ N_XI40/XI11/NET36_XI40/XI11/MM10_g N_VDD_XI40/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI11/MM11 N_XI40/XI11/NET36_XI40/XI11/MM11_d
+ N_XI40/XI11/NET35_XI40/XI11/MM11_g N_VDD_XI40/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI12/MM2 N_XI40/XI12/NET34_XI40/XI12/MM2_d
+ N_XI40/XI12/NET33_XI40/XI12/MM2_g N_VSS_XI40/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI12/MM3 N_XI40/XI12/NET33_XI40/XI12/MM3_d N_WL<76>_XI40/XI12/MM3_g
+ N_BLN<3>_XI40/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI12/MM0 N_XI40/XI12/NET34_XI40/XI12/MM0_d N_WL<76>_XI40/XI12/MM0_g
+ N_BL<3>_XI40/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI12/MM1 N_XI40/XI12/NET33_XI40/XI12/MM1_d
+ N_XI40/XI12/NET34_XI40/XI12/MM1_g N_VSS_XI40/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI12/MM9 N_XI40/XI12/NET36_XI40/XI12/MM9_d N_WL<77>_XI40/XI12/MM9_g
+ N_BL<3>_XI40/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI12/MM6 N_XI40/XI12/NET35_XI40/XI12/MM6_d
+ N_XI40/XI12/NET36_XI40/XI12/MM6_g N_VSS_XI40/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI12/MM7 N_XI40/XI12/NET36_XI40/XI12/MM7_d
+ N_XI40/XI12/NET35_XI40/XI12/MM7_g N_VSS_XI40/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI12/MM8 N_XI40/XI12/NET35_XI40/XI12/MM8_d N_WL<77>_XI40/XI12/MM8_g
+ N_BLN<3>_XI40/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI12/MM5 N_XI40/XI12/NET34_XI40/XI12/MM5_d
+ N_XI40/XI12/NET33_XI40/XI12/MM5_g N_VDD_XI40/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI12/MM4 N_XI40/XI12/NET33_XI40/XI12/MM4_d
+ N_XI40/XI12/NET34_XI40/XI12/MM4_g N_VDD_XI40/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI12/MM10 N_XI40/XI12/NET35_XI40/XI12/MM10_d
+ N_XI40/XI12/NET36_XI40/XI12/MM10_g N_VDD_XI40/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI12/MM11 N_XI40/XI12/NET36_XI40/XI12/MM11_d
+ N_XI40/XI12/NET35_XI40/XI12/MM11_g N_VDD_XI40/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI13/MM2 N_XI40/XI13/NET34_XI40/XI13/MM2_d
+ N_XI40/XI13/NET33_XI40/XI13/MM2_g N_VSS_XI40/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI13/MM3 N_XI40/XI13/NET33_XI40/XI13/MM3_d N_WL<76>_XI40/XI13/MM3_g
+ N_BLN<2>_XI40/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI13/MM0 N_XI40/XI13/NET34_XI40/XI13/MM0_d N_WL<76>_XI40/XI13/MM0_g
+ N_BL<2>_XI40/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI13/MM1 N_XI40/XI13/NET33_XI40/XI13/MM1_d
+ N_XI40/XI13/NET34_XI40/XI13/MM1_g N_VSS_XI40/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI13/MM9 N_XI40/XI13/NET36_XI40/XI13/MM9_d N_WL<77>_XI40/XI13/MM9_g
+ N_BL<2>_XI40/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI13/MM6 N_XI40/XI13/NET35_XI40/XI13/MM6_d
+ N_XI40/XI13/NET36_XI40/XI13/MM6_g N_VSS_XI40/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI13/MM7 N_XI40/XI13/NET36_XI40/XI13/MM7_d
+ N_XI40/XI13/NET35_XI40/XI13/MM7_g N_VSS_XI40/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI13/MM8 N_XI40/XI13/NET35_XI40/XI13/MM8_d N_WL<77>_XI40/XI13/MM8_g
+ N_BLN<2>_XI40/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI13/MM5 N_XI40/XI13/NET34_XI40/XI13/MM5_d
+ N_XI40/XI13/NET33_XI40/XI13/MM5_g N_VDD_XI40/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI13/MM4 N_XI40/XI13/NET33_XI40/XI13/MM4_d
+ N_XI40/XI13/NET34_XI40/XI13/MM4_g N_VDD_XI40/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI13/MM10 N_XI40/XI13/NET35_XI40/XI13/MM10_d
+ N_XI40/XI13/NET36_XI40/XI13/MM10_g N_VDD_XI40/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI13/MM11 N_XI40/XI13/NET36_XI40/XI13/MM11_d
+ N_XI40/XI13/NET35_XI40/XI13/MM11_g N_VDD_XI40/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI14/MM2 N_XI40/XI14/NET34_XI40/XI14/MM2_d
+ N_XI40/XI14/NET33_XI40/XI14/MM2_g N_VSS_XI40/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI14/MM3 N_XI40/XI14/NET33_XI40/XI14/MM3_d N_WL<76>_XI40/XI14/MM3_g
+ N_BLN<1>_XI40/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI14/MM0 N_XI40/XI14/NET34_XI40/XI14/MM0_d N_WL<76>_XI40/XI14/MM0_g
+ N_BL<1>_XI40/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI14/MM1 N_XI40/XI14/NET33_XI40/XI14/MM1_d
+ N_XI40/XI14/NET34_XI40/XI14/MM1_g N_VSS_XI40/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI14/MM9 N_XI40/XI14/NET36_XI40/XI14/MM9_d N_WL<77>_XI40/XI14/MM9_g
+ N_BL<1>_XI40/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI14/MM6 N_XI40/XI14/NET35_XI40/XI14/MM6_d
+ N_XI40/XI14/NET36_XI40/XI14/MM6_g N_VSS_XI40/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI14/MM7 N_XI40/XI14/NET36_XI40/XI14/MM7_d
+ N_XI40/XI14/NET35_XI40/XI14/MM7_g N_VSS_XI40/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI14/MM8 N_XI40/XI14/NET35_XI40/XI14/MM8_d N_WL<77>_XI40/XI14/MM8_g
+ N_BLN<1>_XI40/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI14/MM5 N_XI40/XI14/NET34_XI40/XI14/MM5_d
+ N_XI40/XI14/NET33_XI40/XI14/MM5_g N_VDD_XI40/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI14/MM4 N_XI40/XI14/NET33_XI40/XI14/MM4_d
+ N_XI40/XI14/NET34_XI40/XI14/MM4_g N_VDD_XI40/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI14/MM10 N_XI40/XI14/NET35_XI40/XI14/MM10_d
+ N_XI40/XI14/NET36_XI40/XI14/MM10_g N_VDD_XI40/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI14/MM11 N_XI40/XI14/NET36_XI40/XI14/MM11_d
+ N_XI40/XI14/NET35_XI40/XI14/MM11_g N_VDD_XI40/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI15/MM2 N_XI40/XI15/NET34_XI40/XI15/MM2_d
+ N_XI40/XI15/NET33_XI40/XI15/MM2_g N_VSS_XI40/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI15/MM3 N_XI40/XI15/NET33_XI40/XI15/MM3_d N_WL<76>_XI40/XI15/MM3_g
+ N_BLN<0>_XI40/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI15/MM0 N_XI40/XI15/NET34_XI40/XI15/MM0_d N_WL<76>_XI40/XI15/MM0_g
+ N_BL<0>_XI40/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI15/MM1 N_XI40/XI15/NET33_XI40/XI15/MM1_d
+ N_XI40/XI15/NET34_XI40/XI15/MM1_g N_VSS_XI40/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI15/MM9 N_XI40/XI15/NET36_XI40/XI15/MM9_d N_WL<77>_XI40/XI15/MM9_g
+ N_BL<0>_XI40/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI15/MM6 N_XI40/XI15/NET35_XI40/XI15/MM6_d
+ N_XI40/XI15/NET36_XI40/XI15/MM6_g N_VSS_XI40/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI15/MM7 N_XI40/XI15/NET36_XI40/XI15/MM7_d
+ N_XI40/XI15/NET35_XI40/XI15/MM7_g N_VSS_XI40/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI40/XI15/MM8 N_XI40/XI15/NET35_XI40/XI15/MM8_d N_WL<77>_XI40/XI15/MM8_g
+ N_BLN<0>_XI40/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI40/XI15/MM5 N_XI40/XI15/NET34_XI40/XI15/MM5_d
+ N_XI40/XI15/NET33_XI40/XI15/MM5_g N_VDD_XI40/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI15/MM4 N_XI40/XI15/NET33_XI40/XI15/MM4_d
+ N_XI40/XI15/NET34_XI40/XI15/MM4_g N_VDD_XI40/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI15/MM10 N_XI40/XI15/NET35_XI40/XI15/MM10_d
+ N_XI40/XI15/NET36_XI40/XI15/MM10_g N_VDD_XI40/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI40/XI15/MM11 N_XI40/XI15/NET36_XI40/XI15/MM11_d
+ N_XI40/XI15/NET35_XI40/XI15/MM11_g N_VDD_XI40/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI0/MM2 N_XI41/XI0/NET34_XI41/XI0/MM2_d N_XI41/XI0/NET33_XI41/XI0/MM2_g
+ N_VSS_XI41/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI0/MM3 N_XI41/XI0/NET33_XI41/XI0/MM3_d N_WL<78>_XI41/XI0/MM3_g
+ N_BLN<15>_XI41/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI0/MM0 N_XI41/XI0/NET34_XI41/XI0/MM0_d N_WL<78>_XI41/XI0/MM0_g
+ N_BL<15>_XI41/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI0/MM1 N_XI41/XI0/NET33_XI41/XI0/MM1_d N_XI41/XI0/NET34_XI41/XI0/MM1_g
+ N_VSS_XI41/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI0/MM9 N_XI41/XI0/NET36_XI41/XI0/MM9_d N_WL<79>_XI41/XI0/MM9_g
+ N_BL<15>_XI41/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI0/MM6 N_XI41/XI0/NET35_XI41/XI0/MM6_d N_XI41/XI0/NET36_XI41/XI0/MM6_g
+ N_VSS_XI41/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI0/MM7 N_XI41/XI0/NET36_XI41/XI0/MM7_d N_XI41/XI0/NET35_XI41/XI0/MM7_g
+ N_VSS_XI41/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI0/MM8 N_XI41/XI0/NET35_XI41/XI0/MM8_d N_WL<79>_XI41/XI0/MM8_g
+ N_BLN<15>_XI41/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI0/MM5 N_XI41/XI0/NET34_XI41/XI0/MM5_d N_XI41/XI0/NET33_XI41/XI0/MM5_g
+ N_VDD_XI41/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI0/MM4 N_XI41/XI0/NET33_XI41/XI0/MM4_d N_XI41/XI0/NET34_XI41/XI0/MM4_g
+ N_VDD_XI41/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI0/MM10 N_XI41/XI0/NET35_XI41/XI0/MM10_d N_XI41/XI0/NET36_XI41/XI0/MM10_g
+ N_VDD_XI41/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI0/MM11 N_XI41/XI0/NET36_XI41/XI0/MM11_d N_XI41/XI0/NET35_XI41/XI0/MM11_g
+ N_VDD_XI41/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI1/MM2 N_XI41/XI1/NET34_XI41/XI1/MM2_d N_XI41/XI1/NET33_XI41/XI1/MM2_g
+ N_VSS_XI41/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI1/MM3 N_XI41/XI1/NET33_XI41/XI1/MM3_d N_WL<78>_XI41/XI1/MM3_g
+ N_BLN<14>_XI41/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI1/MM0 N_XI41/XI1/NET34_XI41/XI1/MM0_d N_WL<78>_XI41/XI1/MM0_g
+ N_BL<14>_XI41/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI1/MM1 N_XI41/XI1/NET33_XI41/XI1/MM1_d N_XI41/XI1/NET34_XI41/XI1/MM1_g
+ N_VSS_XI41/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI1/MM9 N_XI41/XI1/NET36_XI41/XI1/MM9_d N_WL<79>_XI41/XI1/MM9_g
+ N_BL<14>_XI41/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI1/MM6 N_XI41/XI1/NET35_XI41/XI1/MM6_d N_XI41/XI1/NET36_XI41/XI1/MM6_g
+ N_VSS_XI41/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI1/MM7 N_XI41/XI1/NET36_XI41/XI1/MM7_d N_XI41/XI1/NET35_XI41/XI1/MM7_g
+ N_VSS_XI41/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI1/MM8 N_XI41/XI1/NET35_XI41/XI1/MM8_d N_WL<79>_XI41/XI1/MM8_g
+ N_BLN<14>_XI41/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI1/MM5 N_XI41/XI1/NET34_XI41/XI1/MM5_d N_XI41/XI1/NET33_XI41/XI1/MM5_g
+ N_VDD_XI41/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI1/MM4 N_XI41/XI1/NET33_XI41/XI1/MM4_d N_XI41/XI1/NET34_XI41/XI1/MM4_g
+ N_VDD_XI41/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI1/MM10 N_XI41/XI1/NET35_XI41/XI1/MM10_d N_XI41/XI1/NET36_XI41/XI1/MM10_g
+ N_VDD_XI41/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI1/MM11 N_XI41/XI1/NET36_XI41/XI1/MM11_d N_XI41/XI1/NET35_XI41/XI1/MM11_g
+ N_VDD_XI41/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI2/MM2 N_XI41/XI2/NET34_XI41/XI2/MM2_d N_XI41/XI2/NET33_XI41/XI2/MM2_g
+ N_VSS_XI41/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI2/MM3 N_XI41/XI2/NET33_XI41/XI2/MM3_d N_WL<78>_XI41/XI2/MM3_g
+ N_BLN<13>_XI41/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI2/MM0 N_XI41/XI2/NET34_XI41/XI2/MM0_d N_WL<78>_XI41/XI2/MM0_g
+ N_BL<13>_XI41/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI2/MM1 N_XI41/XI2/NET33_XI41/XI2/MM1_d N_XI41/XI2/NET34_XI41/XI2/MM1_g
+ N_VSS_XI41/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI2/MM9 N_XI41/XI2/NET36_XI41/XI2/MM9_d N_WL<79>_XI41/XI2/MM9_g
+ N_BL<13>_XI41/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI2/MM6 N_XI41/XI2/NET35_XI41/XI2/MM6_d N_XI41/XI2/NET36_XI41/XI2/MM6_g
+ N_VSS_XI41/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI2/MM7 N_XI41/XI2/NET36_XI41/XI2/MM7_d N_XI41/XI2/NET35_XI41/XI2/MM7_g
+ N_VSS_XI41/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI2/MM8 N_XI41/XI2/NET35_XI41/XI2/MM8_d N_WL<79>_XI41/XI2/MM8_g
+ N_BLN<13>_XI41/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI2/MM5 N_XI41/XI2/NET34_XI41/XI2/MM5_d N_XI41/XI2/NET33_XI41/XI2/MM5_g
+ N_VDD_XI41/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI2/MM4 N_XI41/XI2/NET33_XI41/XI2/MM4_d N_XI41/XI2/NET34_XI41/XI2/MM4_g
+ N_VDD_XI41/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI2/MM10 N_XI41/XI2/NET35_XI41/XI2/MM10_d N_XI41/XI2/NET36_XI41/XI2/MM10_g
+ N_VDD_XI41/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI2/MM11 N_XI41/XI2/NET36_XI41/XI2/MM11_d N_XI41/XI2/NET35_XI41/XI2/MM11_g
+ N_VDD_XI41/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI3/MM2 N_XI41/XI3/NET34_XI41/XI3/MM2_d N_XI41/XI3/NET33_XI41/XI3/MM2_g
+ N_VSS_XI41/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI3/MM3 N_XI41/XI3/NET33_XI41/XI3/MM3_d N_WL<78>_XI41/XI3/MM3_g
+ N_BLN<12>_XI41/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI3/MM0 N_XI41/XI3/NET34_XI41/XI3/MM0_d N_WL<78>_XI41/XI3/MM0_g
+ N_BL<12>_XI41/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI3/MM1 N_XI41/XI3/NET33_XI41/XI3/MM1_d N_XI41/XI3/NET34_XI41/XI3/MM1_g
+ N_VSS_XI41/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI3/MM9 N_XI41/XI3/NET36_XI41/XI3/MM9_d N_WL<79>_XI41/XI3/MM9_g
+ N_BL<12>_XI41/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI3/MM6 N_XI41/XI3/NET35_XI41/XI3/MM6_d N_XI41/XI3/NET36_XI41/XI3/MM6_g
+ N_VSS_XI41/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI3/MM7 N_XI41/XI3/NET36_XI41/XI3/MM7_d N_XI41/XI3/NET35_XI41/XI3/MM7_g
+ N_VSS_XI41/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI3/MM8 N_XI41/XI3/NET35_XI41/XI3/MM8_d N_WL<79>_XI41/XI3/MM8_g
+ N_BLN<12>_XI41/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI3/MM5 N_XI41/XI3/NET34_XI41/XI3/MM5_d N_XI41/XI3/NET33_XI41/XI3/MM5_g
+ N_VDD_XI41/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI3/MM4 N_XI41/XI3/NET33_XI41/XI3/MM4_d N_XI41/XI3/NET34_XI41/XI3/MM4_g
+ N_VDD_XI41/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI3/MM10 N_XI41/XI3/NET35_XI41/XI3/MM10_d N_XI41/XI3/NET36_XI41/XI3/MM10_g
+ N_VDD_XI41/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI3/MM11 N_XI41/XI3/NET36_XI41/XI3/MM11_d N_XI41/XI3/NET35_XI41/XI3/MM11_g
+ N_VDD_XI41/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI4/MM2 N_XI41/XI4/NET34_XI41/XI4/MM2_d N_XI41/XI4/NET33_XI41/XI4/MM2_g
+ N_VSS_XI41/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI4/MM3 N_XI41/XI4/NET33_XI41/XI4/MM3_d N_WL<78>_XI41/XI4/MM3_g
+ N_BLN<11>_XI41/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI4/MM0 N_XI41/XI4/NET34_XI41/XI4/MM0_d N_WL<78>_XI41/XI4/MM0_g
+ N_BL<11>_XI41/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI4/MM1 N_XI41/XI4/NET33_XI41/XI4/MM1_d N_XI41/XI4/NET34_XI41/XI4/MM1_g
+ N_VSS_XI41/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI4/MM9 N_XI41/XI4/NET36_XI41/XI4/MM9_d N_WL<79>_XI41/XI4/MM9_g
+ N_BL<11>_XI41/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI4/MM6 N_XI41/XI4/NET35_XI41/XI4/MM6_d N_XI41/XI4/NET36_XI41/XI4/MM6_g
+ N_VSS_XI41/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI4/MM7 N_XI41/XI4/NET36_XI41/XI4/MM7_d N_XI41/XI4/NET35_XI41/XI4/MM7_g
+ N_VSS_XI41/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI4/MM8 N_XI41/XI4/NET35_XI41/XI4/MM8_d N_WL<79>_XI41/XI4/MM8_g
+ N_BLN<11>_XI41/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI4/MM5 N_XI41/XI4/NET34_XI41/XI4/MM5_d N_XI41/XI4/NET33_XI41/XI4/MM5_g
+ N_VDD_XI41/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI4/MM4 N_XI41/XI4/NET33_XI41/XI4/MM4_d N_XI41/XI4/NET34_XI41/XI4/MM4_g
+ N_VDD_XI41/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI4/MM10 N_XI41/XI4/NET35_XI41/XI4/MM10_d N_XI41/XI4/NET36_XI41/XI4/MM10_g
+ N_VDD_XI41/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI4/MM11 N_XI41/XI4/NET36_XI41/XI4/MM11_d N_XI41/XI4/NET35_XI41/XI4/MM11_g
+ N_VDD_XI41/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI5/MM2 N_XI41/XI5/NET34_XI41/XI5/MM2_d N_XI41/XI5/NET33_XI41/XI5/MM2_g
+ N_VSS_XI41/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI5/MM3 N_XI41/XI5/NET33_XI41/XI5/MM3_d N_WL<78>_XI41/XI5/MM3_g
+ N_BLN<10>_XI41/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI5/MM0 N_XI41/XI5/NET34_XI41/XI5/MM0_d N_WL<78>_XI41/XI5/MM0_g
+ N_BL<10>_XI41/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI5/MM1 N_XI41/XI5/NET33_XI41/XI5/MM1_d N_XI41/XI5/NET34_XI41/XI5/MM1_g
+ N_VSS_XI41/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI5/MM9 N_XI41/XI5/NET36_XI41/XI5/MM9_d N_WL<79>_XI41/XI5/MM9_g
+ N_BL<10>_XI41/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI5/MM6 N_XI41/XI5/NET35_XI41/XI5/MM6_d N_XI41/XI5/NET36_XI41/XI5/MM6_g
+ N_VSS_XI41/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI5/MM7 N_XI41/XI5/NET36_XI41/XI5/MM7_d N_XI41/XI5/NET35_XI41/XI5/MM7_g
+ N_VSS_XI41/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI5/MM8 N_XI41/XI5/NET35_XI41/XI5/MM8_d N_WL<79>_XI41/XI5/MM8_g
+ N_BLN<10>_XI41/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI5/MM5 N_XI41/XI5/NET34_XI41/XI5/MM5_d N_XI41/XI5/NET33_XI41/XI5/MM5_g
+ N_VDD_XI41/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI5/MM4 N_XI41/XI5/NET33_XI41/XI5/MM4_d N_XI41/XI5/NET34_XI41/XI5/MM4_g
+ N_VDD_XI41/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI5/MM10 N_XI41/XI5/NET35_XI41/XI5/MM10_d N_XI41/XI5/NET36_XI41/XI5/MM10_g
+ N_VDD_XI41/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI5/MM11 N_XI41/XI5/NET36_XI41/XI5/MM11_d N_XI41/XI5/NET35_XI41/XI5/MM11_g
+ N_VDD_XI41/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI6/MM2 N_XI41/XI6/NET34_XI41/XI6/MM2_d N_XI41/XI6/NET33_XI41/XI6/MM2_g
+ N_VSS_XI41/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM3 N_XI41/XI6/NET33_XI41/XI6/MM3_d N_WL<78>_XI41/XI6/MM3_g
+ N_BLN<9>_XI41/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM0 N_XI41/XI6/NET34_XI41/XI6/MM0_d N_WL<78>_XI41/XI6/MM0_g
+ N_BL<9>_XI41/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM1 N_XI41/XI6/NET33_XI41/XI6/MM1_d N_XI41/XI6/NET34_XI41/XI6/MM1_g
+ N_VSS_XI41/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM9 N_XI41/XI6/NET36_XI41/XI6/MM9_d N_WL<79>_XI41/XI6/MM9_g
+ N_BL<9>_XI41/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM6 N_XI41/XI6/NET35_XI41/XI6/MM6_d N_XI41/XI6/NET36_XI41/XI6/MM6_g
+ N_VSS_XI41/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM7 N_XI41/XI6/NET36_XI41/XI6/MM7_d N_XI41/XI6/NET35_XI41/XI6/MM7_g
+ N_VSS_XI41/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM8 N_XI41/XI6/NET35_XI41/XI6/MM8_d N_WL<79>_XI41/XI6/MM8_g
+ N_BLN<9>_XI41/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI6/MM5 N_XI41/XI6/NET34_XI41/XI6/MM5_d N_XI41/XI6/NET33_XI41/XI6/MM5_g
+ N_VDD_XI41/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI6/MM4 N_XI41/XI6/NET33_XI41/XI6/MM4_d N_XI41/XI6/NET34_XI41/XI6/MM4_g
+ N_VDD_XI41/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI6/MM10 N_XI41/XI6/NET35_XI41/XI6/MM10_d N_XI41/XI6/NET36_XI41/XI6/MM10_g
+ N_VDD_XI41/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI6/MM11 N_XI41/XI6/NET36_XI41/XI6/MM11_d N_XI41/XI6/NET35_XI41/XI6/MM11_g
+ N_VDD_XI41/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI7/MM2 N_XI41/XI7/NET34_XI41/XI7/MM2_d N_XI41/XI7/NET33_XI41/XI7/MM2_g
+ N_VSS_XI41/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM3 N_XI41/XI7/NET33_XI41/XI7/MM3_d N_WL<78>_XI41/XI7/MM3_g
+ N_BLN<8>_XI41/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM0 N_XI41/XI7/NET34_XI41/XI7/MM0_d N_WL<78>_XI41/XI7/MM0_g
+ N_BL<8>_XI41/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM1 N_XI41/XI7/NET33_XI41/XI7/MM1_d N_XI41/XI7/NET34_XI41/XI7/MM1_g
+ N_VSS_XI41/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM9 N_XI41/XI7/NET36_XI41/XI7/MM9_d N_WL<79>_XI41/XI7/MM9_g
+ N_BL<8>_XI41/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM6 N_XI41/XI7/NET35_XI41/XI7/MM6_d N_XI41/XI7/NET36_XI41/XI7/MM6_g
+ N_VSS_XI41/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM7 N_XI41/XI7/NET36_XI41/XI7/MM7_d N_XI41/XI7/NET35_XI41/XI7/MM7_g
+ N_VSS_XI41/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM8 N_XI41/XI7/NET35_XI41/XI7/MM8_d N_WL<79>_XI41/XI7/MM8_g
+ N_BLN<8>_XI41/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI7/MM5 N_XI41/XI7/NET34_XI41/XI7/MM5_d N_XI41/XI7/NET33_XI41/XI7/MM5_g
+ N_VDD_XI41/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI7/MM4 N_XI41/XI7/NET33_XI41/XI7/MM4_d N_XI41/XI7/NET34_XI41/XI7/MM4_g
+ N_VDD_XI41/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI7/MM10 N_XI41/XI7/NET35_XI41/XI7/MM10_d N_XI41/XI7/NET36_XI41/XI7/MM10_g
+ N_VDD_XI41/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI7/MM11 N_XI41/XI7/NET36_XI41/XI7/MM11_d N_XI41/XI7/NET35_XI41/XI7/MM11_g
+ N_VDD_XI41/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI8/MM2 N_XI41/XI8/NET34_XI41/XI8/MM2_d N_XI41/XI8/NET33_XI41/XI8/MM2_g
+ N_VSS_XI41/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM3 N_XI41/XI8/NET33_XI41/XI8/MM3_d N_WL<78>_XI41/XI8/MM3_g
+ N_BLN<7>_XI41/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM0 N_XI41/XI8/NET34_XI41/XI8/MM0_d N_WL<78>_XI41/XI8/MM0_g
+ N_BL<7>_XI41/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM1 N_XI41/XI8/NET33_XI41/XI8/MM1_d N_XI41/XI8/NET34_XI41/XI8/MM1_g
+ N_VSS_XI41/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM9 N_XI41/XI8/NET36_XI41/XI8/MM9_d N_WL<79>_XI41/XI8/MM9_g
+ N_BL<7>_XI41/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM6 N_XI41/XI8/NET35_XI41/XI8/MM6_d N_XI41/XI8/NET36_XI41/XI8/MM6_g
+ N_VSS_XI41/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM7 N_XI41/XI8/NET36_XI41/XI8/MM7_d N_XI41/XI8/NET35_XI41/XI8/MM7_g
+ N_VSS_XI41/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM8 N_XI41/XI8/NET35_XI41/XI8/MM8_d N_WL<79>_XI41/XI8/MM8_g
+ N_BLN<7>_XI41/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI8/MM5 N_XI41/XI8/NET34_XI41/XI8/MM5_d N_XI41/XI8/NET33_XI41/XI8/MM5_g
+ N_VDD_XI41/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI8/MM4 N_XI41/XI8/NET33_XI41/XI8/MM4_d N_XI41/XI8/NET34_XI41/XI8/MM4_g
+ N_VDD_XI41/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI8/MM10 N_XI41/XI8/NET35_XI41/XI8/MM10_d N_XI41/XI8/NET36_XI41/XI8/MM10_g
+ N_VDD_XI41/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI8/MM11 N_XI41/XI8/NET36_XI41/XI8/MM11_d N_XI41/XI8/NET35_XI41/XI8/MM11_g
+ N_VDD_XI41/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI9/MM2 N_XI41/XI9/NET34_XI41/XI9/MM2_d N_XI41/XI9/NET33_XI41/XI9/MM2_g
+ N_VSS_XI41/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM3 N_XI41/XI9/NET33_XI41/XI9/MM3_d N_WL<78>_XI41/XI9/MM3_g
+ N_BLN<6>_XI41/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM0 N_XI41/XI9/NET34_XI41/XI9/MM0_d N_WL<78>_XI41/XI9/MM0_g
+ N_BL<6>_XI41/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM1 N_XI41/XI9/NET33_XI41/XI9/MM1_d N_XI41/XI9/NET34_XI41/XI9/MM1_g
+ N_VSS_XI41/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM9 N_XI41/XI9/NET36_XI41/XI9/MM9_d N_WL<79>_XI41/XI9/MM9_g
+ N_BL<6>_XI41/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM6 N_XI41/XI9/NET35_XI41/XI9/MM6_d N_XI41/XI9/NET36_XI41/XI9/MM6_g
+ N_VSS_XI41/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM7 N_XI41/XI9/NET36_XI41/XI9/MM7_d N_XI41/XI9/NET35_XI41/XI9/MM7_g
+ N_VSS_XI41/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM8 N_XI41/XI9/NET35_XI41/XI9/MM8_d N_WL<79>_XI41/XI9/MM8_g
+ N_BLN<6>_XI41/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI9/MM5 N_XI41/XI9/NET34_XI41/XI9/MM5_d N_XI41/XI9/NET33_XI41/XI9/MM5_g
+ N_VDD_XI41/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI9/MM4 N_XI41/XI9/NET33_XI41/XI9/MM4_d N_XI41/XI9/NET34_XI41/XI9/MM4_g
+ N_VDD_XI41/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI9/MM10 N_XI41/XI9/NET35_XI41/XI9/MM10_d N_XI41/XI9/NET36_XI41/XI9/MM10_g
+ N_VDD_XI41/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI9/MM11 N_XI41/XI9/NET36_XI41/XI9/MM11_d N_XI41/XI9/NET35_XI41/XI9/MM11_g
+ N_VDD_XI41/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI10/MM2 N_XI41/XI10/NET34_XI41/XI10/MM2_d
+ N_XI41/XI10/NET33_XI41/XI10/MM2_g N_VSS_XI41/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI10/MM3 N_XI41/XI10/NET33_XI41/XI10/MM3_d N_WL<78>_XI41/XI10/MM3_g
+ N_BLN<5>_XI41/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI10/MM0 N_XI41/XI10/NET34_XI41/XI10/MM0_d N_WL<78>_XI41/XI10/MM0_g
+ N_BL<5>_XI41/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI10/MM1 N_XI41/XI10/NET33_XI41/XI10/MM1_d
+ N_XI41/XI10/NET34_XI41/XI10/MM1_g N_VSS_XI41/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI10/MM9 N_XI41/XI10/NET36_XI41/XI10/MM9_d N_WL<79>_XI41/XI10/MM9_g
+ N_BL<5>_XI41/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI10/MM6 N_XI41/XI10/NET35_XI41/XI10/MM6_d
+ N_XI41/XI10/NET36_XI41/XI10/MM6_g N_VSS_XI41/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI10/MM7 N_XI41/XI10/NET36_XI41/XI10/MM7_d
+ N_XI41/XI10/NET35_XI41/XI10/MM7_g N_VSS_XI41/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI10/MM8 N_XI41/XI10/NET35_XI41/XI10/MM8_d N_WL<79>_XI41/XI10/MM8_g
+ N_BLN<5>_XI41/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI10/MM5 N_XI41/XI10/NET34_XI41/XI10/MM5_d
+ N_XI41/XI10/NET33_XI41/XI10/MM5_g N_VDD_XI41/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI10/MM4 N_XI41/XI10/NET33_XI41/XI10/MM4_d
+ N_XI41/XI10/NET34_XI41/XI10/MM4_g N_VDD_XI41/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI10/MM10 N_XI41/XI10/NET35_XI41/XI10/MM10_d
+ N_XI41/XI10/NET36_XI41/XI10/MM10_g N_VDD_XI41/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI10/MM11 N_XI41/XI10/NET36_XI41/XI10/MM11_d
+ N_XI41/XI10/NET35_XI41/XI10/MM11_g N_VDD_XI41/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI11/MM2 N_XI41/XI11/NET34_XI41/XI11/MM2_d
+ N_XI41/XI11/NET33_XI41/XI11/MM2_g N_VSS_XI41/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI11/MM3 N_XI41/XI11/NET33_XI41/XI11/MM3_d N_WL<78>_XI41/XI11/MM3_g
+ N_BLN<4>_XI41/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI11/MM0 N_XI41/XI11/NET34_XI41/XI11/MM0_d N_WL<78>_XI41/XI11/MM0_g
+ N_BL<4>_XI41/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI11/MM1 N_XI41/XI11/NET33_XI41/XI11/MM1_d
+ N_XI41/XI11/NET34_XI41/XI11/MM1_g N_VSS_XI41/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI11/MM9 N_XI41/XI11/NET36_XI41/XI11/MM9_d N_WL<79>_XI41/XI11/MM9_g
+ N_BL<4>_XI41/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI11/MM6 N_XI41/XI11/NET35_XI41/XI11/MM6_d
+ N_XI41/XI11/NET36_XI41/XI11/MM6_g N_VSS_XI41/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI11/MM7 N_XI41/XI11/NET36_XI41/XI11/MM7_d
+ N_XI41/XI11/NET35_XI41/XI11/MM7_g N_VSS_XI41/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI11/MM8 N_XI41/XI11/NET35_XI41/XI11/MM8_d N_WL<79>_XI41/XI11/MM8_g
+ N_BLN<4>_XI41/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI11/MM5 N_XI41/XI11/NET34_XI41/XI11/MM5_d
+ N_XI41/XI11/NET33_XI41/XI11/MM5_g N_VDD_XI41/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI11/MM4 N_XI41/XI11/NET33_XI41/XI11/MM4_d
+ N_XI41/XI11/NET34_XI41/XI11/MM4_g N_VDD_XI41/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI11/MM10 N_XI41/XI11/NET35_XI41/XI11/MM10_d
+ N_XI41/XI11/NET36_XI41/XI11/MM10_g N_VDD_XI41/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI11/MM11 N_XI41/XI11/NET36_XI41/XI11/MM11_d
+ N_XI41/XI11/NET35_XI41/XI11/MM11_g N_VDD_XI41/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI12/MM2 N_XI41/XI12/NET34_XI41/XI12/MM2_d
+ N_XI41/XI12/NET33_XI41/XI12/MM2_g N_VSS_XI41/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI12/MM3 N_XI41/XI12/NET33_XI41/XI12/MM3_d N_WL<78>_XI41/XI12/MM3_g
+ N_BLN<3>_XI41/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI12/MM0 N_XI41/XI12/NET34_XI41/XI12/MM0_d N_WL<78>_XI41/XI12/MM0_g
+ N_BL<3>_XI41/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI12/MM1 N_XI41/XI12/NET33_XI41/XI12/MM1_d
+ N_XI41/XI12/NET34_XI41/XI12/MM1_g N_VSS_XI41/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI12/MM9 N_XI41/XI12/NET36_XI41/XI12/MM9_d N_WL<79>_XI41/XI12/MM9_g
+ N_BL<3>_XI41/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI12/MM6 N_XI41/XI12/NET35_XI41/XI12/MM6_d
+ N_XI41/XI12/NET36_XI41/XI12/MM6_g N_VSS_XI41/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI12/MM7 N_XI41/XI12/NET36_XI41/XI12/MM7_d
+ N_XI41/XI12/NET35_XI41/XI12/MM7_g N_VSS_XI41/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI12/MM8 N_XI41/XI12/NET35_XI41/XI12/MM8_d N_WL<79>_XI41/XI12/MM8_g
+ N_BLN<3>_XI41/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI12/MM5 N_XI41/XI12/NET34_XI41/XI12/MM5_d
+ N_XI41/XI12/NET33_XI41/XI12/MM5_g N_VDD_XI41/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI12/MM4 N_XI41/XI12/NET33_XI41/XI12/MM4_d
+ N_XI41/XI12/NET34_XI41/XI12/MM4_g N_VDD_XI41/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI12/MM10 N_XI41/XI12/NET35_XI41/XI12/MM10_d
+ N_XI41/XI12/NET36_XI41/XI12/MM10_g N_VDD_XI41/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI12/MM11 N_XI41/XI12/NET36_XI41/XI12/MM11_d
+ N_XI41/XI12/NET35_XI41/XI12/MM11_g N_VDD_XI41/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI13/MM2 N_XI41/XI13/NET34_XI41/XI13/MM2_d
+ N_XI41/XI13/NET33_XI41/XI13/MM2_g N_VSS_XI41/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI13/MM3 N_XI41/XI13/NET33_XI41/XI13/MM3_d N_WL<78>_XI41/XI13/MM3_g
+ N_BLN<2>_XI41/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI13/MM0 N_XI41/XI13/NET34_XI41/XI13/MM0_d N_WL<78>_XI41/XI13/MM0_g
+ N_BL<2>_XI41/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI13/MM1 N_XI41/XI13/NET33_XI41/XI13/MM1_d
+ N_XI41/XI13/NET34_XI41/XI13/MM1_g N_VSS_XI41/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI13/MM9 N_XI41/XI13/NET36_XI41/XI13/MM9_d N_WL<79>_XI41/XI13/MM9_g
+ N_BL<2>_XI41/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI13/MM6 N_XI41/XI13/NET35_XI41/XI13/MM6_d
+ N_XI41/XI13/NET36_XI41/XI13/MM6_g N_VSS_XI41/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI13/MM7 N_XI41/XI13/NET36_XI41/XI13/MM7_d
+ N_XI41/XI13/NET35_XI41/XI13/MM7_g N_VSS_XI41/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI13/MM8 N_XI41/XI13/NET35_XI41/XI13/MM8_d N_WL<79>_XI41/XI13/MM8_g
+ N_BLN<2>_XI41/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI13/MM5 N_XI41/XI13/NET34_XI41/XI13/MM5_d
+ N_XI41/XI13/NET33_XI41/XI13/MM5_g N_VDD_XI41/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI13/MM4 N_XI41/XI13/NET33_XI41/XI13/MM4_d
+ N_XI41/XI13/NET34_XI41/XI13/MM4_g N_VDD_XI41/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI13/MM10 N_XI41/XI13/NET35_XI41/XI13/MM10_d
+ N_XI41/XI13/NET36_XI41/XI13/MM10_g N_VDD_XI41/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI13/MM11 N_XI41/XI13/NET36_XI41/XI13/MM11_d
+ N_XI41/XI13/NET35_XI41/XI13/MM11_g N_VDD_XI41/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI14/MM2 N_XI41/XI14/NET34_XI41/XI14/MM2_d
+ N_XI41/XI14/NET33_XI41/XI14/MM2_g N_VSS_XI41/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI14/MM3 N_XI41/XI14/NET33_XI41/XI14/MM3_d N_WL<78>_XI41/XI14/MM3_g
+ N_BLN<1>_XI41/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI14/MM0 N_XI41/XI14/NET34_XI41/XI14/MM0_d N_WL<78>_XI41/XI14/MM0_g
+ N_BL<1>_XI41/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI14/MM1 N_XI41/XI14/NET33_XI41/XI14/MM1_d
+ N_XI41/XI14/NET34_XI41/XI14/MM1_g N_VSS_XI41/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI14/MM9 N_XI41/XI14/NET36_XI41/XI14/MM9_d N_WL<79>_XI41/XI14/MM9_g
+ N_BL<1>_XI41/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI14/MM6 N_XI41/XI14/NET35_XI41/XI14/MM6_d
+ N_XI41/XI14/NET36_XI41/XI14/MM6_g N_VSS_XI41/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI14/MM7 N_XI41/XI14/NET36_XI41/XI14/MM7_d
+ N_XI41/XI14/NET35_XI41/XI14/MM7_g N_VSS_XI41/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI14/MM8 N_XI41/XI14/NET35_XI41/XI14/MM8_d N_WL<79>_XI41/XI14/MM8_g
+ N_BLN<1>_XI41/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI14/MM5 N_XI41/XI14/NET34_XI41/XI14/MM5_d
+ N_XI41/XI14/NET33_XI41/XI14/MM5_g N_VDD_XI41/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI14/MM4 N_XI41/XI14/NET33_XI41/XI14/MM4_d
+ N_XI41/XI14/NET34_XI41/XI14/MM4_g N_VDD_XI41/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI14/MM10 N_XI41/XI14/NET35_XI41/XI14/MM10_d
+ N_XI41/XI14/NET36_XI41/XI14/MM10_g N_VDD_XI41/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI14/MM11 N_XI41/XI14/NET36_XI41/XI14/MM11_d
+ N_XI41/XI14/NET35_XI41/XI14/MM11_g N_VDD_XI41/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI15/MM2 N_XI41/XI15/NET34_XI41/XI15/MM2_d
+ N_XI41/XI15/NET33_XI41/XI15/MM2_g N_VSS_XI41/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI15/MM3 N_XI41/XI15/NET33_XI41/XI15/MM3_d N_WL<78>_XI41/XI15/MM3_g
+ N_BLN<0>_XI41/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI15/MM0 N_XI41/XI15/NET34_XI41/XI15/MM0_d N_WL<78>_XI41/XI15/MM0_g
+ N_BL<0>_XI41/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI15/MM1 N_XI41/XI15/NET33_XI41/XI15/MM1_d
+ N_XI41/XI15/NET34_XI41/XI15/MM1_g N_VSS_XI41/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI15/MM9 N_XI41/XI15/NET36_XI41/XI15/MM9_d N_WL<79>_XI41/XI15/MM9_g
+ N_BL<0>_XI41/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI15/MM6 N_XI41/XI15/NET35_XI41/XI15/MM6_d
+ N_XI41/XI15/NET36_XI41/XI15/MM6_g N_VSS_XI41/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI15/MM7 N_XI41/XI15/NET36_XI41/XI15/MM7_d
+ N_XI41/XI15/NET35_XI41/XI15/MM7_g N_VSS_XI41/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI41/XI15/MM8 N_XI41/XI15/NET35_XI41/XI15/MM8_d N_WL<79>_XI41/XI15/MM8_g
+ N_BLN<0>_XI41/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI41/XI15/MM5 N_XI41/XI15/NET34_XI41/XI15/MM5_d
+ N_XI41/XI15/NET33_XI41/XI15/MM5_g N_VDD_XI41/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI15/MM4 N_XI41/XI15/NET33_XI41/XI15/MM4_d
+ N_XI41/XI15/NET34_XI41/XI15/MM4_g N_VDD_XI41/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI15/MM10 N_XI41/XI15/NET35_XI41/XI15/MM10_d
+ N_XI41/XI15/NET36_XI41/XI15/MM10_g N_VDD_XI41/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI41/XI15/MM11 N_XI41/XI15/NET36_XI41/XI15/MM11_d
+ N_XI41/XI15/NET35_XI41/XI15/MM11_g N_VDD_XI41/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI0/MM2 N_XI42/XI0/NET34_XI42/XI0/MM2_d N_XI42/XI0/NET33_XI42/XI0/MM2_g
+ N_VSS_XI42/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI0/MM3 N_XI42/XI0/NET33_XI42/XI0/MM3_d N_WL<80>_XI42/XI0/MM3_g
+ N_BLN<15>_XI42/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI0/MM0 N_XI42/XI0/NET34_XI42/XI0/MM0_d N_WL<80>_XI42/XI0/MM0_g
+ N_BL<15>_XI42/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI0/MM1 N_XI42/XI0/NET33_XI42/XI0/MM1_d N_XI42/XI0/NET34_XI42/XI0/MM1_g
+ N_VSS_XI42/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI0/MM9 N_XI42/XI0/NET36_XI42/XI0/MM9_d N_WL<81>_XI42/XI0/MM9_g
+ N_BL<15>_XI42/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI0/MM6 N_XI42/XI0/NET35_XI42/XI0/MM6_d N_XI42/XI0/NET36_XI42/XI0/MM6_g
+ N_VSS_XI42/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI0/MM7 N_XI42/XI0/NET36_XI42/XI0/MM7_d N_XI42/XI0/NET35_XI42/XI0/MM7_g
+ N_VSS_XI42/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI0/MM8 N_XI42/XI0/NET35_XI42/XI0/MM8_d N_WL<81>_XI42/XI0/MM8_g
+ N_BLN<15>_XI42/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI0/MM5 N_XI42/XI0/NET34_XI42/XI0/MM5_d N_XI42/XI0/NET33_XI42/XI0/MM5_g
+ N_VDD_XI42/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI0/MM4 N_XI42/XI0/NET33_XI42/XI0/MM4_d N_XI42/XI0/NET34_XI42/XI0/MM4_g
+ N_VDD_XI42/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI0/MM10 N_XI42/XI0/NET35_XI42/XI0/MM10_d N_XI42/XI0/NET36_XI42/XI0/MM10_g
+ N_VDD_XI42/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI0/MM11 N_XI42/XI0/NET36_XI42/XI0/MM11_d N_XI42/XI0/NET35_XI42/XI0/MM11_g
+ N_VDD_XI42/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI1/MM2 N_XI42/XI1/NET34_XI42/XI1/MM2_d N_XI42/XI1/NET33_XI42/XI1/MM2_g
+ N_VSS_XI42/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI1/MM3 N_XI42/XI1/NET33_XI42/XI1/MM3_d N_WL<80>_XI42/XI1/MM3_g
+ N_BLN<14>_XI42/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI1/MM0 N_XI42/XI1/NET34_XI42/XI1/MM0_d N_WL<80>_XI42/XI1/MM0_g
+ N_BL<14>_XI42/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI1/MM1 N_XI42/XI1/NET33_XI42/XI1/MM1_d N_XI42/XI1/NET34_XI42/XI1/MM1_g
+ N_VSS_XI42/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI1/MM9 N_XI42/XI1/NET36_XI42/XI1/MM9_d N_WL<81>_XI42/XI1/MM9_g
+ N_BL<14>_XI42/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI1/MM6 N_XI42/XI1/NET35_XI42/XI1/MM6_d N_XI42/XI1/NET36_XI42/XI1/MM6_g
+ N_VSS_XI42/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI1/MM7 N_XI42/XI1/NET36_XI42/XI1/MM7_d N_XI42/XI1/NET35_XI42/XI1/MM7_g
+ N_VSS_XI42/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI1/MM8 N_XI42/XI1/NET35_XI42/XI1/MM8_d N_WL<81>_XI42/XI1/MM8_g
+ N_BLN<14>_XI42/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI1/MM5 N_XI42/XI1/NET34_XI42/XI1/MM5_d N_XI42/XI1/NET33_XI42/XI1/MM5_g
+ N_VDD_XI42/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI1/MM4 N_XI42/XI1/NET33_XI42/XI1/MM4_d N_XI42/XI1/NET34_XI42/XI1/MM4_g
+ N_VDD_XI42/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI1/MM10 N_XI42/XI1/NET35_XI42/XI1/MM10_d N_XI42/XI1/NET36_XI42/XI1/MM10_g
+ N_VDD_XI42/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI1/MM11 N_XI42/XI1/NET36_XI42/XI1/MM11_d N_XI42/XI1/NET35_XI42/XI1/MM11_g
+ N_VDD_XI42/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI2/MM2 N_XI42/XI2/NET34_XI42/XI2/MM2_d N_XI42/XI2/NET33_XI42/XI2/MM2_g
+ N_VSS_XI42/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI2/MM3 N_XI42/XI2/NET33_XI42/XI2/MM3_d N_WL<80>_XI42/XI2/MM3_g
+ N_BLN<13>_XI42/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI2/MM0 N_XI42/XI2/NET34_XI42/XI2/MM0_d N_WL<80>_XI42/XI2/MM0_g
+ N_BL<13>_XI42/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI2/MM1 N_XI42/XI2/NET33_XI42/XI2/MM1_d N_XI42/XI2/NET34_XI42/XI2/MM1_g
+ N_VSS_XI42/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI2/MM9 N_XI42/XI2/NET36_XI42/XI2/MM9_d N_WL<81>_XI42/XI2/MM9_g
+ N_BL<13>_XI42/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI2/MM6 N_XI42/XI2/NET35_XI42/XI2/MM6_d N_XI42/XI2/NET36_XI42/XI2/MM6_g
+ N_VSS_XI42/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI2/MM7 N_XI42/XI2/NET36_XI42/XI2/MM7_d N_XI42/XI2/NET35_XI42/XI2/MM7_g
+ N_VSS_XI42/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI2/MM8 N_XI42/XI2/NET35_XI42/XI2/MM8_d N_WL<81>_XI42/XI2/MM8_g
+ N_BLN<13>_XI42/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI2/MM5 N_XI42/XI2/NET34_XI42/XI2/MM5_d N_XI42/XI2/NET33_XI42/XI2/MM5_g
+ N_VDD_XI42/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI2/MM4 N_XI42/XI2/NET33_XI42/XI2/MM4_d N_XI42/XI2/NET34_XI42/XI2/MM4_g
+ N_VDD_XI42/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI2/MM10 N_XI42/XI2/NET35_XI42/XI2/MM10_d N_XI42/XI2/NET36_XI42/XI2/MM10_g
+ N_VDD_XI42/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI2/MM11 N_XI42/XI2/NET36_XI42/XI2/MM11_d N_XI42/XI2/NET35_XI42/XI2/MM11_g
+ N_VDD_XI42/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI3/MM2 N_XI42/XI3/NET34_XI42/XI3/MM2_d N_XI42/XI3/NET33_XI42/XI3/MM2_g
+ N_VSS_XI42/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI3/MM3 N_XI42/XI3/NET33_XI42/XI3/MM3_d N_WL<80>_XI42/XI3/MM3_g
+ N_BLN<12>_XI42/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI3/MM0 N_XI42/XI3/NET34_XI42/XI3/MM0_d N_WL<80>_XI42/XI3/MM0_g
+ N_BL<12>_XI42/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI3/MM1 N_XI42/XI3/NET33_XI42/XI3/MM1_d N_XI42/XI3/NET34_XI42/XI3/MM1_g
+ N_VSS_XI42/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI3/MM9 N_XI42/XI3/NET36_XI42/XI3/MM9_d N_WL<81>_XI42/XI3/MM9_g
+ N_BL<12>_XI42/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI3/MM6 N_XI42/XI3/NET35_XI42/XI3/MM6_d N_XI42/XI3/NET36_XI42/XI3/MM6_g
+ N_VSS_XI42/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI3/MM7 N_XI42/XI3/NET36_XI42/XI3/MM7_d N_XI42/XI3/NET35_XI42/XI3/MM7_g
+ N_VSS_XI42/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI3/MM8 N_XI42/XI3/NET35_XI42/XI3/MM8_d N_WL<81>_XI42/XI3/MM8_g
+ N_BLN<12>_XI42/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI3/MM5 N_XI42/XI3/NET34_XI42/XI3/MM5_d N_XI42/XI3/NET33_XI42/XI3/MM5_g
+ N_VDD_XI42/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI3/MM4 N_XI42/XI3/NET33_XI42/XI3/MM4_d N_XI42/XI3/NET34_XI42/XI3/MM4_g
+ N_VDD_XI42/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI3/MM10 N_XI42/XI3/NET35_XI42/XI3/MM10_d N_XI42/XI3/NET36_XI42/XI3/MM10_g
+ N_VDD_XI42/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI3/MM11 N_XI42/XI3/NET36_XI42/XI3/MM11_d N_XI42/XI3/NET35_XI42/XI3/MM11_g
+ N_VDD_XI42/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI4/MM2 N_XI42/XI4/NET34_XI42/XI4/MM2_d N_XI42/XI4/NET33_XI42/XI4/MM2_g
+ N_VSS_XI42/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI4/MM3 N_XI42/XI4/NET33_XI42/XI4/MM3_d N_WL<80>_XI42/XI4/MM3_g
+ N_BLN<11>_XI42/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI4/MM0 N_XI42/XI4/NET34_XI42/XI4/MM0_d N_WL<80>_XI42/XI4/MM0_g
+ N_BL<11>_XI42/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI4/MM1 N_XI42/XI4/NET33_XI42/XI4/MM1_d N_XI42/XI4/NET34_XI42/XI4/MM1_g
+ N_VSS_XI42/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI4/MM9 N_XI42/XI4/NET36_XI42/XI4/MM9_d N_WL<81>_XI42/XI4/MM9_g
+ N_BL<11>_XI42/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI4/MM6 N_XI42/XI4/NET35_XI42/XI4/MM6_d N_XI42/XI4/NET36_XI42/XI4/MM6_g
+ N_VSS_XI42/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI4/MM7 N_XI42/XI4/NET36_XI42/XI4/MM7_d N_XI42/XI4/NET35_XI42/XI4/MM7_g
+ N_VSS_XI42/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI4/MM8 N_XI42/XI4/NET35_XI42/XI4/MM8_d N_WL<81>_XI42/XI4/MM8_g
+ N_BLN<11>_XI42/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI4/MM5 N_XI42/XI4/NET34_XI42/XI4/MM5_d N_XI42/XI4/NET33_XI42/XI4/MM5_g
+ N_VDD_XI42/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI4/MM4 N_XI42/XI4/NET33_XI42/XI4/MM4_d N_XI42/XI4/NET34_XI42/XI4/MM4_g
+ N_VDD_XI42/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI4/MM10 N_XI42/XI4/NET35_XI42/XI4/MM10_d N_XI42/XI4/NET36_XI42/XI4/MM10_g
+ N_VDD_XI42/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI4/MM11 N_XI42/XI4/NET36_XI42/XI4/MM11_d N_XI42/XI4/NET35_XI42/XI4/MM11_g
+ N_VDD_XI42/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI5/MM2 N_XI42/XI5/NET34_XI42/XI5/MM2_d N_XI42/XI5/NET33_XI42/XI5/MM2_g
+ N_VSS_XI42/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI5/MM3 N_XI42/XI5/NET33_XI42/XI5/MM3_d N_WL<80>_XI42/XI5/MM3_g
+ N_BLN<10>_XI42/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI5/MM0 N_XI42/XI5/NET34_XI42/XI5/MM0_d N_WL<80>_XI42/XI5/MM0_g
+ N_BL<10>_XI42/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI5/MM1 N_XI42/XI5/NET33_XI42/XI5/MM1_d N_XI42/XI5/NET34_XI42/XI5/MM1_g
+ N_VSS_XI42/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI5/MM9 N_XI42/XI5/NET36_XI42/XI5/MM9_d N_WL<81>_XI42/XI5/MM9_g
+ N_BL<10>_XI42/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI5/MM6 N_XI42/XI5/NET35_XI42/XI5/MM6_d N_XI42/XI5/NET36_XI42/XI5/MM6_g
+ N_VSS_XI42/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI5/MM7 N_XI42/XI5/NET36_XI42/XI5/MM7_d N_XI42/XI5/NET35_XI42/XI5/MM7_g
+ N_VSS_XI42/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI5/MM8 N_XI42/XI5/NET35_XI42/XI5/MM8_d N_WL<81>_XI42/XI5/MM8_g
+ N_BLN<10>_XI42/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI5/MM5 N_XI42/XI5/NET34_XI42/XI5/MM5_d N_XI42/XI5/NET33_XI42/XI5/MM5_g
+ N_VDD_XI42/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI5/MM4 N_XI42/XI5/NET33_XI42/XI5/MM4_d N_XI42/XI5/NET34_XI42/XI5/MM4_g
+ N_VDD_XI42/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI5/MM10 N_XI42/XI5/NET35_XI42/XI5/MM10_d N_XI42/XI5/NET36_XI42/XI5/MM10_g
+ N_VDD_XI42/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI5/MM11 N_XI42/XI5/NET36_XI42/XI5/MM11_d N_XI42/XI5/NET35_XI42/XI5/MM11_g
+ N_VDD_XI42/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI6/MM2 N_XI42/XI6/NET34_XI42/XI6/MM2_d N_XI42/XI6/NET33_XI42/XI6/MM2_g
+ N_VSS_XI42/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM3 N_XI42/XI6/NET33_XI42/XI6/MM3_d N_WL<80>_XI42/XI6/MM3_g
+ N_BLN<9>_XI42/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM0 N_XI42/XI6/NET34_XI42/XI6/MM0_d N_WL<80>_XI42/XI6/MM0_g
+ N_BL<9>_XI42/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM1 N_XI42/XI6/NET33_XI42/XI6/MM1_d N_XI42/XI6/NET34_XI42/XI6/MM1_g
+ N_VSS_XI42/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM9 N_XI42/XI6/NET36_XI42/XI6/MM9_d N_WL<81>_XI42/XI6/MM9_g
+ N_BL<9>_XI42/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM6 N_XI42/XI6/NET35_XI42/XI6/MM6_d N_XI42/XI6/NET36_XI42/XI6/MM6_g
+ N_VSS_XI42/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM7 N_XI42/XI6/NET36_XI42/XI6/MM7_d N_XI42/XI6/NET35_XI42/XI6/MM7_g
+ N_VSS_XI42/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM8 N_XI42/XI6/NET35_XI42/XI6/MM8_d N_WL<81>_XI42/XI6/MM8_g
+ N_BLN<9>_XI42/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI6/MM5 N_XI42/XI6/NET34_XI42/XI6/MM5_d N_XI42/XI6/NET33_XI42/XI6/MM5_g
+ N_VDD_XI42/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI6/MM4 N_XI42/XI6/NET33_XI42/XI6/MM4_d N_XI42/XI6/NET34_XI42/XI6/MM4_g
+ N_VDD_XI42/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI6/MM10 N_XI42/XI6/NET35_XI42/XI6/MM10_d N_XI42/XI6/NET36_XI42/XI6/MM10_g
+ N_VDD_XI42/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI6/MM11 N_XI42/XI6/NET36_XI42/XI6/MM11_d N_XI42/XI6/NET35_XI42/XI6/MM11_g
+ N_VDD_XI42/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI7/MM2 N_XI42/XI7/NET34_XI42/XI7/MM2_d N_XI42/XI7/NET33_XI42/XI7/MM2_g
+ N_VSS_XI42/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM3 N_XI42/XI7/NET33_XI42/XI7/MM3_d N_WL<80>_XI42/XI7/MM3_g
+ N_BLN<8>_XI42/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM0 N_XI42/XI7/NET34_XI42/XI7/MM0_d N_WL<80>_XI42/XI7/MM0_g
+ N_BL<8>_XI42/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM1 N_XI42/XI7/NET33_XI42/XI7/MM1_d N_XI42/XI7/NET34_XI42/XI7/MM1_g
+ N_VSS_XI42/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM9 N_XI42/XI7/NET36_XI42/XI7/MM9_d N_WL<81>_XI42/XI7/MM9_g
+ N_BL<8>_XI42/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM6 N_XI42/XI7/NET35_XI42/XI7/MM6_d N_XI42/XI7/NET36_XI42/XI7/MM6_g
+ N_VSS_XI42/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM7 N_XI42/XI7/NET36_XI42/XI7/MM7_d N_XI42/XI7/NET35_XI42/XI7/MM7_g
+ N_VSS_XI42/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM8 N_XI42/XI7/NET35_XI42/XI7/MM8_d N_WL<81>_XI42/XI7/MM8_g
+ N_BLN<8>_XI42/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI7/MM5 N_XI42/XI7/NET34_XI42/XI7/MM5_d N_XI42/XI7/NET33_XI42/XI7/MM5_g
+ N_VDD_XI42/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI7/MM4 N_XI42/XI7/NET33_XI42/XI7/MM4_d N_XI42/XI7/NET34_XI42/XI7/MM4_g
+ N_VDD_XI42/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI7/MM10 N_XI42/XI7/NET35_XI42/XI7/MM10_d N_XI42/XI7/NET36_XI42/XI7/MM10_g
+ N_VDD_XI42/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI7/MM11 N_XI42/XI7/NET36_XI42/XI7/MM11_d N_XI42/XI7/NET35_XI42/XI7/MM11_g
+ N_VDD_XI42/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI8/MM2 N_XI42/XI8/NET34_XI42/XI8/MM2_d N_XI42/XI8/NET33_XI42/XI8/MM2_g
+ N_VSS_XI42/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM3 N_XI42/XI8/NET33_XI42/XI8/MM3_d N_WL<80>_XI42/XI8/MM3_g
+ N_BLN<7>_XI42/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM0 N_XI42/XI8/NET34_XI42/XI8/MM0_d N_WL<80>_XI42/XI8/MM0_g
+ N_BL<7>_XI42/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM1 N_XI42/XI8/NET33_XI42/XI8/MM1_d N_XI42/XI8/NET34_XI42/XI8/MM1_g
+ N_VSS_XI42/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM9 N_XI42/XI8/NET36_XI42/XI8/MM9_d N_WL<81>_XI42/XI8/MM9_g
+ N_BL<7>_XI42/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM6 N_XI42/XI8/NET35_XI42/XI8/MM6_d N_XI42/XI8/NET36_XI42/XI8/MM6_g
+ N_VSS_XI42/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM7 N_XI42/XI8/NET36_XI42/XI8/MM7_d N_XI42/XI8/NET35_XI42/XI8/MM7_g
+ N_VSS_XI42/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM8 N_XI42/XI8/NET35_XI42/XI8/MM8_d N_WL<81>_XI42/XI8/MM8_g
+ N_BLN<7>_XI42/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI8/MM5 N_XI42/XI8/NET34_XI42/XI8/MM5_d N_XI42/XI8/NET33_XI42/XI8/MM5_g
+ N_VDD_XI42/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI8/MM4 N_XI42/XI8/NET33_XI42/XI8/MM4_d N_XI42/XI8/NET34_XI42/XI8/MM4_g
+ N_VDD_XI42/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI8/MM10 N_XI42/XI8/NET35_XI42/XI8/MM10_d N_XI42/XI8/NET36_XI42/XI8/MM10_g
+ N_VDD_XI42/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI8/MM11 N_XI42/XI8/NET36_XI42/XI8/MM11_d N_XI42/XI8/NET35_XI42/XI8/MM11_g
+ N_VDD_XI42/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI9/MM2 N_XI42/XI9/NET34_XI42/XI9/MM2_d N_XI42/XI9/NET33_XI42/XI9/MM2_g
+ N_VSS_XI42/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM3 N_XI42/XI9/NET33_XI42/XI9/MM3_d N_WL<80>_XI42/XI9/MM3_g
+ N_BLN<6>_XI42/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM0 N_XI42/XI9/NET34_XI42/XI9/MM0_d N_WL<80>_XI42/XI9/MM0_g
+ N_BL<6>_XI42/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM1 N_XI42/XI9/NET33_XI42/XI9/MM1_d N_XI42/XI9/NET34_XI42/XI9/MM1_g
+ N_VSS_XI42/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM9 N_XI42/XI9/NET36_XI42/XI9/MM9_d N_WL<81>_XI42/XI9/MM9_g
+ N_BL<6>_XI42/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM6 N_XI42/XI9/NET35_XI42/XI9/MM6_d N_XI42/XI9/NET36_XI42/XI9/MM6_g
+ N_VSS_XI42/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM7 N_XI42/XI9/NET36_XI42/XI9/MM7_d N_XI42/XI9/NET35_XI42/XI9/MM7_g
+ N_VSS_XI42/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM8 N_XI42/XI9/NET35_XI42/XI9/MM8_d N_WL<81>_XI42/XI9/MM8_g
+ N_BLN<6>_XI42/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI9/MM5 N_XI42/XI9/NET34_XI42/XI9/MM5_d N_XI42/XI9/NET33_XI42/XI9/MM5_g
+ N_VDD_XI42/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI9/MM4 N_XI42/XI9/NET33_XI42/XI9/MM4_d N_XI42/XI9/NET34_XI42/XI9/MM4_g
+ N_VDD_XI42/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI9/MM10 N_XI42/XI9/NET35_XI42/XI9/MM10_d N_XI42/XI9/NET36_XI42/XI9/MM10_g
+ N_VDD_XI42/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI9/MM11 N_XI42/XI9/NET36_XI42/XI9/MM11_d N_XI42/XI9/NET35_XI42/XI9/MM11_g
+ N_VDD_XI42/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI10/MM2 N_XI42/XI10/NET34_XI42/XI10/MM2_d
+ N_XI42/XI10/NET33_XI42/XI10/MM2_g N_VSS_XI42/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI10/MM3 N_XI42/XI10/NET33_XI42/XI10/MM3_d N_WL<80>_XI42/XI10/MM3_g
+ N_BLN<5>_XI42/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI10/MM0 N_XI42/XI10/NET34_XI42/XI10/MM0_d N_WL<80>_XI42/XI10/MM0_g
+ N_BL<5>_XI42/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI10/MM1 N_XI42/XI10/NET33_XI42/XI10/MM1_d
+ N_XI42/XI10/NET34_XI42/XI10/MM1_g N_VSS_XI42/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI10/MM9 N_XI42/XI10/NET36_XI42/XI10/MM9_d N_WL<81>_XI42/XI10/MM9_g
+ N_BL<5>_XI42/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI10/MM6 N_XI42/XI10/NET35_XI42/XI10/MM6_d
+ N_XI42/XI10/NET36_XI42/XI10/MM6_g N_VSS_XI42/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI10/MM7 N_XI42/XI10/NET36_XI42/XI10/MM7_d
+ N_XI42/XI10/NET35_XI42/XI10/MM7_g N_VSS_XI42/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI10/MM8 N_XI42/XI10/NET35_XI42/XI10/MM8_d N_WL<81>_XI42/XI10/MM8_g
+ N_BLN<5>_XI42/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI10/MM5 N_XI42/XI10/NET34_XI42/XI10/MM5_d
+ N_XI42/XI10/NET33_XI42/XI10/MM5_g N_VDD_XI42/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI10/MM4 N_XI42/XI10/NET33_XI42/XI10/MM4_d
+ N_XI42/XI10/NET34_XI42/XI10/MM4_g N_VDD_XI42/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI10/MM10 N_XI42/XI10/NET35_XI42/XI10/MM10_d
+ N_XI42/XI10/NET36_XI42/XI10/MM10_g N_VDD_XI42/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI10/MM11 N_XI42/XI10/NET36_XI42/XI10/MM11_d
+ N_XI42/XI10/NET35_XI42/XI10/MM11_g N_VDD_XI42/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI11/MM2 N_XI42/XI11/NET34_XI42/XI11/MM2_d
+ N_XI42/XI11/NET33_XI42/XI11/MM2_g N_VSS_XI42/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI11/MM3 N_XI42/XI11/NET33_XI42/XI11/MM3_d N_WL<80>_XI42/XI11/MM3_g
+ N_BLN<4>_XI42/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI11/MM0 N_XI42/XI11/NET34_XI42/XI11/MM0_d N_WL<80>_XI42/XI11/MM0_g
+ N_BL<4>_XI42/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI11/MM1 N_XI42/XI11/NET33_XI42/XI11/MM1_d
+ N_XI42/XI11/NET34_XI42/XI11/MM1_g N_VSS_XI42/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI11/MM9 N_XI42/XI11/NET36_XI42/XI11/MM9_d N_WL<81>_XI42/XI11/MM9_g
+ N_BL<4>_XI42/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI11/MM6 N_XI42/XI11/NET35_XI42/XI11/MM6_d
+ N_XI42/XI11/NET36_XI42/XI11/MM6_g N_VSS_XI42/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI11/MM7 N_XI42/XI11/NET36_XI42/XI11/MM7_d
+ N_XI42/XI11/NET35_XI42/XI11/MM7_g N_VSS_XI42/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI11/MM8 N_XI42/XI11/NET35_XI42/XI11/MM8_d N_WL<81>_XI42/XI11/MM8_g
+ N_BLN<4>_XI42/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI11/MM5 N_XI42/XI11/NET34_XI42/XI11/MM5_d
+ N_XI42/XI11/NET33_XI42/XI11/MM5_g N_VDD_XI42/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI11/MM4 N_XI42/XI11/NET33_XI42/XI11/MM4_d
+ N_XI42/XI11/NET34_XI42/XI11/MM4_g N_VDD_XI42/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI11/MM10 N_XI42/XI11/NET35_XI42/XI11/MM10_d
+ N_XI42/XI11/NET36_XI42/XI11/MM10_g N_VDD_XI42/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI11/MM11 N_XI42/XI11/NET36_XI42/XI11/MM11_d
+ N_XI42/XI11/NET35_XI42/XI11/MM11_g N_VDD_XI42/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI12/MM2 N_XI42/XI12/NET34_XI42/XI12/MM2_d
+ N_XI42/XI12/NET33_XI42/XI12/MM2_g N_VSS_XI42/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI12/MM3 N_XI42/XI12/NET33_XI42/XI12/MM3_d N_WL<80>_XI42/XI12/MM3_g
+ N_BLN<3>_XI42/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI12/MM0 N_XI42/XI12/NET34_XI42/XI12/MM0_d N_WL<80>_XI42/XI12/MM0_g
+ N_BL<3>_XI42/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI12/MM1 N_XI42/XI12/NET33_XI42/XI12/MM1_d
+ N_XI42/XI12/NET34_XI42/XI12/MM1_g N_VSS_XI42/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI12/MM9 N_XI42/XI12/NET36_XI42/XI12/MM9_d N_WL<81>_XI42/XI12/MM9_g
+ N_BL<3>_XI42/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI12/MM6 N_XI42/XI12/NET35_XI42/XI12/MM6_d
+ N_XI42/XI12/NET36_XI42/XI12/MM6_g N_VSS_XI42/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI12/MM7 N_XI42/XI12/NET36_XI42/XI12/MM7_d
+ N_XI42/XI12/NET35_XI42/XI12/MM7_g N_VSS_XI42/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI12/MM8 N_XI42/XI12/NET35_XI42/XI12/MM8_d N_WL<81>_XI42/XI12/MM8_g
+ N_BLN<3>_XI42/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI12/MM5 N_XI42/XI12/NET34_XI42/XI12/MM5_d
+ N_XI42/XI12/NET33_XI42/XI12/MM5_g N_VDD_XI42/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI12/MM4 N_XI42/XI12/NET33_XI42/XI12/MM4_d
+ N_XI42/XI12/NET34_XI42/XI12/MM4_g N_VDD_XI42/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI12/MM10 N_XI42/XI12/NET35_XI42/XI12/MM10_d
+ N_XI42/XI12/NET36_XI42/XI12/MM10_g N_VDD_XI42/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI12/MM11 N_XI42/XI12/NET36_XI42/XI12/MM11_d
+ N_XI42/XI12/NET35_XI42/XI12/MM11_g N_VDD_XI42/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI13/MM2 N_XI42/XI13/NET34_XI42/XI13/MM2_d
+ N_XI42/XI13/NET33_XI42/XI13/MM2_g N_VSS_XI42/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI13/MM3 N_XI42/XI13/NET33_XI42/XI13/MM3_d N_WL<80>_XI42/XI13/MM3_g
+ N_BLN<2>_XI42/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI13/MM0 N_XI42/XI13/NET34_XI42/XI13/MM0_d N_WL<80>_XI42/XI13/MM0_g
+ N_BL<2>_XI42/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI13/MM1 N_XI42/XI13/NET33_XI42/XI13/MM1_d
+ N_XI42/XI13/NET34_XI42/XI13/MM1_g N_VSS_XI42/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI13/MM9 N_XI42/XI13/NET36_XI42/XI13/MM9_d N_WL<81>_XI42/XI13/MM9_g
+ N_BL<2>_XI42/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI13/MM6 N_XI42/XI13/NET35_XI42/XI13/MM6_d
+ N_XI42/XI13/NET36_XI42/XI13/MM6_g N_VSS_XI42/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI13/MM7 N_XI42/XI13/NET36_XI42/XI13/MM7_d
+ N_XI42/XI13/NET35_XI42/XI13/MM7_g N_VSS_XI42/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI13/MM8 N_XI42/XI13/NET35_XI42/XI13/MM8_d N_WL<81>_XI42/XI13/MM8_g
+ N_BLN<2>_XI42/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI13/MM5 N_XI42/XI13/NET34_XI42/XI13/MM5_d
+ N_XI42/XI13/NET33_XI42/XI13/MM5_g N_VDD_XI42/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI13/MM4 N_XI42/XI13/NET33_XI42/XI13/MM4_d
+ N_XI42/XI13/NET34_XI42/XI13/MM4_g N_VDD_XI42/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI13/MM10 N_XI42/XI13/NET35_XI42/XI13/MM10_d
+ N_XI42/XI13/NET36_XI42/XI13/MM10_g N_VDD_XI42/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI13/MM11 N_XI42/XI13/NET36_XI42/XI13/MM11_d
+ N_XI42/XI13/NET35_XI42/XI13/MM11_g N_VDD_XI42/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI14/MM2 N_XI42/XI14/NET34_XI42/XI14/MM2_d
+ N_XI42/XI14/NET33_XI42/XI14/MM2_g N_VSS_XI42/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI14/MM3 N_XI42/XI14/NET33_XI42/XI14/MM3_d N_WL<80>_XI42/XI14/MM3_g
+ N_BLN<1>_XI42/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI14/MM0 N_XI42/XI14/NET34_XI42/XI14/MM0_d N_WL<80>_XI42/XI14/MM0_g
+ N_BL<1>_XI42/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI14/MM1 N_XI42/XI14/NET33_XI42/XI14/MM1_d
+ N_XI42/XI14/NET34_XI42/XI14/MM1_g N_VSS_XI42/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI14/MM9 N_XI42/XI14/NET36_XI42/XI14/MM9_d N_WL<81>_XI42/XI14/MM9_g
+ N_BL<1>_XI42/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI14/MM6 N_XI42/XI14/NET35_XI42/XI14/MM6_d
+ N_XI42/XI14/NET36_XI42/XI14/MM6_g N_VSS_XI42/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI14/MM7 N_XI42/XI14/NET36_XI42/XI14/MM7_d
+ N_XI42/XI14/NET35_XI42/XI14/MM7_g N_VSS_XI42/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI14/MM8 N_XI42/XI14/NET35_XI42/XI14/MM8_d N_WL<81>_XI42/XI14/MM8_g
+ N_BLN<1>_XI42/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI14/MM5 N_XI42/XI14/NET34_XI42/XI14/MM5_d
+ N_XI42/XI14/NET33_XI42/XI14/MM5_g N_VDD_XI42/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI14/MM4 N_XI42/XI14/NET33_XI42/XI14/MM4_d
+ N_XI42/XI14/NET34_XI42/XI14/MM4_g N_VDD_XI42/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI14/MM10 N_XI42/XI14/NET35_XI42/XI14/MM10_d
+ N_XI42/XI14/NET36_XI42/XI14/MM10_g N_VDD_XI42/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI14/MM11 N_XI42/XI14/NET36_XI42/XI14/MM11_d
+ N_XI42/XI14/NET35_XI42/XI14/MM11_g N_VDD_XI42/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI15/MM2 N_XI42/XI15/NET34_XI42/XI15/MM2_d
+ N_XI42/XI15/NET33_XI42/XI15/MM2_g N_VSS_XI42/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI15/MM3 N_XI42/XI15/NET33_XI42/XI15/MM3_d N_WL<80>_XI42/XI15/MM3_g
+ N_BLN<0>_XI42/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI15/MM0 N_XI42/XI15/NET34_XI42/XI15/MM0_d N_WL<80>_XI42/XI15/MM0_g
+ N_BL<0>_XI42/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI15/MM1 N_XI42/XI15/NET33_XI42/XI15/MM1_d
+ N_XI42/XI15/NET34_XI42/XI15/MM1_g N_VSS_XI42/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI15/MM9 N_XI42/XI15/NET36_XI42/XI15/MM9_d N_WL<81>_XI42/XI15/MM9_g
+ N_BL<0>_XI42/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI15/MM6 N_XI42/XI15/NET35_XI42/XI15/MM6_d
+ N_XI42/XI15/NET36_XI42/XI15/MM6_g N_VSS_XI42/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI15/MM7 N_XI42/XI15/NET36_XI42/XI15/MM7_d
+ N_XI42/XI15/NET35_XI42/XI15/MM7_g N_VSS_XI42/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI42/XI15/MM8 N_XI42/XI15/NET35_XI42/XI15/MM8_d N_WL<81>_XI42/XI15/MM8_g
+ N_BLN<0>_XI42/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI42/XI15/MM5 N_XI42/XI15/NET34_XI42/XI15/MM5_d
+ N_XI42/XI15/NET33_XI42/XI15/MM5_g N_VDD_XI42/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI15/MM4 N_XI42/XI15/NET33_XI42/XI15/MM4_d
+ N_XI42/XI15/NET34_XI42/XI15/MM4_g N_VDD_XI42/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI15/MM10 N_XI42/XI15/NET35_XI42/XI15/MM10_d
+ N_XI42/XI15/NET36_XI42/XI15/MM10_g N_VDD_XI42/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI42/XI15/MM11 N_XI42/XI15/NET36_XI42/XI15/MM11_d
+ N_XI42/XI15/NET35_XI42/XI15/MM11_g N_VDD_XI42/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI0/MM2 N_XI43/XI0/NET34_XI43/XI0/MM2_d N_XI43/XI0/NET33_XI43/XI0/MM2_g
+ N_VSS_XI43/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI0/MM3 N_XI43/XI0/NET33_XI43/XI0/MM3_d N_WL<82>_XI43/XI0/MM3_g
+ N_BLN<15>_XI43/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI0/MM0 N_XI43/XI0/NET34_XI43/XI0/MM0_d N_WL<82>_XI43/XI0/MM0_g
+ N_BL<15>_XI43/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI0/MM1 N_XI43/XI0/NET33_XI43/XI0/MM1_d N_XI43/XI0/NET34_XI43/XI0/MM1_g
+ N_VSS_XI43/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI0/MM9 N_XI43/XI0/NET36_XI43/XI0/MM9_d N_WL<83>_XI43/XI0/MM9_g
+ N_BL<15>_XI43/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI0/MM6 N_XI43/XI0/NET35_XI43/XI0/MM6_d N_XI43/XI0/NET36_XI43/XI0/MM6_g
+ N_VSS_XI43/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI0/MM7 N_XI43/XI0/NET36_XI43/XI0/MM7_d N_XI43/XI0/NET35_XI43/XI0/MM7_g
+ N_VSS_XI43/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI0/MM8 N_XI43/XI0/NET35_XI43/XI0/MM8_d N_WL<83>_XI43/XI0/MM8_g
+ N_BLN<15>_XI43/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI0/MM5 N_XI43/XI0/NET34_XI43/XI0/MM5_d N_XI43/XI0/NET33_XI43/XI0/MM5_g
+ N_VDD_XI43/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI0/MM4 N_XI43/XI0/NET33_XI43/XI0/MM4_d N_XI43/XI0/NET34_XI43/XI0/MM4_g
+ N_VDD_XI43/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI0/MM10 N_XI43/XI0/NET35_XI43/XI0/MM10_d N_XI43/XI0/NET36_XI43/XI0/MM10_g
+ N_VDD_XI43/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI0/MM11 N_XI43/XI0/NET36_XI43/XI0/MM11_d N_XI43/XI0/NET35_XI43/XI0/MM11_g
+ N_VDD_XI43/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI1/MM2 N_XI43/XI1/NET34_XI43/XI1/MM2_d N_XI43/XI1/NET33_XI43/XI1/MM2_g
+ N_VSS_XI43/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI1/MM3 N_XI43/XI1/NET33_XI43/XI1/MM3_d N_WL<82>_XI43/XI1/MM3_g
+ N_BLN<14>_XI43/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI1/MM0 N_XI43/XI1/NET34_XI43/XI1/MM0_d N_WL<82>_XI43/XI1/MM0_g
+ N_BL<14>_XI43/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI1/MM1 N_XI43/XI1/NET33_XI43/XI1/MM1_d N_XI43/XI1/NET34_XI43/XI1/MM1_g
+ N_VSS_XI43/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI1/MM9 N_XI43/XI1/NET36_XI43/XI1/MM9_d N_WL<83>_XI43/XI1/MM9_g
+ N_BL<14>_XI43/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI1/MM6 N_XI43/XI1/NET35_XI43/XI1/MM6_d N_XI43/XI1/NET36_XI43/XI1/MM6_g
+ N_VSS_XI43/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI1/MM7 N_XI43/XI1/NET36_XI43/XI1/MM7_d N_XI43/XI1/NET35_XI43/XI1/MM7_g
+ N_VSS_XI43/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI1/MM8 N_XI43/XI1/NET35_XI43/XI1/MM8_d N_WL<83>_XI43/XI1/MM8_g
+ N_BLN<14>_XI43/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI1/MM5 N_XI43/XI1/NET34_XI43/XI1/MM5_d N_XI43/XI1/NET33_XI43/XI1/MM5_g
+ N_VDD_XI43/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI1/MM4 N_XI43/XI1/NET33_XI43/XI1/MM4_d N_XI43/XI1/NET34_XI43/XI1/MM4_g
+ N_VDD_XI43/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI1/MM10 N_XI43/XI1/NET35_XI43/XI1/MM10_d N_XI43/XI1/NET36_XI43/XI1/MM10_g
+ N_VDD_XI43/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI1/MM11 N_XI43/XI1/NET36_XI43/XI1/MM11_d N_XI43/XI1/NET35_XI43/XI1/MM11_g
+ N_VDD_XI43/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI2/MM2 N_XI43/XI2/NET34_XI43/XI2/MM2_d N_XI43/XI2/NET33_XI43/XI2/MM2_g
+ N_VSS_XI43/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI2/MM3 N_XI43/XI2/NET33_XI43/XI2/MM3_d N_WL<82>_XI43/XI2/MM3_g
+ N_BLN<13>_XI43/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI2/MM0 N_XI43/XI2/NET34_XI43/XI2/MM0_d N_WL<82>_XI43/XI2/MM0_g
+ N_BL<13>_XI43/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI2/MM1 N_XI43/XI2/NET33_XI43/XI2/MM1_d N_XI43/XI2/NET34_XI43/XI2/MM1_g
+ N_VSS_XI43/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI2/MM9 N_XI43/XI2/NET36_XI43/XI2/MM9_d N_WL<83>_XI43/XI2/MM9_g
+ N_BL<13>_XI43/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI2/MM6 N_XI43/XI2/NET35_XI43/XI2/MM6_d N_XI43/XI2/NET36_XI43/XI2/MM6_g
+ N_VSS_XI43/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI2/MM7 N_XI43/XI2/NET36_XI43/XI2/MM7_d N_XI43/XI2/NET35_XI43/XI2/MM7_g
+ N_VSS_XI43/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI2/MM8 N_XI43/XI2/NET35_XI43/XI2/MM8_d N_WL<83>_XI43/XI2/MM8_g
+ N_BLN<13>_XI43/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI2/MM5 N_XI43/XI2/NET34_XI43/XI2/MM5_d N_XI43/XI2/NET33_XI43/XI2/MM5_g
+ N_VDD_XI43/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI2/MM4 N_XI43/XI2/NET33_XI43/XI2/MM4_d N_XI43/XI2/NET34_XI43/XI2/MM4_g
+ N_VDD_XI43/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI2/MM10 N_XI43/XI2/NET35_XI43/XI2/MM10_d N_XI43/XI2/NET36_XI43/XI2/MM10_g
+ N_VDD_XI43/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI2/MM11 N_XI43/XI2/NET36_XI43/XI2/MM11_d N_XI43/XI2/NET35_XI43/XI2/MM11_g
+ N_VDD_XI43/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI3/MM2 N_XI43/XI3/NET34_XI43/XI3/MM2_d N_XI43/XI3/NET33_XI43/XI3/MM2_g
+ N_VSS_XI43/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI3/MM3 N_XI43/XI3/NET33_XI43/XI3/MM3_d N_WL<82>_XI43/XI3/MM3_g
+ N_BLN<12>_XI43/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI3/MM0 N_XI43/XI3/NET34_XI43/XI3/MM0_d N_WL<82>_XI43/XI3/MM0_g
+ N_BL<12>_XI43/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI3/MM1 N_XI43/XI3/NET33_XI43/XI3/MM1_d N_XI43/XI3/NET34_XI43/XI3/MM1_g
+ N_VSS_XI43/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI3/MM9 N_XI43/XI3/NET36_XI43/XI3/MM9_d N_WL<83>_XI43/XI3/MM9_g
+ N_BL<12>_XI43/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI3/MM6 N_XI43/XI3/NET35_XI43/XI3/MM6_d N_XI43/XI3/NET36_XI43/XI3/MM6_g
+ N_VSS_XI43/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI3/MM7 N_XI43/XI3/NET36_XI43/XI3/MM7_d N_XI43/XI3/NET35_XI43/XI3/MM7_g
+ N_VSS_XI43/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI3/MM8 N_XI43/XI3/NET35_XI43/XI3/MM8_d N_WL<83>_XI43/XI3/MM8_g
+ N_BLN<12>_XI43/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI3/MM5 N_XI43/XI3/NET34_XI43/XI3/MM5_d N_XI43/XI3/NET33_XI43/XI3/MM5_g
+ N_VDD_XI43/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI3/MM4 N_XI43/XI3/NET33_XI43/XI3/MM4_d N_XI43/XI3/NET34_XI43/XI3/MM4_g
+ N_VDD_XI43/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI3/MM10 N_XI43/XI3/NET35_XI43/XI3/MM10_d N_XI43/XI3/NET36_XI43/XI3/MM10_g
+ N_VDD_XI43/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI3/MM11 N_XI43/XI3/NET36_XI43/XI3/MM11_d N_XI43/XI3/NET35_XI43/XI3/MM11_g
+ N_VDD_XI43/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI4/MM2 N_XI43/XI4/NET34_XI43/XI4/MM2_d N_XI43/XI4/NET33_XI43/XI4/MM2_g
+ N_VSS_XI43/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI4/MM3 N_XI43/XI4/NET33_XI43/XI4/MM3_d N_WL<82>_XI43/XI4/MM3_g
+ N_BLN<11>_XI43/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI4/MM0 N_XI43/XI4/NET34_XI43/XI4/MM0_d N_WL<82>_XI43/XI4/MM0_g
+ N_BL<11>_XI43/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI4/MM1 N_XI43/XI4/NET33_XI43/XI4/MM1_d N_XI43/XI4/NET34_XI43/XI4/MM1_g
+ N_VSS_XI43/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI4/MM9 N_XI43/XI4/NET36_XI43/XI4/MM9_d N_WL<83>_XI43/XI4/MM9_g
+ N_BL<11>_XI43/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI4/MM6 N_XI43/XI4/NET35_XI43/XI4/MM6_d N_XI43/XI4/NET36_XI43/XI4/MM6_g
+ N_VSS_XI43/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI4/MM7 N_XI43/XI4/NET36_XI43/XI4/MM7_d N_XI43/XI4/NET35_XI43/XI4/MM7_g
+ N_VSS_XI43/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI4/MM8 N_XI43/XI4/NET35_XI43/XI4/MM8_d N_WL<83>_XI43/XI4/MM8_g
+ N_BLN<11>_XI43/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI4/MM5 N_XI43/XI4/NET34_XI43/XI4/MM5_d N_XI43/XI4/NET33_XI43/XI4/MM5_g
+ N_VDD_XI43/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI4/MM4 N_XI43/XI4/NET33_XI43/XI4/MM4_d N_XI43/XI4/NET34_XI43/XI4/MM4_g
+ N_VDD_XI43/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI4/MM10 N_XI43/XI4/NET35_XI43/XI4/MM10_d N_XI43/XI4/NET36_XI43/XI4/MM10_g
+ N_VDD_XI43/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI4/MM11 N_XI43/XI4/NET36_XI43/XI4/MM11_d N_XI43/XI4/NET35_XI43/XI4/MM11_g
+ N_VDD_XI43/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI5/MM2 N_XI43/XI5/NET34_XI43/XI5/MM2_d N_XI43/XI5/NET33_XI43/XI5/MM2_g
+ N_VSS_XI43/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI5/MM3 N_XI43/XI5/NET33_XI43/XI5/MM3_d N_WL<82>_XI43/XI5/MM3_g
+ N_BLN<10>_XI43/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI5/MM0 N_XI43/XI5/NET34_XI43/XI5/MM0_d N_WL<82>_XI43/XI5/MM0_g
+ N_BL<10>_XI43/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI5/MM1 N_XI43/XI5/NET33_XI43/XI5/MM1_d N_XI43/XI5/NET34_XI43/XI5/MM1_g
+ N_VSS_XI43/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI5/MM9 N_XI43/XI5/NET36_XI43/XI5/MM9_d N_WL<83>_XI43/XI5/MM9_g
+ N_BL<10>_XI43/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI5/MM6 N_XI43/XI5/NET35_XI43/XI5/MM6_d N_XI43/XI5/NET36_XI43/XI5/MM6_g
+ N_VSS_XI43/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI5/MM7 N_XI43/XI5/NET36_XI43/XI5/MM7_d N_XI43/XI5/NET35_XI43/XI5/MM7_g
+ N_VSS_XI43/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI5/MM8 N_XI43/XI5/NET35_XI43/XI5/MM8_d N_WL<83>_XI43/XI5/MM8_g
+ N_BLN<10>_XI43/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI5/MM5 N_XI43/XI5/NET34_XI43/XI5/MM5_d N_XI43/XI5/NET33_XI43/XI5/MM5_g
+ N_VDD_XI43/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI5/MM4 N_XI43/XI5/NET33_XI43/XI5/MM4_d N_XI43/XI5/NET34_XI43/XI5/MM4_g
+ N_VDD_XI43/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI5/MM10 N_XI43/XI5/NET35_XI43/XI5/MM10_d N_XI43/XI5/NET36_XI43/XI5/MM10_g
+ N_VDD_XI43/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI5/MM11 N_XI43/XI5/NET36_XI43/XI5/MM11_d N_XI43/XI5/NET35_XI43/XI5/MM11_g
+ N_VDD_XI43/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI6/MM2 N_XI43/XI6/NET34_XI43/XI6/MM2_d N_XI43/XI6/NET33_XI43/XI6/MM2_g
+ N_VSS_XI43/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM3 N_XI43/XI6/NET33_XI43/XI6/MM3_d N_WL<82>_XI43/XI6/MM3_g
+ N_BLN<9>_XI43/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM0 N_XI43/XI6/NET34_XI43/XI6/MM0_d N_WL<82>_XI43/XI6/MM0_g
+ N_BL<9>_XI43/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM1 N_XI43/XI6/NET33_XI43/XI6/MM1_d N_XI43/XI6/NET34_XI43/XI6/MM1_g
+ N_VSS_XI43/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM9 N_XI43/XI6/NET36_XI43/XI6/MM9_d N_WL<83>_XI43/XI6/MM9_g
+ N_BL<9>_XI43/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM6 N_XI43/XI6/NET35_XI43/XI6/MM6_d N_XI43/XI6/NET36_XI43/XI6/MM6_g
+ N_VSS_XI43/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM7 N_XI43/XI6/NET36_XI43/XI6/MM7_d N_XI43/XI6/NET35_XI43/XI6/MM7_g
+ N_VSS_XI43/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM8 N_XI43/XI6/NET35_XI43/XI6/MM8_d N_WL<83>_XI43/XI6/MM8_g
+ N_BLN<9>_XI43/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI6/MM5 N_XI43/XI6/NET34_XI43/XI6/MM5_d N_XI43/XI6/NET33_XI43/XI6/MM5_g
+ N_VDD_XI43/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI6/MM4 N_XI43/XI6/NET33_XI43/XI6/MM4_d N_XI43/XI6/NET34_XI43/XI6/MM4_g
+ N_VDD_XI43/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI6/MM10 N_XI43/XI6/NET35_XI43/XI6/MM10_d N_XI43/XI6/NET36_XI43/XI6/MM10_g
+ N_VDD_XI43/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI6/MM11 N_XI43/XI6/NET36_XI43/XI6/MM11_d N_XI43/XI6/NET35_XI43/XI6/MM11_g
+ N_VDD_XI43/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI7/MM2 N_XI43/XI7/NET34_XI43/XI7/MM2_d N_XI43/XI7/NET33_XI43/XI7/MM2_g
+ N_VSS_XI43/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM3 N_XI43/XI7/NET33_XI43/XI7/MM3_d N_WL<82>_XI43/XI7/MM3_g
+ N_BLN<8>_XI43/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM0 N_XI43/XI7/NET34_XI43/XI7/MM0_d N_WL<82>_XI43/XI7/MM0_g
+ N_BL<8>_XI43/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM1 N_XI43/XI7/NET33_XI43/XI7/MM1_d N_XI43/XI7/NET34_XI43/XI7/MM1_g
+ N_VSS_XI43/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM9 N_XI43/XI7/NET36_XI43/XI7/MM9_d N_WL<83>_XI43/XI7/MM9_g
+ N_BL<8>_XI43/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM6 N_XI43/XI7/NET35_XI43/XI7/MM6_d N_XI43/XI7/NET36_XI43/XI7/MM6_g
+ N_VSS_XI43/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM7 N_XI43/XI7/NET36_XI43/XI7/MM7_d N_XI43/XI7/NET35_XI43/XI7/MM7_g
+ N_VSS_XI43/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM8 N_XI43/XI7/NET35_XI43/XI7/MM8_d N_WL<83>_XI43/XI7/MM8_g
+ N_BLN<8>_XI43/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI7/MM5 N_XI43/XI7/NET34_XI43/XI7/MM5_d N_XI43/XI7/NET33_XI43/XI7/MM5_g
+ N_VDD_XI43/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI7/MM4 N_XI43/XI7/NET33_XI43/XI7/MM4_d N_XI43/XI7/NET34_XI43/XI7/MM4_g
+ N_VDD_XI43/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI7/MM10 N_XI43/XI7/NET35_XI43/XI7/MM10_d N_XI43/XI7/NET36_XI43/XI7/MM10_g
+ N_VDD_XI43/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI7/MM11 N_XI43/XI7/NET36_XI43/XI7/MM11_d N_XI43/XI7/NET35_XI43/XI7/MM11_g
+ N_VDD_XI43/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI8/MM2 N_XI43/XI8/NET34_XI43/XI8/MM2_d N_XI43/XI8/NET33_XI43/XI8/MM2_g
+ N_VSS_XI43/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM3 N_XI43/XI8/NET33_XI43/XI8/MM3_d N_WL<82>_XI43/XI8/MM3_g
+ N_BLN<7>_XI43/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM0 N_XI43/XI8/NET34_XI43/XI8/MM0_d N_WL<82>_XI43/XI8/MM0_g
+ N_BL<7>_XI43/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM1 N_XI43/XI8/NET33_XI43/XI8/MM1_d N_XI43/XI8/NET34_XI43/XI8/MM1_g
+ N_VSS_XI43/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM9 N_XI43/XI8/NET36_XI43/XI8/MM9_d N_WL<83>_XI43/XI8/MM9_g
+ N_BL<7>_XI43/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM6 N_XI43/XI8/NET35_XI43/XI8/MM6_d N_XI43/XI8/NET36_XI43/XI8/MM6_g
+ N_VSS_XI43/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM7 N_XI43/XI8/NET36_XI43/XI8/MM7_d N_XI43/XI8/NET35_XI43/XI8/MM7_g
+ N_VSS_XI43/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM8 N_XI43/XI8/NET35_XI43/XI8/MM8_d N_WL<83>_XI43/XI8/MM8_g
+ N_BLN<7>_XI43/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI8/MM5 N_XI43/XI8/NET34_XI43/XI8/MM5_d N_XI43/XI8/NET33_XI43/XI8/MM5_g
+ N_VDD_XI43/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI8/MM4 N_XI43/XI8/NET33_XI43/XI8/MM4_d N_XI43/XI8/NET34_XI43/XI8/MM4_g
+ N_VDD_XI43/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI8/MM10 N_XI43/XI8/NET35_XI43/XI8/MM10_d N_XI43/XI8/NET36_XI43/XI8/MM10_g
+ N_VDD_XI43/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI8/MM11 N_XI43/XI8/NET36_XI43/XI8/MM11_d N_XI43/XI8/NET35_XI43/XI8/MM11_g
+ N_VDD_XI43/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI9/MM2 N_XI43/XI9/NET34_XI43/XI9/MM2_d N_XI43/XI9/NET33_XI43/XI9/MM2_g
+ N_VSS_XI43/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM3 N_XI43/XI9/NET33_XI43/XI9/MM3_d N_WL<82>_XI43/XI9/MM3_g
+ N_BLN<6>_XI43/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM0 N_XI43/XI9/NET34_XI43/XI9/MM0_d N_WL<82>_XI43/XI9/MM0_g
+ N_BL<6>_XI43/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM1 N_XI43/XI9/NET33_XI43/XI9/MM1_d N_XI43/XI9/NET34_XI43/XI9/MM1_g
+ N_VSS_XI43/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM9 N_XI43/XI9/NET36_XI43/XI9/MM9_d N_WL<83>_XI43/XI9/MM9_g
+ N_BL<6>_XI43/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM6 N_XI43/XI9/NET35_XI43/XI9/MM6_d N_XI43/XI9/NET36_XI43/XI9/MM6_g
+ N_VSS_XI43/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM7 N_XI43/XI9/NET36_XI43/XI9/MM7_d N_XI43/XI9/NET35_XI43/XI9/MM7_g
+ N_VSS_XI43/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM8 N_XI43/XI9/NET35_XI43/XI9/MM8_d N_WL<83>_XI43/XI9/MM8_g
+ N_BLN<6>_XI43/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI9/MM5 N_XI43/XI9/NET34_XI43/XI9/MM5_d N_XI43/XI9/NET33_XI43/XI9/MM5_g
+ N_VDD_XI43/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI9/MM4 N_XI43/XI9/NET33_XI43/XI9/MM4_d N_XI43/XI9/NET34_XI43/XI9/MM4_g
+ N_VDD_XI43/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI9/MM10 N_XI43/XI9/NET35_XI43/XI9/MM10_d N_XI43/XI9/NET36_XI43/XI9/MM10_g
+ N_VDD_XI43/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI9/MM11 N_XI43/XI9/NET36_XI43/XI9/MM11_d N_XI43/XI9/NET35_XI43/XI9/MM11_g
+ N_VDD_XI43/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI10/MM2 N_XI43/XI10/NET34_XI43/XI10/MM2_d
+ N_XI43/XI10/NET33_XI43/XI10/MM2_g N_VSS_XI43/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI10/MM3 N_XI43/XI10/NET33_XI43/XI10/MM3_d N_WL<82>_XI43/XI10/MM3_g
+ N_BLN<5>_XI43/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI10/MM0 N_XI43/XI10/NET34_XI43/XI10/MM0_d N_WL<82>_XI43/XI10/MM0_g
+ N_BL<5>_XI43/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI10/MM1 N_XI43/XI10/NET33_XI43/XI10/MM1_d
+ N_XI43/XI10/NET34_XI43/XI10/MM1_g N_VSS_XI43/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI10/MM9 N_XI43/XI10/NET36_XI43/XI10/MM9_d N_WL<83>_XI43/XI10/MM9_g
+ N_BL<5>_XI43/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI10/MM6 N_XI43/XI10/NET35_XI43/XI10/MM6_d
+ N_XI43/XI10/NET36_XI43/XI10/MM6_g N_VSS_XI43/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI10/MM7 N_XI43/XI10/NET36_XI43/XI10/MM7_d
+ N_XI43/XI10/NET35_XI43/XI10/MM7_g N_VSS_XI43/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI10/MM8 N_XI43/XI10/NET35_XI43/XI10/MM8_d N_WL<83>_XI43/XI10/MM8_g
+ N_BLN<5>_XI43/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI10/MM5 N_XI43/XI10/NET34_XI43/XI10/MM5_d
+ N_XI43/XI10/NET33_XI43/XI10/MM5_g N_VDD_XI43/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI10/MM4 N_XI43/XI10/NET33_XI43/XI10/MM4_d
+ N_XI43/XI10/NET34_XI43/XI10/MM4_g N_VDD_XI43/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI10/MM10 N_XI43/XI10/NET35_XI43/XI10/MM10_d
+ N_XI43/XI10/NET36_XI43/XI10/MM10_g N_VDD_XI43/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI10/MM11 N_XI43/XI10/NET36_XI43/XI10/MM11_d
+ N_XI43/XI10/NET35_XI43/XI10/MM11_g N_VDD_XI43/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI11/MM2 N_XI43/XI11/NET34_XI43/XI11/MM2_d
+ N_XI43/XI11/NET33_XI43/XI11/MM2_g N_VSS_XI43/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI11/MM3 N_XI43/XI11/NET33_XI43/XI11/MM3_d N_WL<82>_XI43/XI11/MM3_g
+ N_BLN<4>_XI43/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI11/MM0 N_XI43/XI11/NET34_XI43/XI11/MM0_d N_WL<82>_XI43/XI11/MM0_g
+ N_BL<4>_XI43/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI11/MM1 N_XI43/XI11/NET33_XI43/XI11/MM1_d
+ N_XI43/XI11/NET34_XI43/XI11/MM1_g N_VSS_XI43/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI11/MM9 N_XI43/XI11/NET36_XI43/XI11/MM9_d N_WL<83>_XI43/XI11/MM9_g
+ N_BL<4>_XI43/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI11/MM6 N_XI43/XI11/NET35_XI43/XI11/MM6_d
+ N_XI43/XI11/NET36_XI43/XI11/MM6_g N_VSS_XI43/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI11/MM7 N_XI43/XI11/NET36_XI43/XI11/MM7_d
+ N_XI43/XI11/NET35_XI43/XI11/MM7_g N_VSS_XI43/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI11/MM8 N_XI43/XI11/NET35_XI43/XI11/MM8_d N_WL<83>_XI43/XI11/MM8_g
+ N_BLN<4>_XI43/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI11/MM5 N_XI43/XI11/NET34_XI43/XI11/MM5_d
+ N_XI43/XI11/NET33_XI43/XI11/MM5_g N_VDD_XI43/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI11/MM4 N_XI43/XI11/NET33_XI43/XI11/MM4_d
+ N_XI43/XI11/NET34_XI43/XI11/MM4_g N_VDD_XI43/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI11/MM10 N_XI43/XI11/NET35_XI43/XI11/MM10_d
+ N_XI43/XI11/NET36_XI43/XI11/MM10_g N_VDD_XI43/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI11/MM11 N_XI43/XI11/NET36_XI43/XI11/MM11_d
+ N_XI43/XI11/NET35_XI43/XI11/MM11_g N_VDD_XI43/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI12/MM2 N_XI43/XI12/NET34_XI43/XI12/MM2_d
+ N_XI43/XI12/NET33_XI43/XI12/MM2_g N_VSS_XI43/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI12/MM3 N_XI43/XI12/NET33_XI43/XI12/MM3_d N_WL<82>_XI43/XI12/MM3_g
+ N_BLN<3>_XI43/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI12/MM0 N_XI43/XI12/NET34_XI43/XI12/MM0_d N_WL<82>_XI43/XI12/MM0_g
+ N_BL<3>_XI43/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI12/MM1 N_XI43/XI12/NET33_XI43/XI12/MM1_d
+ N_XI43/XI12/NET34_XI43/XI12/MM1_g N_VSS_XI43/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI12/MM9 N_XI43/XI12/NET36_XI43/XI12/MM9_d N_WL<83>_XI43/XI12/MM9_g
+ N_BL<3>_XI43/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI12/MM6 N_XI43/XI12/NET35_XI43/XI12/MM6_d
+ N_XI43/XI12/NET36_XI43/XI12/MM6_g N_VSS_XI43/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI12/MM7 N_XI43/XI12/NET36_XI43/XI12/MM7_d
+ N_XI43/XI12/NET35_XI43/XI12/MM7_g N_VSS_XI43/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI12/MM8 N_XI43/XI12/NET35_XI43/XI12/MM8_d N_WL<83>_XI43/XI12/MM8_g
+ N_BLN<3>_XI43/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI12/MM5 N_XI43/XI12/NET34_XI43/XI12/MM5_d
+ N_XI43/XI12/NET33_XI43/XI12/MM5_g N_VDD_XI43/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI12/MM4 N_XI43/XI12/NET33_XI43/XI12/MM4_d
+ N_XI43/XI12/NET34_XI43/XI12/MM4_g N_VDD_XI43/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI12/MM10 N_XI43/XI12/NET35_XI43/XI12/MM10_d
+ N_XI43/XI12/NET36_XI43/XI12/MM10_g N_VDD_XI43/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI12/MM11 N_XI43/XI12/NET36_XI43/XI12/MM11_d
+ N_XI43/XI12/NET35_XI43/XI12/MM11_g N_VDD_XI43/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI13/MM2 N_XI43/XI13/NET34_XI43/XI13/MM2_d
+ N_XI43/XI13/NET33_XI43/XI13/MM2_g N_VSS_XI43/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI13/MM3 N_XI43/XI13/NET33_XI43/XI13/MM3_d N_WL<82>_XI43/XI13/MM3_g
+ N_BLN<2>_XI43/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI13/MM0 N_XI43/XI13/NET34_XI43/XI13/MM0_d N_WL<82>_XI43/XI13/MM0_g
+ N_BL<2>_XI43/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI13/MM1 N_XI43/XI13/NET33_XI43/XI13/MM1_d
+ N_XI43/XI13/NET34_XI43/XI13/MM1_g N_VSS_XI43/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI13/MM9 N_XI43/XI13/NET36_XI43/XI13/MM9_d N_WL<83>_XI43/XI13/MM9_g
+ N_BL<2>_XI43/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI13/MM6 N_XI43/XI13/NET35_XI43/XI13/MM6_d
+ N_XI43/XI13/NET36_XI43/XI13/MM6_g N_VSS_XI43/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI13/MM7 N_XI43/XI13/NET36_XI43/XI13/MM7_d
+ N_XI43/XI13/NET35_XI43/XI13/MM7_g N_VSS_XI43/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI13/MM8 N_XI43/XI13/NET35_XI43/XI13/MM8_d N_WL<83>_XI43/XI13/MM8_g
+ N_BLN<2>_XI43/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI13/MM5 N_XI43/XI13/NET34_XI43/XI13/MM5_d
+ N_XI43/XI13/NET33_XI43/XI13/MM5_g N_VDD_XI43/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI13/MM4 N_XI43/XI13/NET33_XI43/XI13/MM4_d
+ N_XI43/XI13/NET34_XI43/XI13/MM4_g N_VDD_XI43/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI13/MM10 N_XI43/XI13/NET35_XI43/XI13/MM10_d
+ N_XI43/XI13/NET36_XI43/XI13/MM10_g N_VDD_XI43/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI13/MM11 N_XI43/XI13/NET36_XI43/XI13/MM11_d
+ N_XI43/XI13/NET35_XI43/XI13/MM11_g N_VDD_XI43/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI14/MM2 N_XI43/XI14/NET34_XI43/XI14/MM2_d
+ N_XI43/XI14/NET33_XI43/XI14/MM2_g N_VSS_XI43/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI14/MM3 N_XI43/XI14/NET33_XI43/XI14/MM3_d N_WL<82>_XI43/XI14/MM3_g
+ N_BLN<1>_XI43/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI14/MM0 N_XI43/XI14/NET34_XI43/XI14/MM0_d N_WL<82>_XI43/XI14/MM0_g
+ N_BL<1>_XI43/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI14/MM1 N_XI43/XI14/NET33_XI43/XI14/MM1_d
+ N_XI43/XI14/NET34_XI43/XI14/MM1_g N_VSS_XI43/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI14/MM9 N_XI43/XI14/NET36_XI43/XI14/MM9_d N_WL<83>_XI43/XI14/MM9_g
+ N_BL<1>_XI43/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI14/MM6 N_XI43/XI14/NET35_XI43/XI14/MM6_d
+ N_XI43/XI14/NET36_XI43/XI14/MM6_g N_VSS_XI43/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI14/MM7 N_XI43/XI14/NET36_XI43/XI14/MM7_d
+ N_XI43/XI14/NET35_XI43/XI14/MM7_g N_VSS_XI43/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI14/MM8 N_XI43/XI14/NET35_XI43/XI14/MM8_d N_WL<83>_XI43/XI14/MM8_g
+ N_BLN<1>_XI43/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI14/MM5 N_XI43/XI14/NET34_XI43/XI14/MM5_d
+ N_XI43/XI14/NET33_XI43/XI14/MM5_g N_VDD_XI43/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI14/MM4 N_XI43/XI14/NET33_XI43/XI14/MM4_d
+ N_XI43/XI14/NET34_XI43/XI14/MM4_g N_VDD_XI43/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI14/MM10 N_XI43/XI14/NET35_XI43/XI14/MM10_d
+ N_XI43/XI14/NET36_XI43/XI14/MM10_g N_VDD_XI43/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI14/MM11 N_XI43/XI14/NET36_XI43/XI14/MM11_d
+ N_XI43/XI14/NET35_XI43/XI14/MM11_g N_VDD_XI43/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI15/MM2 N_XI43/XI15/NET34_XI43/XI15/MM2_d
+ N_XI43/XI15/NET33_XI43/XI15/MM2_g N_VSS_XI43/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI15/MM3 N_XI43/XI15/NET33_XI43/XI15/MM3_d N_WL<82>_XI43/XI15/MM3_g
+ N_BLN<0>_XI43/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI15/MM0 N_XI43/XI15/NET34_XI43/XI15/MM0_d N_WL<82>_XI43/XI15/MM0_g
+ N_BL<0>_XI43/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI15/MM1 N_XI43/XI15/NET33_XI43/XI15/MM1_d
+ N_XI43/XI15/NET34_XI43/XI15/MM1_g N_VSS_XI43/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI15/MM9 N_XI43/XI15/NET36_XI43/XI15/MM9_d N_WL<83>_XI43/XI15/MM9_g
+ N_BL<0>_XI43/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI15/MM6 N_XI43/XI15/NET35_XI43/XI15/MM6_d
+ N_XI43/XI15/NET36_XI43/XI15/MM6_g N_VSS_XI43/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI15/MM7 N_XI43/XI15/NET36_XI43/XI15/MM7_d
+ N_XI43/XI15/NET35_XI43/XI15/MM7_g N_VSS_XI43/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI43/XI15/MM8 N_XI43/XI15/NET35_XI43/XI15/MM8_d N_WL<83>_XI43/XI15/MM8_g
+ N_BLN<0>_XI43/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI43/XI15/MM5 N_XI43/XI15/NET34_XI43/XI15/MM5_d
+ N_XI43/XI15/NET33_XI43/XI15/MM5_g N_VDD_XI43/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI15/MM4 N_XI43/XI15/NET33_XI43/XI15/MM4_d
+ N_XI43/XI15/NET34_XI43/XI15/MM4_g N_VDD_XI43/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI15/MM10 N_XI43/XI15/NET35_XI43/XI15/MM10_d
+ N_XI43/XI15/NET36_XI43/XI15/MM10_g N_VDD_XI43/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI43/XI15/MM11 N_XI43/XI15/NET36_XI43/XI15/MM11_d
+ N_XI43/XI15/NET35_XI43/XI15/MM11_g N_VDD_XI43/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI0/MM2 N_XI44/XI0/NET34_XI44/XI0/MM2_d N_XI44/XI0/NET33_XI44/XI0/MM2_g
+ N_VSS_XI44/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI0/MM3 N_XI44/XI0/NET33_XI44/XI0/MM3_d N_WL<84>_XI44/XI0/MM3_g
+ N_BLN<15>_XI44/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI0/MM0 N_XI44/XI0/NET34_XI44/XI0/MM0_d N_WL<84>_XI44/XI0/MM0_g
+ N_BL<15>_XI44/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI0/MM1 N_XI44/XI0/NET33_XI44/XI0/MM1_d N_XI44/XI0/NET34_XI44/XI0/MM1_g
+ N_VSS_XI44/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI0/MM9 N_XI44/XI0/NET36_XI44/XI0/MM9_d N_WL<85>_XI44/XI0/MM9_g
+ N_BL<15>_XI44/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI0/MM6 N_XI44/XI0/NET35_XI44/XI0/MM6_d N_XI44/XI0/NET36_XI44/XI0/MM6_g
+ N_VSS_XI44/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI0/MM7 N_XI44/XI0/NET36_XI44/XI0/MM7_d N_XI44/XI0/NET35_XI44/XI0/MM7_g
+ N_VSS_XI44/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI0/MM8 N_XI44/XI0/NET35_XI44/XI0/MM8_d N_WL<85>_XI44/XI0/MM8_g
+ N_BLN<15>_XI44/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI0/MM5 N_XI44/XI0/NET34_XI44/XI0/MM5_d N_XI44/XI0/NET33_XI44/XI0/MM5_g
+ N_VDD_XI44/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI0/MM4 N_XI44/XI0/NET33_XI44/XI0/MM4_d N_XI44/XI0/NET34_XI44/XI0/MM4_g
+ N_VDD_XI44/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI0/MM10 N_XI44/XI0/NET35_XI44/XI0/MM10_d N_XI44/XI0/NET36_XI44/XI0/MM10_g
+ N_VDD_XI44/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI0/MM11 N_XI44/XI0/NET36_XI44/XI0/MM11_d N_XI44/XI0/NET35_XI44/XI0/MM11_g
+ N_VDD_XI44/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI1/MM2 N_XI44/XI1/NET34_XI44/XI1/MM2_d N_XI44/XI1/NET33_XI44/XI1/MM2_g
+ N_VSS_XI44/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI1/MM3 N_XI44/XI1/NET33_XI44/XI1/MM3_d N_WL<84>_XI44/XI1/MM3_g
+ N_BLN<14>_XI44/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI1/MM0 N_XI44/XI1/NET34_XI44/XI1/MM0_d N_WL<84>_XI44/XI1/MM0_g
+ N_BL<14>_XI44/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI1/MM1 N_XI44/XI1/NET33_XI44/XI1/MM1_d N_XI44/XI1/NET34_XI44/XI1/MM1_g
+ N_VSS_XI44/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI1/MM9 N_XI44/XI1/NET36_XI44/XI1/MM9_d N_WL<85>_XI44/XI1/MM9_g
+ N_BL<14>_XI44/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI1/MM6 N_XI44/XI1/NET35_XI44/XI1/MM6_d N_XI44/XI1/NET36_XI44/XI1/MM6_g
+ N_VSS_XI44/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI1/MM7 N_XI44/XI1/NET36_XI44/XI1/MM7_d N_XI44/XI1/NET35_XI44/XI1/MM7_g
+ N_VSS_XI44/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI1/MM8 N_XI44/XI1/NET35_XI44/XI1/MM8_d N_WL<85>_XI44/XI1/MM8_g
+ N_BLN<14>_XI44/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI1/MM5 N_XI44/XI1/NET34_XI44/XI1/MM5_d N_XI44/XI1/NET33_XI44/XI1/MM5_g
+ N_VDD_XI44/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI1/MM4 N_XI44/XI1/NET33_XI44/XI1/MM4_d N_XI44/XI1/NET34_XI44/XI1/MM4_g
+ N_VDD_XI44/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI1/MM10 N_XI44/XI1/NET35_XI44/XI1/MM10_d N_XI44/XI1/NET36_XI44/XI1/MM10_g
+ N_VDD_XI44/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI1/MM11 N_XI44/XI1/NET36_XI44/XI1/MM11_d N_XI44/XI1/NET35_XI44/XI1/MM11_g
+ N_VDD_XI44/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI2/MM2 N_XI44/XI2/NET34_XI44/XI2/MM2_d N_XI44/XI2/NET33_XI44/XI2/MM2_g
+ N_VSS_XI44/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI2/MM3 N_XI44/XI2/NET33_XI44/XI2/MM3_d N_WL<84>_XI44/XI2/MM3_g
+ N_BLN<13>_XI44/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI2/MM0 N_XI44/XI2/NET34_XI44/XI2/MM0_d N_WL<84>_XI44/XI2/MM0_g
+ N_BL<13>_XI44/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI2/MM1 N_XI44/XI2/NET33_XI44/XI2/MM1_d N_XI44/XI2/NET34_XI44/XI2/MM1_g
+ N_VSS_XI44/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI2/MM9 N_XI44/XI2/NET36_XI44/XI2/MM9_d N_WL<85>_XI44/XI2/MM9_g
+ N_BL<13>_XI44/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI2/MM6 N_XI44/XI2/NET35_XI44/XI2/MM6_d N_XI44/XI2/NET36_XI44/XI2/MM6_g
+ N_VSS_XI44/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI2/MM7 N_XI44/XI2/NET36_XI44/XI2/MM7_d N_XI44/XI2/NET35_XI44/XI2/MM7_g
+ N_VSS_XI44/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI2/MM8 N_XI44/XI2/NET35_XI44/XI2/MM8_d N_WL<85>_XI44/XI2/MM8_g
+ N_BLN<13>_XI44/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI2/MM5 N_XI44/XI2/NET34_XI44/XI2/MM5_d N_XI44/XI2/NET33_XI44/XI2/MM5_g
+ N_VDD_XI44/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI2/MM4 N_XI44/XI2/NET33_XI44/XI2/MM4_d N_XI44/XI2/NET34_XI44/XI2/MM4_g
+ N_VDD_XI44/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI2/MM10 N_XI44/XI2/NET35_XI44/XI2/MM10_d N_XI44/XI2/NET36_XI44/XI2/MM10_g
+ N_VDD_XI44/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI2/MM11 N_XI44/XI2/NET36_XI44/XI2/MM11_d N_XI44/XI2/NET35_XI44/XI2/MM11_g
+ N_VDD_XI44/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI3/MM2 N_XI44/XI3/NET34_XI44/XI3/MM2_d N_XI44/XI3/NET33_XI44/XI3/MM2_g
+ N_VSS_XI44/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI3/MM3 N_XI44/XI3/NET33_XI44/XI3/MM3_d N_WL<84>_XI44/XI3/MM3_g
+ N_BLN<12>_XI44/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI3/MM0 N_XI44/XI3/NET34_XI44/XI3/MM0_d N_WL<84>_XI44/XI3/MM0_g
+ N_BL<12>_XI44/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI3/MM1 N_XI44/XI3/NET33_XI44/XI3/MM1_d N_XI44/XI3/NET34_XI44/XI3/MM1_g
+ N_VSS_XI44/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI3/MM9 N_XI44/XI3/NET36_XI44/XI3/MM9_d N_WL<85>_XI44/XI3/MM9_g
+ N_BL<12>_XI44/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI3/MM6 N_XI44/XI3/NET35_XI44/XI3/MM6_d N_XI44/XI3/NET36_XI44/XI3/MM6_g
+ N_VSS_XI44/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI3/MM7 N_XI44/XI3/NET36_XI44/XI3/MM7_d N_XI44/XI3/NET35_XI44/XI3/MM7_g
+ N_VSS_XI44/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI3/MM8 N_XI44/XI3/NET35_XI44/XI3/MM8_d N_WL<85>_XI44/XI3/MM8_g
+ N_BLN<12>_XI44/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI3/MM5 N_XI44/XI3/NET34_XI44/XI3/MM5_d N_XI44/XI3/NET33_XI44/XI3/MM5_g
+ N_VDD_XI44/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI3/MM4 N_XI44/XI3/NET33_XI44/XI3/MM4_d N_XI44/XI3/NET34_XI44/XI3/MM4_g
+ N_VDD_XI44/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI3/MM10 N_XI44/XI3/NET35_XI44/XI3/MM10_d N_XI44/XI3/NET36_XI44/XI3/MM10_g
+ N_VDD_XI44/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI3/MM11 N_XI44/XI3/NET36_XI44/XI3/MM11_d N_XI44/XI3/NET35_XI44/XI3/MM11_g
+ N_VDD_XI44/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI4/MM2 N_XI44/XI4/NET34_XI44/XI4/MM2_d N_XI44/XI4/NET33_XI44/XI4/MM2_g
+ N_VSS_XI44/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI4/MM3 N_XI44/XI4/NET33_XI44/XI4/MM3_d N_WL<84>_XI44/XI4/MM3_g
+ N_BLN<11>_XI44/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI4/MM0 N_XI44/XI4/NET34_XI44/XI4/MM0_d N_WL<84>_XI44/XI4/MM0_g
+ N_BL<11>_XI44/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI4/MM1 N_XI44/XI4/NET33_XI44/XI4/MM1_d N_XI44/XI4/NET34_XI44/XI4/MM1_g
+ N_VSS_XI44/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI4/MM9 N_XI44/XI4/NET36_XI44/XI4/MM9_d N_WL<85>_XI44/XI4/MM9_g
+ N_BL<11>_XI44/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI4/MM6 N_XI44/XI4/NET35_XI44/XI4/MM6_d N_XI44/XI4/NET36_XI44/XI4/MM6_g
+ N_VSS_XI44/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI4/MM7 N_XI44/XI4/NET36_XI44/XI4/MM7_d N_XI44/XI4/NET35_XI44/XI4/MM7_g
+ N_VSS_XI44/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI4/MM8 N_XI44/XI4/NET35_XI44/XI4/MM8_d N_WL<85>_XI44/XI4/MM8_g
+ N_BLN<11>_XI44/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI4/MM5 N_XI44/XI4/NET34_XI44/XI4/MM5_d N_XI44/XI4/NET33_XI44/XI4/MM5_g
+ N_VDD_XI44/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI4/MM4 N_XI44/XI4/NET33_XI44/XI4/MM4_d N_XI44/XI4/NET34_XI44/XI4/MM4_g
+ N_VDD_XI44/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI4/MM10 N_XI44/XI4/NET35_XI44/XI4/MM10_d N_XI44/XI4/NET36_XI44/XI4/MM10_g
+ N_VDD_XI44/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI4/MM11 N_XI44/XI4/NET36_XI44/XI4/MM11_d N_XI44/XI4/NET35_XI44/XI4/MM11_g
+ N_VDD_XI44/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI5/MM2 N_XI44/XI5/NET34_XI44/XI5/MM2_d N_XI44/XI5/NET33_XI44/XI5/MM2_g
+ N_VSS_XI44/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI5/MM3 N_XI44/XI5/NET33_XI44/XI5/MM3_d N_WL<84>_XI44/XI5/MM3_g
+ N_BLN<10>_XI44/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI5/MM0 N_XI44/XI5/NET34_XI44/XI5/MM0_d N_WL<84>_XI44/XI5/MM0_g
+ N_BL<10>_XI44/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI5/MM1 N_XI44/XI5/NET33_XI44/XI5/MM1_d N_XI44/XI5/NET34_XI44/XI5/MM1_g
+ N_VSS_XI44/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI5/MM9 N_XI44/XI5/NET36_XI44/XI5/MM9_d N_WL<85>_XI44/XI5/MM9_g
+ N_BL<10>_XI44/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI5/MM6 N_XI44/XI5/NET35_XI44/XI5/MM6_d N_XI44/XI5/NET36_XI44/XI5/MM6_g
+ N_VSS_XI44/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI5/MM7 N_XI44/XI5/NET36_XI44/XI5/MM7_d N_XI44/XI5/NET35_XI44/XI5/MM7_g
+ N_VSS_XI44/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI5/MM8 N_XI44/XI5/NET35_XI44/XI5/MM8_d N_WL<85>_XI44/XI5/MM8_g
+ N_BLN<10>_XI44/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI5/MM5 N_XI44/XI5/NET34_XI44/XI5/MM5_d N_XI44/XI5/NET33_XI44/XI5/MM5_g
+ N_VDD_XI44/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI5/MM4 N_XI44/XI5/NET33_XI44/XI5/MM4_d N_XI44/XI5/NET34_XI44/XI5/MM4_g
+ N_VDD_XI44/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI5/MM10 N_XI44/XI5/NET35_XI44/XI5/MM10_d N_XI44/XI5/NET36_XI44/XI5/MM10_g
+ N_VDD_XI44/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI5/MM11 N_XI44/XI5/NET36_XI44/XI5/MM11_d N_XI44/XI5/NET35_XI44/XI5/MM11_g
+ N_VDD_XI44/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI6/MM2 N_XI44/XI6/NET34_XI44/XI6/MM2_d N_XI44/XI6/NET33_XI44/XI6/MM2_g
+ N_VSS_XI44/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM3 N_XI44/XI6/NET33_XI44/XI6/MM3_d N_WL<84>_XI44/XI6/MM3_g
+ N_BLN<9>_XI44/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM0 N_XI44/XI6/NET34_XI44/XI6/MM0_d N_WL<84>_XI44/XI6/MM0_g
+ N_BL<9>_XI44/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM1 N_XI44/XI6/NET33_XI44/XI6/MM1_d N_XI44/XI6/NET34_XI44/XI6/MM1_g
+ N_VSS_XI44/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM9 N_XI44/XI6/NET36_XI44/XI6/MM9_d N_WL<85>_XI44/XI6/MM9_g
+ N_BL<9>_XI44/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM6 N_XI44/XI6/NET35_XI44/XI6/MM6_d N_XI44/XI6/NET36_XI44/XI6/MM6_g
+ N_VSS_XI44/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM7 N_XI44/XI6/NET36_XI44/XI6/MM7_d N_XI44/XI6/NET35_XI44/XI6/MM7_g
+ N_VSS_XI44/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM8 N_XI44/XI6/NET35_XI44/XI6/MM8_d N_WL<85>_XI44/XI6/MM8_g
+ N_BLN<9>_XI44/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI6/MM5 N_XI44/XI6/NET34_XI44/XI6/MM5_d N_XI44/XI6/NET33_XI44/XI6/MM5_g
+ N_VDD_XI44/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI6/MM4 N_XI44/XI6/NET33_XI44/XI6/MM4_d N_XI44/XI6/NET34_XI44/XI6/MM4_g
+ N_VDD_XI44/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI6/MM10 N_XI44/XI6/NET35_XI44/XI6/MM10_d N_XI44/XI6/NET36_XI44/XI6/MM10_g
+ N_VDD_XI44/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI6/MM11 N_XI44/XI6/NET36_XI44/XI6/MM11_d N_XI44/XI6/NET35_XI44/XI6/MM11_g
+ N_VDD_XI44/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI7/MM2 N_XI44/XI7/NET34_XI44/XI7/MM2_d N_XI44/XI7/NET33_XI44/XI7/MM2_g
+ N_VSS_XI44/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM3 N_XI44/XI7/NET33_XI44/XI7/MM3_d N_WL<84>_XI44/XI7/MM3_g
+ N_BLN<8>_XI44/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM0 N_XI44/XI7/NET34_XI44/XI7/MM0_d N_WL<84>_XI44/XI7/MM0_g
+ N_BL<8>_XI44/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM1 N_XI44/XI7/NET33_XI44/XI7/MM1_d N_XI44/XI7/NET34_XI44/XI7/MM1_g
+ N_VSS_XI44/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM9 N_XI44/XI7/NET36_XI44/XI7/MM9_d N_WL<85>_XI44/XI7/MM9_g
+ N_BL<8>_XI44/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM6 N_XI44/XI7/NET35_XI44/XI7/MM6_d N_XI44/XI7/NET36_XI44/XI7/MM6_g
+ N_VSS_XI44/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM7 N_XI44/XI7/NET36_XI44/XI7/MM7_d N_XI44/XI7/NET35_XI44/XI7/MM7_g
+ N_VSS_XI44/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM8 N_XI44/XI7/NET35_XI44/XI7/MM8_d N_WL<85>_XI44/XI7/MM8_g
+ N_BLN<8>_XI44/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI7/MM5 N_XI44/XI7/NET34_XI44/XI7/MM5_d N_XI44/XI7/NET33_XI44/XI7/MM5_g
+ N_VDD_XI44/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI7/MM4 N_XI44/XI7/NET33_XI44/XI7/MM4_d N_XI44/XI7/NET34_XI44/XI7/MM4_g
+ N_VDD_XI44/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI7/MM10 N_XI44/XI7/NET35_XI44/XI7/MM10_d N_XI44/XI7/NET36_XI44/XI7/MM10_g
+ N_VDD_XI44/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI7/MM11 N_XI44/XI7/NET36_XI44/XI7/MM11_d N_XI44/XI7/NET35_XI44/XI7/MM11_g
+ N_VDD_XI44/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI8/MM2 N_XI44/XI8/NET34_XI44/XI8/MM2_d N_XI44/XI8/NET33_XI44/XI8/MM2_g
+ N_VSS_XI44/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM3 N_XI44/XI8/NET33_XI44/XI8/MM3_d N_WL<84>_XI44/XI8/MM3_g
+ N_BLN<7>_XI44/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM0 N_XI44/XI8/NET34_XI44/XI8/MM0_d N_WL<84>_XI44/XI8/MM0_g
+ N_BL<7>_XI44/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM1 N_XI44/XI8/NET33_XI44/XI8/MM1_d N_XI44/XI8/NET34_XI44/XI8/MM1_g
+ N_VSS_XI44/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM9 N_XI44/XI8/NET36_XI44/XI8/MM9_d N_WL<85>_XI44/XI8/MM9_g
+ N_BL<7>_XI44/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM6 N_XI44/XI8/NET35_XI44/XI8/MM6_d N_XI44/XI8/NET36_XI44/XI8/MM6_g
+ N_VSS_XI44/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM7 N_XI44/XI8/NET36_XI44/XI8/MM7_d N_XI44/XI8/NET35_XI44/XI8/MM7_g
+ N_VSS_XI44/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM8 N_XI44/XI8/NET35_XI44/XI8/MM8_d N_WL<85>_XI44/XI8/MM8_g
+ N_BLN<7>_XI44/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI8/MM5 N_XI44/XI8/NET34_XI44/XI8/MM5_d N_XI44/XI8/NET33_XI44/XI8/MM5_g
+ N_VDD_XI44/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI8/MM4 N_XI44/XI8/NET33_XI44/XI8/MM4_d N_XI44/XI8/NET34_XI44/XI8/MM4_g
+ N_VDD_XI44/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI8/MM10 N_XI44/XI8/NET35_XI44/XI8/MM10_d N_XI44/XI8/NET36_XI44/XI8/MM10_g
+ N_VDD_XI44/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI8/MM11 N_XI44/XI8/NET36_XI44/XI8/MM11_d N_XI44/XI8/NET35_XI44/XI8/MM11_g
+ N_VDD_XI44/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI9/MM2 N_XI44/XI9/NET34_XI44/XI9/MM2_d N_XI44/XI9/NET33_XI44/XI9/MM2_g
+ N_VSS_XI44/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM3 N_XI44/XI9/NET33_XI44/XI9/MM3_d N_WL<84>_XI44/XI9/MM3_g
+ N_BLN<6>_XI44/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM0 N_XI44/XI9/NET34_XI44/XI9/MM0_d N_WL<84>_XI44/XI9/MM0_g
+ N_BL<6>_XI44/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM1 N_XI44/XI9/NET33_XI44/XI9/MM1_d N_XI44/XI9/NET34_XI44/XI9/MM1_g
+ N_VSS_XI44/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM9 N_XI44/XI9/NET36_XI44/XI9/MM9_d N_WL<85>_XI44/XI9/MM9_g
+ N_BL<6>_XI44/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM6 N_XI44/XI9/NET35_XI44/XI9/MM6_d N_XI44/XI9/NET36_XI44/XI9/MM6_g
+ N_VSS_XI44/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM7 N_XI44/XI9/NET36_XI44/XI9/MM7_d N_XI44/XI9/NET35_XI44/XI9/MM7_g
+ N_VSS_XI44/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM8 N_XI44/XI9/NET35_XI44/XI9/MM8_d N_WL<85>_XI44/XI9/MM8_g
+ N_BLN<6>_XI44/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI9/MM5 N_XI44/XI9/NET34_XI44/XI9/MM5_d N_XI44/XI9/NET33_XI44/XI9/MM5_g
+ N_VDD_XI44/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI9/MM4 N_XI44/XI9/NET33_XI44/XI9/MM4_d N_XI44/XI9/NET34_XI44/XI9/MM4_g
+ N_VDD_XI44/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI9/MM10 N_XI44/XI9/NET35_XI44/XI9/MM10_d N_XI44/XI9/NET36_XI44/XI9/MM10_g
+ N_VDD_XI44/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI9/MM11 N_XI44/XI9/NET36_XI44/XI9/MM11_d N_XI44/XI9/NET35_XI44/XI9/MM11_g
+ N_VDD_XI44/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI10/MM2 N_XI44/XI10/NET34_XI44/XI10/MM2_d
+ N_XI44/XI10/NET33_XI44/XI10/MM2_g N_VSS_XI44/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI10/MM3 N_XI44/XI10/NET33_XI44/XI10/MM3_d N_WL<84>_XI44/XI10/MM3_g
+ N_BLN<5>_XI44/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI10/MM0 N_XI44/XI10/NET34_XI44/XI10/MM0_d N_WL<84>_XI44/XI10/MM0_g
+ N_BL<5>_XI44/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI10/MM1 N_XI44/XI10/NET33_XI44/XI10/MM1_d
+ N_XI44/XI10/NET34_XI44/XI10/MM1_g N_VSS_XI44/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI10/MM9 N_XI44/XI10/NET36_XI44/XI10/MM9_d N_WL<85>_XI44/XI10/MM9_g
+ N_BL<5>_XI44/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI10/MM6 N_XI44/XI10/NET35_XI44/XI10/MM6_d
+ N_XI44/XI10/NET36_XI44/XI10/MM6_g N_VSS_XI44/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI10/MM7 N_XI44/XI10/NET36_XI44/XI10/MM7_d
+ N_XI44/XI10/NET35_XI44/XI10/MM7_g N_VSS_XI44/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI10/MM8 N_XI44/XI10/NET35_XI44/XI10/MM8_d N_WL<85>_XI44/XI10/MM8_g
+ N_BLN<5>_XI44/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI10/MM5 N_XI44/XI10/NET34_XI44/XI10/MM5_d
+ N_XI44/XI10/NET33_XI44/XI10/MM5_g N_VDD_XI44/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI10/MM4 N_XI44/XI10/NET33_XI44/XI10/MM4_d
+ N_XI44/XI10/NET34_XI44/XI10/MM4_g N_VDD_XI44/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI10/MM10 N_XI44/XI10/NET35_XI44/XI10/MM10_d
+ N_XI44/XI10/NET36_XI44/XI10/MM10_g N_VDD_XI44/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI10/MM11 N_XI44/XI10/NET36_XI44/XI10/MM11_d
+ N_XI44/XI10/NET35_XI44/XI10/MM11_g N_VDD_XI44/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI11/MM2 N_XI44/XI11/NET34_XI44/XI11/MM2_d
+ N_XI44/XI11/NET33_XI44/XI11/MM2_g N_VSS_XI44/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI11/MM3 N_XI44/XI11/NET33_XI44/XI11/MM3_d N_WL<84>_XI44/XI11/MM3_g
+ N_BLN<4>_XI44/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI11/MM0 N_XI44/XI11/NET34_XI44/XI11/MM0_d N_WL<84>_XI44/XI11/MM0_g
+ N_BL<4>_XI44/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI11/MM1 N_XI44/XI11/NET33_XI44/XI11/MM1_d
+ N_XI44/XI11/NET34_XI44/XI11/MM1_g N_VSS_XI44/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI11/MM9 N_XI44/XI11/NET36_XI44/XI11/MM9_d N_WL<85>_XI44/XI11/MM9_g
+ N_BL<4>_XI44/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI11/MM6 N_XI44/XI11/NET35_XI44/XI11/MM6_d
+ N_XI44/XI11/NET36_XI44/XI11/MM6_g N_VSS_XI44/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI11/MM7 N_XI44/XI11/NET36_XI44/XI11/MM7_d
+ N_XI44/XI11/NET35_XI44/XI11/MM7_g N_VSS_XI44/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI11/MM8 N_XI44/XI11/NET35_XI44/XI11/MM8_d N_WL<85>_XI44/XI11/MM8_g
+ N_BLN<4>_XI44/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI11/MM5 N_XI44/XI11/NET34_XI44/XI11/MM5_d
+ N_XI44/XI11/NET33_XI44/XI11/MM5_g N_VDD_XI44/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI11/MM4 N_XI44/XI11/NET33_XI44/XI11/MM4_d
+ N_XI44/XI11/NET34_XI44/XI11/MM4_g N_VDD_XI44/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI11/MM10 N_XI44/XI11/NET35_XI44/XI11/MM10_d
+ N_XI44/XI11/NET36_XI44/XI11/MM10_g N_VDD_XI44/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI11/MM11 N_XI44/XI11/NET36_XI44/XI11/MM11_d
+ N_XI44/XI11/NET35_XI44/XI11/MM11_g N_VDD_XI44/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI12/MM2 N_XI44/XI12/NET34_XI44/XI12/MM2_d
+ N_XI44/XI12/NET33_XI44/XI12/MM2_g N_VSS_XI44/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI12/MM3 N_XI44/XI12/NET33_XI44/XI12/MM3_d N_WL<84>_XI44/XI12/MM3_g
+ N_BLN<3>_XI44/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI12/MM0 N_XI44/XI12/NET34_XI44/XI12/MM0_d N_WL<84>_XI44/XI12/MM0_g
+ N_BL<3>_XI44/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI12/MM1 N_XI44/XI12/NET33_XI44/XI12/MM1_d
+ N_XI44/XI12/NET34_XI44/XI12/MM1_g N_VSS_XI44/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI12/MM9 N_XI44/XI12/NET36_XI44/XI12/MM9_d N_WL<85>_XI44/XI12/MM9_g
+ N_BL<3>_XI44/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI12/MM6 N_XI44/XI12/NET35_XI44/XI12/MM6_d
+ N_XI44/XI12/NET36_XI44/XI12/MM6_g N_VSS_XI44/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI12/MM7 N_XI44/XI12/NET36_XI44/XI12/MM7_d
+ N_XI44/XI12/NET35_XI44/XI12/MM7_g N_VSS_XI44/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI12/MM8 N_XI44/XI12/NET35_XI44/XI12/MM8_d N_WL<85>_XI44/XI12/MM8_g
+ N_BLN<3>_XI44/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI12/MM5 N_XI44/XI12/NET34_XI44/XI12/MM5_d
+ N_XI44/XI12/NET33_XI44/XI12/MM5_g N_VDD_XI44/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI12/MM4 N_XI44/XI12/NET33_XI44/XI12/MM4_d
+ N_XI44/XI12/NET34_XI44/XI12/MM4_g N_VDD_XI44/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI12/MM10 N_XI44/XI12/NET35_XI44/XI12/MM10_d
+ N_XI44/XI12/NET36_XI44/XI12/MM10_g N_VDD_XI44/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI12/MM11 N_XI44/XI12/NET36_XI44/XI12/MM11_d
+ N_XI44/XI12/NET35_XI44/XI12/MM11_g N_VDD_XI44/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI13/MM2 N_XI44/XI13/NET34_XI44/XI13/MM2_d
+ N_XI44/XI13/NET33_XI44/XI13/MM2_g N_VSS_XI44/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI13/MM3 N_XI44/XI13/NET33_XI44/XI13/MM3_d N_WL<84>_XI44/XI13/MM3_g
+ N_BLN<2>_XI44/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI13/MM0 N_XI44/XI13/NET34_XI44/XI13/MM0_d N_WL<84>_XI44/XI13/MM0_g
+ N_BL<2>_XI44/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI13/MM1 N_XI44/XI13/NET33_XI44/XI13/MM1_d
+ N_XI44/XI13/NET34_XI44/XI13/MM1_g N_VSS_XI44/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI13/MM9 N_XI44/XI13/NET36_XI44/XI13/MM9_d N_WL<85>_XI44/XI13/MM9_g
+ N_BL<2>_XI44/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI13/MM6 N_XI44/XI13/NET35_XI44/XI13/MM6_d
+ N_XI44/XI13/NET36_XI44/XI13/MM6_g N_VSS_XI44/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI13/MM7 N_XI44/XI13/NET36_XI44/XI13/MM7_d
+ N_XI44/XI13/NET35_XI44/XI13/MM7_g N_VSS_XI44/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI13/MM8 N_XI44/XI13/NET35_XI44/XI13/MM8_d N_WL<85>_XI44/XI13/MM8_g
+ N_BLN<2>_XI44/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI13/MM5 N_XI44/XI13/NET34_XI44/XI13/MM5_d
+ N_XI44/XI13/NET33_XI44/XI13/MM5_g N_VDD_XI44/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI13/MM4 N_XI44/XI13/NET33_XI44/XI13/MM4_d
+ N_XI44/XI13/NET34_XI44/XI13/MM4_g N_VDD_XI44/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI13/MM10 N_XI44/XI13/NET35_XI44/XI13/MM10_d
+ N_XI44/XI13/NET36_XI44/XI13/MM10_g N_VDD_XI44/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI13/MM11 N_XI44/XI13/NET36_XI44/XI13/MM11_d
+ N_XI44/XI13/NET35_XI44/XI13/MM11_g N_VDD_XI44/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI14/MM2 N_XI44/XI14/NET34_XI44/XI14/MM2_d
+ N_XI44/XI14/NET33_XI44/XI14/MM2_g N_VSS_XI44/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI14/MM3 N_XI44/XI14/NET33_XI44/XI14/MM3_d N_WL<84>_XI44/XI14/MM3_g
+ N_BLN<1>_XI44/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI14/MM0 N_XI44/XI14/NET34_XI44/XI14/MM0_d N_WL<84>_XI44/XI14/MM0_g
+ N_BL<1>_XI44/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI14/MM1 N_XI44/XI14/NET33_XI44/XI14/MM1_d
+ N_XI44/XI14/NET34_XI44/XI14/MM1_g N_VSS_XI44/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI14/MM9 N_XI44/XI14/NET36_XI44/XI14/MM9_d N_WL<85>_XI44/XI14/MM9_g
+ N_BL<1>_XI44/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI14/MM6 N_XI44/XI14/NET35_XI44/XI14/MM6_d
+ N_XI44/XI14/NET36_XI44/XI14/MM6_g N_VSS_XI44/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI14/MM7 N_XI44/XI14/NET36_XI44/XI14/MM7_d
+ N_XI44/XI14/NET35_XI44/XI14/MM7_g N_VSS_XI44/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI14/MM8 N_XI44/XI14/NET35_XI44/XI14/MM8_d N_WL<85>_XI44/XI14/MM8_g
+ N_BLN<1>_XI44/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI14/MM5 N_XI44/XI14/NET34_XI44/XI14/MM5_d
+ N_XI44/XI14/NET33_XI44/XI14/MM5_g N_VDD_XI44/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI14/MM4 N_XI44/XI14/NET33_XI44/XI14/MM4_d
+ N_XI44/XI14/NET34_XI44/XI14/MM4_g N_VDD_XI44/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI14/MM10 N_XI44/XI14/NET35_XI44/XI14/MM10_d
+ N_XI44/XI14/NET36_XI44/XI14/MM10_g N_VDD_XI44/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI14/MM11 N_XI44/XI14/NET36_XI44/XI14/MM11_d
+ N_XI44/XI14/NET35_XI44/XI14/MM11_g N_VDD_XI44/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI15/MM2 N_XI44/XI15/NET34_XI44/XI15/MM2_d
+ N_XI44/XI15/NET33_XI44/XI15/MM2_g N_VSS_XI44/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI15/MM3 N_XI44/XI15/NET33_XI44/XI15/MM3_d N_WL<84>_XI44/XI15/MM3_g
+ N_BLN<0>_XI44/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI15/MM0 N_XI44/XI15/NET34_XI44/XI15/MM0_d N_WL<84>_XI44/XI15/MM0_g
+ N_BL<0>_XI44/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI15/MM1 N_XI44/XI15/NET33_XI44/XI15/MM1_d
+ N_XI44/XI15/NET34_XI44/XI15/MM1_g N_VSS_XI44/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI15/MM9 N_XI44/XI15/NET36_XI44/XI15/MM9_d N_WL<85>_XI44/XI15/MM9_g
+ N_BL<0>_XI44/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI15/MM6 N_XI44/XI15/NET35_XI44/XI15/MM6_d
+ N_XI44/XI15/NET36_XI44/XI15/MM6_g N_VSS_XI44/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI15/MM7 N_XI44/XI15/NET36_XI44/XI15/MM7_d
+ N_XI44/XI15/NET35_XI44/XI15/MM7_g N_VSS_XI44/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI44/XI15/MM8 N_XI44/XI15/NET35_XI44/XI15/MM8_d N_WL<85>_XI44/XI15/MM8_g
+ N_BLN<0>_XI44/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI44/XI15/MM5 N_XI44/XI15/NET34_XI44/XI15/MM5_d
+ N_XI44/XI15/NET33_XI44/XI15/MM5_g N_VDD_XI44/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI15/MM4 N_XI44/XI15/NET33_XI44/XI15/MM4_d
+ N_XI44/XI15/NET34_XI44/XI15/MM4_g N_VDD_XI44/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI15/MM10 N_XI44/XI15/NET35_XI44/XI15/MM10_d
+ N_XI44/XI15/NET36_XI44/XI15/MM10_g N_VDD_XI44/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI44/XI15/MM11 N_XI44/XI15/NET36_XI44/XI15/MM11_d
+ N_XI44/XI15/NET35_XI44/XI15/MM11_g N_VDD_XI44/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI0/MM2 N_XI45/XI0/NET34_XI45/XI0/MM2_d N_XI45/XI0/NET33_XI45/XI0/MM2_g
+ N_VSS_XI45/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI0/MM3 N_XI45/XI0/NET33_XI45/XI0/MM3_d N_WL<86>_XI45/XI0/MM3_g
+ N_BLN<15>_XI45/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI0/MM0 N_XI45/XI0/NET34_XI45/XI0/MM0_d N_WL<86>_XI45/XI0/MM0_g
+ N_BL<15>_XI45/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI0/MM1 N_XI45/XI0/NET33_XI45/XI0/MM1_d N_XI45/XI0/NET34_XI45/XI0/MM1_g
+ N_VSS_XI45/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI0/MM9 N_XI45/XI0/NET36_XI45/XI0/MM9_d N_WL<87>_XI45/XI0/MM9_g
+ N_BL<15>_XI45/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI0/MM6 N_XI45/XI0/NET35_XI45/XI0/MM6_d N_XI45/XI0/NET36_XI45/XI0/MM6_g
+ N_VSS_XI45/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI0/MM7 N_XI45/XI0/NET36_XI45/XI0/MM7_d N_XI45/XI0/NET35_XI45/XI0/MM7_g
+ N_VSS_XI45/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI0/MM8 N_XI45/XI0/NET35_XI45/XI0/MM8_d N_WL<87>_XI45/XI0/MM8_g
+ N_BLN<15>_XI45/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI0/MM5 N_XI45/XI0/NET34_XI45/XI0/MM5_d N_XI45/XI0/NET33_XI45/XI0/MM5_g
+ N_VDD_XI45/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI0/MM4 N_XI45/XI0/NET33_XI45/XI0/MM4_d N_XI45/XI0/NET34_XI45/XI0/MM4_g
+ N_VDD_XI45/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI0/MM10 N_XI45/XI0/NET35_XI45/XI0/MM10_d N_XI45/XI0/NET36_XI45/XI0/MM10_g
+ N_VDD_XI45/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI0/MM11 N_XI45/XI0/NET36_XI45/XI0/MM11_d N_XI45/XI0/NET35_XI45/XI0/MM11_g
+ N_VDD_XI45/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI1/MM2 N_XI45/XI1/NET34_XI45/XI1/MM2_d N_XI45/XI1/NET33_XI45/XI1/MM2_g
+ N_VSS_XI45/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI1/MM3 N_XI45/XI1/NET33_XI45/XI1/MM3_d N_WL<86>_XI45/XI1/MM3_g
+ N_BLN<14>_XI45/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI1/MM0 N_XI45/XI1/NET34_XI45/XI1/MM0_d N_WL<86>_XI45/XI1/MM0_g
+ N_BL<14>_XI45/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI1/MM1 N_XI45/XI1/NET33_XI45/XI1/MM1_d N_XI45/XI1/NET34_XI45/XI1/MM1_g
+ N_VSS_XI45/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI1/MM9 N_XI45/XI1/NET36_XI45/XI1/MM9_d N_WL<87>_XI45/XI1/MM9_g
+ N_BL<14>_XI45/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI1/MM6 N_XI45/XI1/NET35_XI45/XI1/MM6_d N_XI45/XI1/NET36_XI45/XI1/MM6_g
+ N_VSS_XI45/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI1/MM7 N_XI45/XI1/NET36_XI45/XI1/MM7_d N_XI45/XI1/NET35_XI45/XI1/MM7_g
+ N_VSS_XI45/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI1/MM8 N_XI45/XI1/NET35_XI45/XI1/MM8_d N_WL<87>_XI45/XI1/MM8_g
+ N_BLN<14>_XI45/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI1/MM5 N_XI45/XI1/NET34_XI45/XI1/MM5_d N_XI45/XI1/NET33_XI45/XI1/MM5_g
+ N_VDD_XI45/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI1/MM4 N_XI45/XI1/NET33_XI45/XI1/MM4_d N_XI45/XI1/NET34_XI45/XI1/MM4_g
+ N_VDD_XI45/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI1/MM10 N_XI45/XI1/NET35_XI45/XI1/MM10_d N_XI45/XI1/NET36_XI45/XI1/MM10_g
+ N_VDD_XI45/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI1/MM11 N_XI45/XI1/NET36_XI45/XI1/MM11_d N_XI45/XI1/NET35_XI45/XI1/MM11_g
+ N_VDD_XI45/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI2/MM2 N_XI45/XI2/NET34_XI45/XI2/MM2_d N_XI45/XI2/NET33_XI45/XI2/MM2_g
+ N_VSS_XI45/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI2/MM3 N_XI45/XI2/NET33_XI45/XI2/MM3_d N_WL<86>_XI45/XI2/MM3_g
+ N_BLN<13>_XI45/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI2/MM0 N_XI45/XI2/NET34_XI45/XI2/MM0_d N_WL<86>_XI45/XI2/MM0_g
+ N_BL<13>_XI45/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI2/MM1 N_XI45/XI2/NET33_XI45/XI2/MM1_d N_XI45/XI2/NET34_XI45/XI2/MM1_g
+ N_VSS_XI45/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI2/MM9 N_XI45/XI2/NET36_XI45/XI2/MM9_d N_WL<87>_XI45/XI2/MM9_g
+ N_BL<13>_XI45/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI2/MM6 N_XI45/XI2/NET35_XI45/XI2/MM6_d N_XI45/XI2/NET36_XI45/XI2/MM6_g
+ N_VSS_XI45/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI2/MM7 N_XI45/XI2/NET36_XI45/XI2/MM7_d N_XI45/XI2/NET35_XI45/XI2/MM7_g
+ N_VSS_XI45/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI2/MM8 N_XI45/XI2/NET35_XI45/XI2/MM8_d N_WL<87>_XI45/XI2/MM8_g
+ N_BLN<13>_XI45/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI2/MM5 N_XI45/XI2/NET34_XI45/XI2/MM5_d N_XI45/XI2/NET33_XI45/XI2/MM5_g
+ N_VDD_XI45/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI2/MM4 N_XI45/XI2/NET33_XI45/XI2/MM4_d N_XI45/XI2/NET34_XI45/XI2/MM4_g
+ N_VDD_XI45/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI2/MM10 N_XI45/XI2/NET35_XI45/XI2/MM10_d N_XI45/XI2/NET36_XI45/XI2/MM10_g
+ N_VDD_XI45/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI2/MM11 N_XI45/XI2/NET36_XI45/XI2/MM11_d N_XI45/XI2/NET35_XI45/XI2/MM11_g
+ N_VDD_XI45/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI3/MM2 N_XI45/XI3/NET34_XI45/XI3/MM2_d N_XI45/XI3/NET33_XI45/XI3/MM2_g
+ N_VSS_XI45/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI3/MM3 N_XI45/XI3/NET33_XI45/XI3/MM3_d N_WL<86>_XI45/XI3/MM3_g
+ N_BLN<12>_XI45/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI3/MM0 N_XI45/XI3/NET34_XI45/XI3/MM0_d N_WL<86>_XI45/XI3/MM0_g
+ N_BL<12>_XI45/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI3/MM1 N_XI45/XI3/NET33_XI45/XI3/MM1_d N_XI45/XI3/NET34_XI45/XI3/MM1_g
+ N_VSS_XI45/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI3/MM9 N_XI45/XI3/NET36_XI45/XI3/MM9_d N_WL<87>_XI45/XI3/MM9_g
+ N_BL<12>_XI45/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI3/MM6 N_XI45/XI3/NET35_XI45/XI3/MM6_d N_XI45/XI3/NET36_XI45/XI3/MM6_g
+ N_VSS_XI45/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI3/MM7 N_XI45/XI3/NET36_XI45/XI3/MM7_d N_XI45/XI3/NET35_XI45/XI3/MM7_g
+ N_VSS_XI45/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI3/MM8 N_XI45/XI3/NET35_XI45/XI3/MM8_d N_WL<87>_XI45/XI3/MM8_g
+ N_BLN<12>_XI45/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI3/MM5 N_XI45/XI3/NET34_XI45/XI3/MM5_d N_XI45/XI3/NET33_XI45/XI3/MM5_g
+ N_VDD_XI45/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI3/MM4 N_XI45/XI3/NET33_XI45/XI3/MM4_d N_XI45/XI3/NET34_XI45/XI3/MM4_g
+ N_VDD_XI45/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI3/MM10 N_XI45/XI3/NET35_XI45/XI3/MM10_d N_XI45/XI3/NET36_XI45/XI3/MM10_g
+ N_VDD_XI45/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI3/MM11 N_XI45/XI3/NET36_XI45/XI3/MM11_d N_XI45/XI3/NET35_XI45/XI3/MM11_g
+ N_VDD_XI45/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI4/MM2 N_XI45/XI4/NET34_XI45/XI4/MM2_d N_XI45/XI4/NET33_XI45/XI4/MM2_g
+ N_VSS_XI45/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI4/MM3 N_XI45/XI4/NET33_XI45/XI4/MM3_d N_WL<86>_XI45/XI4/MM3_g
+ N_BLN<11>_XI45/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI4/MM0 N_XI45/XI4/NET34_XI45/XI4/MM0_d N_WL<86>_XI45/XI4/MM0_g
+ N_BL<11>_XI45/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI4/MM1 N_XI45/XI4/NET33_XI45/XI4/MM1_d N_XI45/XI4/NET34_XI45/XI4/MM1_g
+ N_VSS_XI45/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI4/MM9 N_XI45/XI4/NET36_XI45/XI4/MM9_d N_WL<87>_XI45/XI4/MM9_g
+ N_BL<11>_XI45/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI4/MM6 N_XI45/XI4/NET35_XI45/XI4/MM6_d N_XI45/XI4/NET36_XI45/XI4/MM6_g
+ N_VSS_XI45/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI4/MM7 N_XI45/XI4/NET36_XI45/XI4/MM7_d N_XI45/XI4/NET35_XI45/XI4/MM7_g
+ N_VSS_XI45/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI4/MM8 N_XI45/XI4/NET35_XI45/XI4/MM8_d N_WL<87>_XI45/XI4/MM8_g
+ N_BLN<11>_XI45/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI4/MM5 N_XI45/XI4/NET34_XI45/XI4/MM5_d N_XI45/XI4/NET33_XI45/XI4/MM5_g
+ N_VDD_XI45/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI4/MM4 N_XI45/XI4/NET33_XI45/XI4/MM4_d N_XI45/XI4/NET34_XI45/XI4/MM4_g
+ N_VDD_XI45/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI4/MM10 N_XI45/XI4/NET35_XI45/XI4/MM10_d N_XI45/XI4/NET36_XI45/XI4/MM10_g
+ N_VDD_XI45/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI4/MM11 N_XI45/XI4/NET36_XI45/XI4/MM11_d N_XI45/XI4/NET35_XI45/XI4/MM11_g
+ N_VDD_XI45/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI5/MM2 N_XI45/XI5/NET34_XI45/XI5/MM2_d N_XI45/XI5/NET33_XI45/XI5/MM2_g
+ N_VSS_XI45/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI5/MM3 N_XI45/XI5/NET33_XI45/XI5/MM3_d N_WL<86>_XI45/XI5/MM3_g
+ N_BLN<10>_XI45/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI5/MM0 N_XI45/XI5/NET34_XI45/XI5/MM0_d N_WL<86>_XI45/XI5/MM0_g
+ N_BL<10>_XI45/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI5/MM1 N_XI45/XI5/NET33_XI45/XI5/MM1_d N_XI45/XI5/NET34_XI45/XI5/MM1_g
+ N_VSS_XI45/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI5/MM9 N_XI45/XI5/NET36_XI45/XI5/MM9_d N_WL<87>_XI45/XI5/MM9_g
+ N_BL<10>_XI45/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI5/MM6 N_XI45/XI5/NET35_XI45/XI5/MM6_d N_XI45/XI5/NET36_XI45/XI5/MM6_g
+ N_VSS_XI45/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI5/MM7 N_XI45/XI5/NET36_XI45/XI5/MM7_d N_XI45/XI5/NET35_XI45/XI5/MM7_g
+ N_VSS_XI45/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI5/MM8 N_XI45/XI5/NET35_XI45/XI5/MM8_d N_WL<87>_XI45/XI5/MM8_g
+ N_BLN<10>_XI45/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI5/MM5 N_XI45/XI5/NET34_XI45/XI5/MM5_d N_XI45/XI5/NET33_XI45/XI5/MM5_g
+ N_VDD_XI45/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI5/MM4 N_XI45/XI5/NET33_XI45/XI5/MM4_d N_XI45/XI5/NET34_XI45/XI5/MM4_g
+ N_VDD_XI45/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI5/MM10 N_XI45/XI5/NET35_XI45/XI5/MM10_d N_XI45/XI5/NET36_XI45/XI5/MM10_g
+ N_VDD_XI45/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI5/MM11 N_XI45/XI5/NET36_XI45/XI5/MM11_d N_XI45/XI5/NET35_XI45/XI5/MM11_g
+ N_VDD_XI45/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI6/MM2 N_XI45/XI6/NET34_XI45/XI6/MM2_d N_XI45/XI6/NET33_XI45/XI6/MM2_g
+ N_VSS_XI45/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM3 N_XI45/XI6/NET33_XI45/XI6/MM3_d N_WL<86>_XI45/XI6/MM3_g
+ N_BLN<9>_XI45/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM0 N_XI45/XI6/NET34_XI45/XI6/MM0_d N_WL<86>_XI45/XI6/MM0_g
+ N_BL<9>_XI45/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM1 N_XI45/XI6/NET33_XI45/XI6/MM1_d N_XI45/XI6/NET34_XI45/XI6/MM1_g
+ N_VSS_XI45/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM9 N_XI45/XI6/NET36_XI45/XI6/MM9_d N_WL<87>_XI45/XI6/MM9_g
+ N_BL<9>_XI45/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM6 N_XI45/XI6/NET35_XI45/XI6/MM6_d N_XI45/XI6/NET36_XI45/XI6/MM6_g
+ N_VSS_XI45/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM7 N_XI45/XI6/NET36_XI45/XI6/MM7_d N_XI45/XI6/NET35_XI45/XI6/MM7_g
+ N_VSS_XI45/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM8 N_XI45/XI6/NET35_XI45/XI6/MM8_d N_WL<87>_XI45/XI6/MM8_g
+ N_BLN<9>_XI45/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI6/MM5 N_XI45/XI6/NET34_XI45/XI6/MM5_d N_XI45/XI6/NET33_XI45/XI6/MM5_g
+ N_VDD_XI45/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI6/MM4 N_XI45/XI6/NET33_XI45/XI6/MM4_d N_XI45/XI6/NET34_XI45/XI6/MM4_g
+ N_VDD_XI45/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI6/MM10 N_XI45/XI6/NET35_XI45/XI6/MM10_d N_XI45/XI6/NET36_XI45/XI6/MM10_g
+ N_VDD_XI45/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI6/MM11 N_XI45/XI6/NET36_XI45/XI6/MM11_d N_XI45/XI6/NET35_XI45/XI6/MM11_g
+ N_VDD_XI45/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI7/MM2 N_XI45/XI7/NET34_XI45/XI7/MM2_d N_XI45/XI7/NET33_XI45/XI7/MM2_g
+ N_VSS_XI45/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM3 N_XI45/XI7/NET33_XI45/XI7/MM3_d N_WL<86>_XI45/XI7/MM3_g
+ N_BLN<8>_XI45/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM0 N_XI45/XI7/NET34_XI45/XI7/MM0_d N_WL<86>_XI45/XI7/MM0_g
+ N_BL<8>_XI45/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM1 N_XI45/XI7/NET33_XI45/XI7/MM1_d N_XI45/XI7/NET34_XI45/XI7/MM1_g
+ N_VSS_XI45/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM9 N_XI45/XI7/NET36_XI45/XI7/MM9_d N_WL<87>_XI45/XI7/MM9_g
+ N_BL<8>_XI45/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM6 N_XI45/XI7/NET35_XI45/XI7/MM6_d N_XI45/XI7/NET36_XI45/XI7/MM6_g
+ N_VSS_XI45/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM7 N_XI45/XI7/NET36_XI45/XI7/MM7_d N_XI45/XI7/NET35_XI45/XI7/MM7_g
+ N_VSS_XI45/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM8 N_XI45/XI7/NET35_XI45/XI7/MM8_d N_WL<87>_XI45/XI7/MM8_g
+ N_BLN<8>_XI45/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI7/MM5 N_XI45/XI7/NET34_XI45/XI7/MM5_d N_XI45/XI7/NET33_XI45/XI7/MM5_g
+ N_VDD_XI45/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI7/MM4 N_XI45/XI7/NET33_XI45/XI7/MM4_d N_XI45/XI7/NET34_XI45/XI7/MM4_g
+ N_VDD_XI45/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI7/MM10 N_XI45/XI7/NET35_XI45/XI7/MM10_d N_XI45/XI7/NET36_XI45/XI7/MM10_g
+ N_VDD_XI45/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI7/MM11 N_XI45/XI7/NET36_XI45/XI7/MM11_d N_XI45/XI7/NET35_XI45/XI7/MM11_g
+ N_VDD_XI45/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI8/MM2 N_XI45/XI8/NET34_XI45/XI8/MM2_d N_XI45/XI8/NET33_XI45/XI8/MM2_g
+ N_VSS_XI45/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM3 N_XI45/XI8/NET33_XI45/XI8/MM3_d N_WL<86>_XI45/XI8/MM3_g
+ N_BLN<7>_XI45/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM0 N_XI45/XI8/NET34_XI45/XI8/MM0_d N_WL<86>_XI45/XI8/MM0_g
+ N_BL<7>_XI45/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM1 N_XI45/XI8/NET33_XI45/XI8/MM1_d N_XI45/XI8/NET34_XI45/XI8/MM1_g
+ N_VSS_XI45/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM9 N_XI45/XI8/NET36_XI45/XI8/MM9_d N_WL<87>_XI45/XI8/MM9_g
+ N_BL<7>_XI45/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM6 N_XI45/XI8/NET35_XI45/XI8/MM6_d N_XI45/XI8/NET36_XI45/XI8/MM6_g
+ N_VSS_XI45/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM7 N_XI45/XI8/NET36_XI45/XI8/MM7_d N_XI45/XI8/NET35_XI45/XI8/MM7_g
+ N_VSS_XI45/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM8 N_XI45/XI8/NET35_XI45/XI8/MM8_d N_WL<87>_XI45/XI8/MM8_g
+ N_BLN<7>_XI45/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI8/MM5 N_XI45/XI8/NET34_XI45/XI8/MM5_d N_XI45/XI8/NET33_XI45/XI8/MM5_g
+ N_VDD_XI45/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI8/MM4 N_XI45/XI8/NET33_XI45/XI8/MM4_d N_XI45/XI8/NET34_XI45/XI8/MM4_g
+ N_VDD_XI45/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI8/MM10 N_XI45/XI8/NET35_XI45/XI8/MM10_d N_XI45/XI8/NET36_XI45/XI8/MM10_g
+ N_VDD_XI45/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI8/MM11 N_XI45/XI8/NET36_XI45/XI8/MM11_d N_XI45/XI8/NET35_XI45/XI8/MM11_g
+ N_VDD_XI45/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI9/MM2 N_XI45/XI9/NET34_XI45/XI9/MM2_d N_XI45/XI9/NET33_XI45/XI9/MM2_g
+ N_VSS_XI45/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM3 N_XI45/XI9/NET33_XI45/XI9/MM3_d N_WL<86>_XI45/XI9/MM3_g
+ N_BLN<6>_XI45/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM0 N_XI45/XI9/NET34_XI45/XI9/MM0_d N_WL<86>_XI45/XI9/MM0_g
+ N_BL<6>_XI45/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM1 N_XI45/XI9/NET33_XI45/XI9/MM1_d N_XI45/XI9/NET34_XI45/XI9/MM1_g
+ N_VSS_XI45/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM9 N_XI45/XI9/NET36_XI45/XI9/MM9_d N_WL<87>_XI45/XI9/MM9_g
+ N_BL<6>_XI45/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM6 N_XI45/XI9/NET35_XI45/XI9/MM6_d N_XI45/XI9/NET36_XI45/XI9/MM6_g
+ N_VSS_XI45/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM7 N_XI45/XI9/NET36_XI45/XI9/MM7_d N_XI45/XI9/NET35_XI45/XI9/MM7_g
+ N_VSS_XI45/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM8 N_XI45/XI9/NET35_XI45/XI9/MM8_d N_WL<87>_XI45/XI9/MM8_g
+ N_BLN<6>_XI45/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI9/MM5 N_XI45/XI9/NET34_XI45/XI9/MM5_d N_XI45/XI9/NET33_XI45/XI9/MM5_g
+ N_VDD_XI45/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI9/MM4 N_XI45/XI9/NET33_XI45/XI9/MM4_d N_XI45/XI9/NET34_XI45/XI9/MM4_g
+ N_VDD_XI45/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI9/MM10 N_XI45/XI9/NET35_XI45/XI9/MM10_d N_XI45/XI9/NET36_XI45/XI9/MM10_g
+ N_VDD_XI45/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI9/MM11 N_XI45/XI9/NET36_XI45/XI9/MM11_d N_XI45/XI9/NET35_XI45/XI9/MM11_g
+ N_VDD_XI45/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI10/MM2 N_XI45/XI10/NET34_XI45/XI10/MM2_d
+ N_XI45/XI10/NET33_XI45/XI10/MM2_g N_VSS_XI45/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI10/MM3 N_XI45/XI10/NET33_XI45/XI10/MM3_d N_WL<86>_XI45/XI10/MM3_g
+ N_BLN<5>_XI45/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI10/MM0 N_XI45/XI10/NET34_XI45/XI10/MM0_d N_WL<86>_XI45/XI10/MM0_g
+ N_BL<5>_XI45/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI10/MM1 N_XI45/XI10/NET33_XI45/XI10/MM1_d
+ N_XI45/XI10/NET34_XI45/XI10/MM1_g N_VSS_XI45/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI10/MM9 N_XI45/XI10/NET36_XI45/XI10/MM9_d N_WL<87>_XI45/XI10/MM9_g
+ N_BL<5>_XI45/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI10/MM6 N_XI45/XI10/NET35_XI45/XI10/MM6_d
+ N_XI45/XI10/NET36_XI45/XI10/MM6_g N_VSS_XI45/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI10/MM7 N_XI45/XI10/NET36_XI45/XI10/MM7_d
+ N_XI45/XI10/NET35_XI45/XI10/MM7_g N_VSS_XI45/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI10/MM8 N_XI45/XI10/NET35_XI45/XI10/MM8_d N_WL<87>_XI45/XI10/MM8_g
+ N_BLN<5>_XI45/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI10/MM5 N_XI45/XI10/NET34_XI45/XI10/MM5_d
+ N_XI45/XI10/NET33_XI45/XI10/MM5_g N_VDD_XI45/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI10/MM4 N_XI45/XI10/NET33_XI45/XI10/MM4_d
+ N_XI45/XI10/NET34_XI45/XI10/MM4_g N_VDD_XI45/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI10/MM10 N_XI45/XI10/NET35_XI45/XI10/MM10_d
+ N_XI45/XI10/NET36_XI45/XI10/MM10_g N_VDD_XI45/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI10/MM11 N_XI45/XI10/NET36_XI45/XI10/MM11_d
+ N_XI45/XI10/NET35_XI45/XI10/MM11_g N_VDD_XI45/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI11/MM2 N_XI45/XI11/NET34_XI45/XI11/MM2_d
+ N_XI45/XI11/NET33_XI45/XI11/MM2_g N_VSS_XI45/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI11/MM3 N_XI45/XI11/NET33_XI45/XI11/MM3_d N_WL<86>_XI45/XI11/MM3_g
+ N_BLN<4>_XI45/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI11/MM0 N_XI45/XI11/NET34_XI45/XI11/MM0_d N_WL<86>_XI45/XI11/MM0_g
+ N_BL<4>_XI45/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI11/MM1 N_XI45/XI11/NET33_XI45/XI11/MM1_d
+ N_XI45/XI11/NET34_XI45/XI11/MM1_g N_VSS_XI45/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI11/MM9 N_XI45/XI11/NET36_XI45/XI11/MM9_d N_WL<87>_XI45/XI11/MM9_g
+ N_BL<4>_XI45/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI11/MM6 N_XI45/XI11/NET35_XI45/XI11/MM6_d
+ N_XI45/XI11/NET36_XI45/XI11/MM6_g N_VSS_XI45/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI11/MM7 N_XI45/XI11/NET36_XI45/XI11/MM7_d
+ N_XI45/XI11/NET35_XI45/XI11/MM7_g N_VSS_XI45/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI11/MM8 N_XI45/XI11/NET35_XI45/XI11/MM8_d N_WL<87>_XI45/XI11/MM8_g
+ N_BLN<4>_XI45/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI11/MM5 N_XI45/XI11/NET34_XI45/XI11/MM5_d
+ N_XI45/XI11/NET33_XI45/XI11/MM5_g N_VDD_XI45/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI11/MM4 N_XI45/XI11/NET33_XI45/XI11/MM4_d
+ N_XI45/XI11/NET34_XI45/XI11/MM4_g N_VDD_XI45/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI11/MM10 N_XI45/XI11/NET35_XI45/XI11/MM10_d
+ N_XI45/XI11/NET36_XI45/XI11/MM10_g N_VDD_XI45/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI11/MM11 N_XI45/XI11/NET36_XI45/XI11/MM11_d
+ N_XI45/XI11/NET35_XI45/XI11/MM11_g N_VDD_XI45/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI12/MM2 N_XI45/XI12/NET34_XI45/XI12/MM2_d
+ N_XI45/XI12/NET33_XI45/XI12/MM2_g N_VSS_XI45/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI12/MM3 N_XI45/XI12/NET33_XI45/XI12/MM3_d N_WL<86>_XI45/XI12/MM3_g
+ N_BLN<3>_XI45/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI12/MM0 N_XI45/XI12/NET34_XI45/XI12/MM0_d N_WL<86>_XI45/XI12/MM0_g
+ N_BL<3>_XI45/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI12/MM1 N_XI45/XI12/NET33_XI45/XI12/MM1_d
+ N_XI45/XI12/NET34_XI45/XI12/MM1_g N_VSS_XI45/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI12/MM9 N_XI45/XI12/NET36_XI45/XI12/MM9_d N_WL<87>_XI45/XI12/MM9_g
+ N_BL<3>_XI45/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI12/MM6 N_XI45/XI12/NET35_XI45/XI12/MM6_d
+ N_XI45/XI12/NET36_XI45/XI12/MM6_g N_VSS_XI45/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI12/MM7 N_XI45/XI12/NET36_XI45/XI12/MM7_d
+ N_XI45/XI12/NET35_XI45/XI12/MM7_g N_VSS_XI45/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI12/MM8 N_XI45/XI12/NET35_XI45/XI12/MM8_d N_WL<87>_XI45/XI12/MM8_g
+ N_BLN<3>_XI45/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI12/MM5 N_XI45/XI12/NET34_XI45/XI12/MM5_d
+ N_XI45/XI12/NET33_XI45/XI12/MM5_g N_VDD_XI45/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI12/MM4 N_XI45/XI12/NET33_XI45/XI12/MM4_d
+ N_XI45/XI12/NET34_XI45/XI12/MM4_g N_VDD_XI45/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI12/MM10 N_XI45/XI12/NET35_XI45/XI12/MM10_d
+ N_XI45/XI12/NET36_XI45/XI12/MM10_g N_VDD_XI45/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI12/MM11 N_XI45/XI12/NET36_XI45/XI12/MM11_d
+ N_XI45/XI12/NET35_XI45/XI12/MM11_g N_VDD_XI45/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI13/MM2 N_XI45/XI13/NET34_XI45/XI13/MM2_d
+ N_XI45/XI13/NET33_XI45/XI13/MM2_g N_VSS_XI45/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI13/MM3 N_XI45/XI13/NET33_XI45/XI13/MM3_d N_WL<86>_XI45/XI13/MM3_g
+ N_BLN<2>_XI45/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI13/MM0 N_XI45/XI13/NET34_XI45/XI13/MM0_d N_WL<86>_XI45/XI13/MM0_g
+ N_BL<2>_XI45/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI13/MM1 N_XI45/XI13/NET33_XI45/XI13/MM1_d
+ N_XI45/XI13/NET34_XI45/XI13/MM1_g N_VSS_XI45/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI13/MM9 N_XI45/XI13/NET36_XI45/XI13/MM9_d N_WL<87>_XI45/XI13/MM9_g
+ N_BL<2>_XI45/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI13/MM6 N_XI45/XI13/NET35_XI45/XI13/MM6_d
+ N_XI45/XI13/NET36_XI45/XI13/MM6_g N_VSS_XI45/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI13/MM7 N_XI45/XI13/NET36_XI45/XI13/MM7_d
+ N_XI45/XI13/NET35_XI45/XI13/MM7_g N_VSS_XI45/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI13/MM8 N_XI45/XI13/NET35_XI45/XI13/MM8_d N_WL<87>_XI45/XI13/MM8_g
+ N_BLN<2>_XI45/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI13/MM5 N_XI45/XI13/NET34_XI45/XI13/MM5_d
+ N_XI45/XI13/NET33_XI45/XI13/MM5_g N_VDD_XI45/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI13/MM4 N_XI45/XI13/NET33_XI45/XI13/MM4_d
+ N_XI45/XI13/NET34_XI45/XI13/MM4_g N_VDD_XI45/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI13/MM10 N_XI45/XI13/NET35_XI45/XI13/MM10_d
+ N_XI45/XI13/NET36_XI45/XI13/MM10_g N_VDD_XI45/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI13/MM11 N_XI45/XI13/NET36_XI45/XI13/MM11_d
+ N_XI45/XI13/NET35_XI45/XI13/MM11_g N_VDD_XI45/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI14/MM2 N_XI45/XI14/NET34_XI45/XI14/MM2_d
+ N_XI45/XI14/NET33_XI45/XI14/MM2_g N_VSS_XI45/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI14/MM3 N_XI45/XI14/NET33_XI45/XI14/MM3_d N_WL<86>_XI45/XI14/MM3_g
+ N_BLN<1>_XI45/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI14/MM0 N_XI45/XI14/NET34_XI45/XI14/MM0_d N_WL<86>_XI45/XI14/MM0_g
+ N_BL<1>_XI45/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI14/MM1 N_XI45/XI14/NET33_XI45/XI14/MM1_d
+ N_XI45/XI14/NET34_XI45/XI14/MM1_g N_VSS_XI45/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI14/MM9 N_XI45/XI14/NET36_XI45/XI14/MM9_d N_WL<87>_XI45/XI14/MM9_g
+ N_BL<1>_XI45/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI14/MM6 N_XI45/XI14/NET35_XI45/XI14/MM6_d
+ N_XI45/XI14/NET36_XI45/XI14/MM6_g N_VSS_XI45/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI14/MM7 N_XI45/XI14/NET36_XI45/XI14/MM7_d
+ N_XI45/XI14/NET35_XI45/XI14/MM7_g N_VSS_XI45/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI14/MM8 N_XI45/XI14/NET35_XI45/XI14/MM8_d N_WL<87>_XI45/XI14/MM8_g
+ N_BLN<1>_XI45/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI14/MM5 N_XI45/XI14/NET34_XI45/XI14/MM5_d
+ N_XI45/XI14/NET33_XI45/XI14/MM5_g N_VDD_XI45/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI14/MM4 N_XI45/XI14/NET33_XI45/XI14/MM4_d
+ N_XI45/XI14/NET34_XI45/XI14/MM4_g N_VDD_XI45/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI14/MM10 N_XI45/XI14/NET35_XI45/XI14/MM10_d
+ N_XI45/XI14/NET36_XI45/XI14/MM10_g N_VDD_XI45/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI14/MM11 N_XI45/XI14/NET36_XI45/XI14/MM11_d
+ N_XI45/XI14/NET35_XI45/XI14/MM11_g N_VDD_XI45/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI15/MM2 N_XI45/XI15/NET34_XI45/XI15/MM2_d
+ N_XI45/XI15/NET33_XI45/XI15/MM2_g N_VSS_XI45/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI15/MM3 N_XI45/XI15/NET33_XI45/XI15/MM3_d N_WL<86>_XI45/XI15/MM3_g
+ N_BLN<0>_XI45/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI15/MM0 N_XI45/XI15/NET34_XI45/XI15/MM0_d N_WL<86>_XI45/XI15/MM0_g
+ N_BL<0>_XI45/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI15/MM1 N_XI45/XI15/NET33_XI45/XI15/MM1_d
+ N_XI45/XI15/NET34_XI45/XI15/MM1_g N_VSS_XI45/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI15/MM9 N_XI45/XI15/NET36_XI45/XI15/MM9_d N_WL<87>_XI45/XI15/MM9_g
+ N_BL<0>_XI45/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI15/MM6 N_XI45/XI15/NET35_XI45/XI15/MM6_d
+ N_XI45/XI15/NET36_XI45/XI15/MM6_g N_VSS_XI45/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI15/MM7 N_XI45/XI15/NET36_XI45/XI15/MM7_d
+ N_XI45/XI15/NET35_XI45/XI15/MM7_g N_VSS_XI45/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI45/XI15/MM8 N_XI45/XI15/NET35_XI45/XI15/MM8_d N_WL<87>_XI45/XI15/MM8_g
+ N_BLN<0>_XI45/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI45/XI15/MM5 N_XI45/XI15/NET34_XI45/XI15/MM5_d
+ N_XI45/XI15/NET33_XI45/XI15/MM5_g N_VDD_XI45/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI15/MM4 N_XI45/XI15/NET33_XI45/XI15/MM4_d
+ N_XI45/XI15/NET34_XI45/XI15/MM4_g N_VDD_XI45/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI15/MM10 N_XI45/XI15/NET35_XI45/XI15/MM10_d
+ N_XI45/XI15/NET36_XI45/XI15/MM10_g N_VDD_XI45/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI45/XI15/MM11 N_XI45/XI15/NET36_XI45/XI15/MM11_d
+ N_XI45/XI15/NET35_XI45/XI15/MM11_g N_VDD_XI45/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI0/MM2 N_XI46/XI0/NET34_XI46/XI0/MM2_d N_XI46/XI0/NET33_XI46/XI0/MM2_g
+ N_VSS_XI46/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI0/MM3 N_XI46/XI0/NET33_XI46/XI0/MM3_d N_WL<88>_XI46/XI0/MM3_g
+ N_BLN<15>_XI46/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI0/MM0 N_XI46/XI0/NET34_XI46/XI0/MM0_d N_WL<88>_XI46/XI0/MM0_g
+ N_BL<15>_XI46/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI0/MM1 N_XI46/XI0/NET33_XI46/XI0/MM1_d N_XI46/XI0/NET34_XI46/XI0/MM1_g
+ N_VSS_XI46/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI0/MM9 N_XI46/XI0/NET36_XI46/XI0/MM9_d N_WL<89>_XI46/XI0/MM9_g
+ N_BL<15>_XI46/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI0/MM6 N_XI46/XI0/NET35_XI46/XI0/MM6_d N_XI46/XI0/NET36_XI46/XI0/MM6_g
+ N_VSS_XI46/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI0/MM7 N_XI46/XI0/NET36_XI46/XI0/MM7_d N_XI46/XI0/NET35_XI46/XI0/MM7_g
+ N_VSS_XI46/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI0/MM8 N_XI46/XI0/NET35_XI46/XI0/MM8_d N_WL<89>_XI46/XI0/MM8_g
+ N_BLN<15>_XI46/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI0/MM5 N_XI46/XI0/NET34_XI46/XI0/MM5_d N_XI46/XI0/NET33_XI46/XI0/MM5_g
+ N_VDD_XI46/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI0/MM4 N_XI46/XI0/NET33_XI46/XI0/MM4_d N_XI46/XI0/NET34_XI46/XI0/MM4_g
+ N_VDD_XI46/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI0/MM10 N_XI46/XI0/NET35_XI46/XI0/MM10_d N_XI46/XI0/NET36_XI46/XI0/MM10_g
+ N_VDD_XI46/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI0/MM11 N_XI46/XI0/NET36_XI46/XI0/MM11_d N_XI46/XI0/NET35_XI46/XI0/MM11_g
+ N_VDD_XI46/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI1/MM2 N_XI46/XI1/NET34_XI46/XI1/MM2_d N_XI46/XI1/NET33_XI46/XI1/MM2_g
+ N_VSS_XI46/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI1/MM3 N_XI46/XI1/NET33_XI46/XI1/MM3_d N_WL<88>_XI46/XI1/MM3_g
+ N_BLN<14>_XI46/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI1/MM0 N_XI46/XI1/NET34_XI46/XI1/MM0_d N_WL<88>_XI46/XI1/MM0_g
+ N_BL<14>_XI46/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI1/MM1 N_XI46/XI1/NET33_XI46/XI1/MM1_d N_XI46/XI1/NET34_XI46/XI1/MM1_g
+ N_VSS_XI46/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI1/MM9 N_XI46/XI1/NET36_XI46/XI1/MM9_d N_WL<89>_XI46/XI1/MM9_g
+ N_BL<14>_XI46/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI1/MM6 N_XI46/XI1/NET35_XI46/XI1/MM6_d N_XI46/XI1/NET36_XI46/XI1/MM6_g
+ N_VSS_XI46/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI1/MM7 N_XI46/XI1/NET36_XI46/XI1/MM7_d N_XI46/XI1/NET35_XI46/XI1/MM7_g
+ N_VSS_XI46/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI1/MM8 N_XI46/XI1/NET35_XI46/XI1/MM8_d N_WL<89>_XI46/XI1/MM8_g
+ N_BLN<14>_XI46/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI1/MM5 N_XI46/XI1/NET34_XI46/XI1/MM5_d N_XI46/XI1/NET33_XI46/XI1/MM5_g
+ N_VDD_XI46/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI1/MM4 N_XI46/XI1/NET33_XI46/XI1/MM4_d N_XI46/XI1/NET34_XI46/XI1/MM4_g
+ N_VDD_XI46/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI1/MM10 N_XI46/XI1/NET35_XI46/XI1/MM10_d N_XI46/XI1/NET36_XI46/XI1/MM10_g
+ N_VDD_XI46/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI1/MM11 N_XI46/XI1/NET36_XI46/XI1/MM11_d N_XI46/XI1/NET35_XI46/XI1/MM11_g
+ N_VDD_XI46/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI2/MM2 N_XI46/XI2/NET34_XI46/XI2/MM2_d N_XI46/XI2/NET33_XI46/XI2/MM2_g
+ N_VSS_XI46/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI2/MM3 N_XI46/XI2/NET33_XI46/XI2/MM3_d N_WL<88>_XI46/XI2/MM3_g
+ N_BLN<13>_XI46/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI2/MM0 N_XI46/XI2/NET34_XI46/XI2/MM0_d N_WL<88>_XI46/XI2/MM0_g
+ N_BL<13>_XI46/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI2/MM1 N_XI46/XI2/NET33_XI46/XI2/MM1_d N_XI46/XI2/NET34_XI46/XI2/MM1_g
+ N_VSS_XI46/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI2/MM9 N_XI46/XI2/NET36_XI46/XI2/MM9_d N_WL<89>_XI46/XI2/MM9_g
+ N_BL<13>_XI46/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI2/MM6 N_XI46/XI2/NET35_XI46/XI2/MM6_d N_XI46/XI2/NET36_XI46/XI2/MM6_g
+ N_VSS_XI46/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI2/MM7 N_XI46/XI2/NET36_XI46/XI2/MM7_d N_XI46/XI2/NET35_XI46/XI2/MM7_g
+ N_VSS_XI46/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI2/MM8 N_XI46/XI2/NET35_XI46/XI2/MM8_d N_WL<89>_XI46/XI2/MM8_g
+ N_BLN<13>_XI46/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI2/MM5 N_XI46/XI2/NET34_XI46/XI2/MM5_d N_XI46/XI2/NET33_XI46/XI2/MM5_g
+ N_VDD_XI46/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI2/MM4 N_XI46/XI2/NET33_XI46/XI2/MM4_d N_XI46/XI2/NET34_XI46/XI2/MM4_g
+ N_VDD_XI46/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI2/MM10 N_XI46/XI2/NET35_XI46/XI2/MM10_d N_XI46/XI2/NET36_XI46/XI2/MM10_g
+ N_VDD_XI46/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI2/MM11 N_XI46/XI2/NET36_XI46/XI2/MM11_d N_XI46/XI2/NET35_XI46/XI2/MM11_g
+ N_VDD_XI46/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI3/MM2 N_XI46/XI3/NET34_XI46/XI3/MM2_d N_XI46/XI3/NET33_XI46/XI3/MM2_g
+ N_VSS_XI46/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI3/MM3 N_XI46/XI3/NET33_XI46/XI3/MM3_d N_WL<88>_XI46/XI3/MM3_g
+ N_BLN<12>_XI46/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI3/MM0 N_XI46/XI3/NET34_XI46/XI3/MM0_d N_WL<88>_XI46/XI3/MM0_g
+ N_BL<12>_XI46/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI3/MM1 N_XI46/XI3/NET33_XI46/XI3/MM1_d N_XI46/XI3/NET34_XI46/XI3/MM1_g
+ N_VSS_XI46/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI3/MM9 N_XI46/XI3/NET36_XI46/XI3/MM9_d N_WL<89>_XI46/XI3/MM9_g
+ N_BL<12>_XI46/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI3/MM6 N_XI46/XI3/NET35_XI46/XI3/MM6_d N_XI46/XI3/NET36_XI46/XI3/MM6_g
+ N_VSS_XI46/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI3/MM7 N_XI46/XI3/NET36_XI46/XI3/MM7_d N_XI46/XI3/NET35_XI46/XI3/MM7_g
+ N_VSS_XI46/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI3/MM8 N_XI46/XI3/NET35_XI46/XI3/MM8_d N_WL<89>_XI46/XI3/MM8_g
+ N_BLN<12>_XI46/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI3/MM5 N_XI46/XI3/NET34_XI46/XI3/MM5_d N_XI46/XI3/NET33_XI46/XI3/MM5_g
+ N_VDD_XI46/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI3/MM4 N_XI46/XI3/NET33_XI46/XI3/MM4_d N_XI46/XI3/NET34_XI46/XI3/MM4_g
+ N_VDD_XI46/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI3/MM10 N_XI46/XI3/NET35_XI46/XI3/MM10_d N_XI46/XI3/NET36_XI46/XI3/MM10_g
+ N_VDD_XI46/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI3/MM11 N_XI46/XI3/NET36_XI46/XI3/MM11_d N_XI46/XI3/NET35_XI46/XI3/MM11_g
+ N_VDD_XI46/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI4/MM2 N_XI46/XI4/NET34_XI46/XI4/MM2_d N_XI46/XI4/NET33_XI46/XI4/MM2_g
+ N_VSS_XI46/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI4/MM3 N_XI46/XI4/NET33_XI46/XI4/MM3_d N_WL<88>_XI46/XI4/MM3_g
+ N_BLN<11>_XI46/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI4/MM0 N_XI46/XI4/NET34_XI46/XI4/MM0_d N_WL<88>_XI46/XI4/MM0_g
+ N_BL<11>_XI46/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI4/MM1 N_XI46/XI4/NET33_XI46/XI4/MM1_d N_XI46/XI4/NET34_XI46/XI4/MM1_g
+ N_VSS_XI46/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI4/MM9 N_XI46/XI4/NET36_XI46/XI4/MM9_d N_WL<89>_XI46/XI4/MM9_g
+ N_BL<11>_XI46/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI4/MM6 N_XI46/XI4/NET35_XI46/XI4/MM6_d N_XI46/XI4/NET36_XI46/XI4/MM6_g
+ N_VSS_XI46/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI4/MM7 N_XI46/XI4/NET36_XI46/XI4/MM7_d N_XI46/XI4/NET35_XI46/XI4/MM7_g
+ N_VSS_XI46/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI4/MM8 N_XI46/XI4/NET35_XI46/XI4/MM8_d N_WL<89>_XI46/XI4/MM8_g
+ N_BLN<11>_XI46/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI4/MM5 N_XI46/XI4/NET34_XI46/XI4/MM5_d N_XI46/XI4/NET33_XI46/XI4/MM5_g
+ N_VDD_XI46/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI4/MM4 N_XI46/XI4/NET33_XI46/XI4/MM4_d N_XI46/XI4/NET34_XI46/XI4/MM4_g
+ N_VDD_XI46/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI4/MM10 N_XI46/XI4/NET35_XI46/XI4/MM10_d N_XI46/XI4/NET36_XI46/XI4/MM10_g
+ N_VDD_XI46/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI4/MM11 N_XI46/XI4/NET36_XI46/XI4/MM11_d N_XI46/XI4/NET35_XI46/XI4/MM11_g
+ N_VDD_XI46/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI5/MM2 N_XI46/XI5/NET34_XI46/XI5/MM2_d N_XI46/XI5/NET33_XI46/XI5/MM2_g
+ N_VSS_XI46/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI5/MM3 N_XI46/XI5/NET33_XI46/XI5/MM3_d N_WL<88>_XI46/XI5/MM3_g
+ N_BLN<10>_XI46/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI5/MM0 N_XI46/XI5/NET34_XI46/XI5/MM0_d N_WL<88>_XI46/XI5/MM0_g
+ N_BL<10>_XI46/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI5/MM1 N_XI46/XI5/NET33_XI46/XI5/MM1_d N_XI46/XI5/NET34_XI46/XI5/MM1_g
+ N_VSS_XI46/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI5/MM9 N_XI46/XI5/NET36_XI46/XI5/MM9_d N_WL<89>_XI46/XI5/MM9_g
+ N_BL<10>_XI46/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI5/MM6 N_XI46/XI5/NET35_XI46/XI5/MM6_d N_XI46/XI5/NET36_XI46/XI5/MM6_g
+ N_VSS_XI46/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI5/MM7 N_XI46/XI5/NET36_XI46/XI5/MM7_d N_XI46/XI5/NET35_XI46/XI5/MM7_g
+ N_VSS_XI46/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI5/MM8 N_XI46/XI5/NET35_XI46/XI5/MM8_d N_WL<89>_XI46/XI5/MM8_g
+ N_BLN<10>_XI46/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI5/MM5 N_XI46/XI5/NET34_XI46/XI5/MM5_d N_XI46/XI5/NET33_XI46/XI5/MM5_g
+ N_VDD_XI46/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI5/MM4 N_XI46/XI5/NET33_XI46/XI5/MM4_d N_XI46/XI5/NET34_XI46/XI5/MM4_g
+ N_VDD_XI46/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI5/MM10 N_XI46/XI5/NET35_XI46/XI5/MM10_d N_XI46/XI5/NET36_XI46/XI5/MM10_g
+ N_VDD_XI46/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI5/MM11 N_XI46/XI5/NET36_XI46/XI5/MM11_d N_XI46/XI5/NET35_XI46/XI5/MM11_g
+ N_VDD_XI46/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI6/MM2 N_XI46/XI6/NET34_XI46/XI6/MM2_d N_XI46/XI6/NET33_XI46/XI6/MM2_g
+ N_VSS_XI46/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM3 N_XI46/XI6/NET33_XI46/XI6/MM3_d N_WL<88>_XI46/XI6/MM3_g
+ N_BLN<9>_XI46/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM0 N_XI46/XI6/NET34_XI46/XI6/MM0_d N_WL<88>_XI46/XI6/MM0_g
+ N_BL<9>_XI46/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM1 N_XI46/XI6/NET33_XI46/XI6/MM1_d N_XI46/XI6/NET34_XI46/XI6/MM1_g
+ N_VSS_XI46/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM9 N_XI46/XI6/NET36_XI46/XI6/MM9_d N_WL<89>_XI46/XI6/MM9_g
+ N_BL<9>_XI46/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM6 N_XI46/XI6/NET35_XI46/XI6/MM6_d N_XI46/XI6/NET36_XI46/XI6/MM6_g
+ N_VSS_XI46/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM7 N_XI46/XI6/NET36_XI46/XI6/MM7_d N_XI46/XI6/NET35_XI46/XI6/MM7_g
+ N_VSS_XI46/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM8 N_XI46/XI6/NET35_XI46/XI6/MM8_d N_WL<89>_XI46/XI6/MM8_g
+ N_BLN<9>_XI46/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI6/MM5 N_XI46/XI6/NET34_XI46/XI6/MM5_d N_XI46/XI6/NET33_XI46/XI6/MM5_g
+ N_VDD_XI46/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI6/MM4 N_XI46/XI6/NET33_XI46/XI6/MM4_d N_XI46/XI6/NET34_XI46/XI6/MM4_g
+ N_VDD_XI46/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI6/MM10 N_XI46/XI6/NET35_XI46/XI6/MM10_d N_XI46/XI6/NET36_XI46/XI6/MM10_g
+ N_VDD_XI46/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI6/MM11 N_XI46/XI6/NET36_XI46/XI6/MM11_d N_XI46/XI6/NET35_XI46/XI6/MM11_g
+ N_VDD_XI46/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI7/MM2 N_XI46/XI7/NET34_XI46/XI7/MM2_d N_XI46/XI7/NET33_XI46/XI7/MM2_g
+ N_VSS_XI46/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM3 N_XI46/XI7/NET33_XI46/XI7/MM3_d N_WL<88>_XI46/XI7/MM3_g
+ N_BLN<8>_XI46/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM0 N_XI46/XI7/NET34_XI46/XI7/MM0_d N_WL<88>_XI46/XI7/MM0_g
+ N_BL<8>_XI46/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM1 N_XI46/XI7/NET33_XI46/XI7/MM1_d N_XI46/XI7/NET34_XI46/XI7/MM1_g
+ N_VSS_XI46/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM9 N_XI46/XI7/NET36_XI46/XI7/MM9_d N_WL<89>_XI46/XI7/MM9_g
+ N_BL<8>_XI46/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM6 N_XI46/XI7/NET35_XI46/XI7/MM6_d N_XI46/XI7/NET36_XI46/XI7/MM6_g
+ N_VSS_XI46/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM7 N_XI46/XI7/NET36_XI46/XI7/MM7_d N_XI46/XI7/NET35_XI46/XI7/MM7_g
+ N_VSS_XI46/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM8 N_XI46/XI7/NET35_XI46/XI7/MM8_d N_WL<89>_XI46/XI7/MM8_g
+ N_BLN<8>_XI46/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI7/MM5 N_XI46/XI7/NET34_XI46/XI7/MM5_d N_XI46/XI7/NET33_XI46/XI7/MM5_g
+ N_VDD_XI46/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI7/MM4 N_XI46/XI7/NET33_XI46/XI7/MM4_d N_XI46/XI7/NET34_XI46/XI7/MM4_g
+ N_VDD_XI46/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI7/MM10 N_XI46/XI7/NET35_XI46/XI7/MM10_d N_XI46/XI7/NET36_XI46/XI7/MM10_g
+ N_VDD_XI46/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI7/MM11 N_XI46/XI7/NET36_XI46/XI7/MM11_d N_XI46/XI7/NET35_XI46/XI7/MM11_g
+ N_VDD_XI46/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI8/MM2 N_XI46/XI8/NET34_XI46/XI8/MM2_d N_XI46/XI8/NET33_XI46/XI8/MM2_g
+ N_VSS_XI46/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM3 N_XI46/XI8/NET33_XI46/XI8/MM3_d N_WL<88>_XI46/XI8/MM3_g
+ N_BLN<7>_XI46/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM0 N_XI46/XI8/NET34_XI46/XI8/MM0_d N_WL<88>_XI46/XI8/MM0_g
+ N_BL<7>_XI46/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM1 N_XI46/XI8/NET33_XI46/XI8/MM1_d N_XI46/XI8/NET34_XI46/XI8/MM1_g
+ N_VSS_XI46/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM9 N_XI46/XI8/NET36_XI46/XI8/MM9_d N_WL<89>_XI46/XI8/MM9_g
+ N_BL<7>_XI46/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM6 N_XI46/XI8/NET35_XI46/XI8/MM6_d N_XI46/XI8/NET36_XI46/XI8/MM6_g
+ N_VSS_XI46/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM7 N_XI46/XI8/NET36_XI46/XI8/MM7_d N_XI46/XI8/NET35_XI46/XI8/MM7_g
+ N_VSS_XI46/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM8 N_XI46/XI8/NET35_XI46/XI8/MM8_d N_WL<89>_XI46/XI8/MM8_g
+ N_BLN<7>_XI46/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI8/MM5 N_XI46/XI8/NET34_XI46/XI8/MM5_d N_XI46/XI8/NET33_XI46/XI8/MM5_g
+ N_VDD_XI46/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI8/MM4 N_XI46/XI8/NET33_XI46/XI8/MM4_d N_XI46/XI8/NET34_XI46/XI8/MM4_g
+ N_VDD_XI46/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI8/MM10 N_XI46/XI8/NET35_XI46/XI8/MM10_d N_XI46/XI8/NET36_XI46/XI8/MM10_g
+ N_VDD_XI46/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI8/MM11 N_XI46/XI8/NET36_XI46/XI8/MM11_d N_XI46/XI8/NET35_XI46/XI8/MM11_g
+ N_VDD_XI46/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI9/MM2 N_XI46/XI9/NET34_XI46/XI9/MM2_d N_XI46/XI9/NET33_XI46/XI9/MM2_g
+ N_VSS_XI46/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM3 N_XI46/XI9/NET33_XI46/XI9/MM3_d N_WL<88>_XI46/XI9/MM3_g
+ N_BLN<6>_XI46/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM0 N_XI46/XI9/NET34_XI46/XI9/MM0_d N_WL<88>_XI46/XI9/MM0_g
+ N_BL<6>_XI46/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM1 N_XI46/XI9/NET33_XI46/XI9/MM1_d N_XI46/XI9/NET34_XI46/XI9/MM1_g
+ N_VSS_XI46/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM9 N_XI46/XI9/NET36_XI46/XI9/MM9_d N_WL<89>_XI46/XI9/MM9_g
+ N_BL<6>_XI46/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM6 N_XI46/XI9/NET35_XI46/XI9/MM6_d N_XI46/XI9/NET36_XI46/XI9/MM6_g
+ N_VSS_XI46/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM7 N_XI46/XI9/NET36_XI46/XI9/MM7_d N_XI46/XI9/NET35_XI46/XI9/MM7_g
+ N_VSS_XI46/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM8 N_XI46/XI9/NET35_XI46/XI9/MM8_d N_WL<89>_XI46/XI9/MM8_g
+ N_BLN<6>_XI46/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI9/MM5 N_XI46/XI9/NET34_XI46/XI9/MM5_d N_XI46/XI9/NET33_XI46/XI9/MM5_g
+ N_VDD_XI46/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI9/MM4 N_XI46/XI9/NET33_XI46/XI9/MM4_d N_XI46/XI9/NET34_XI46/XI9/MM4_g
+ N_VDD_XI46/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI9/MM10 N_XI46/XI9/NET35_XI46/XI9/MM10_d N_XI46/XI9/NET36_XI46/XI9/MM10_g
+ N_VDD_XI46/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI9/MM11 N_XI46/XI9/NET36_XI46/XI9/MM11_d N_XI46/XI9/NET35_XI46/XI9/MM11_g
+ N_VDD_XI46/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI10/MM2 N_XI46/XI10/NET34_XI46/XI10/MM2_d
+ N_XI46/XI10/NET33_XI46/XI10/MM2_g N_VSS_XI46/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI10/MM3 N_XI46/XI10/NET33_XI46/XI10/MM3_d N_WL<88>_XI46/XI10/MM3_g
+ N_BLN<5>_XI46/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI10/MM0 N_XI46/XI10/NET34_XI46/XI10/MM0_d N_WL<88>_XI46/XI10/MM0_g
+ N_BL<5>_XI46/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI10/MM1 N_XI46/XI10/NET33_XI46/XI10/MM1_d
+ N_XI46/XI10/NET34_XI46/XI10/MM1_g N_VSS_XI46/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI10/MM9 N_XI46/XI10/NET36_XI46/XI10/MM9_d N_WL<89>_XI46/XI10/MM9_g
+ N_BL<5>_XI46/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI10/MM6 N_XI46/XI10/NET35_XI46/XI10/MM6_d
+ N_XI46/XI10/NET36_XI46/XI10/MM6_g N_VSS_XI46/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI10/MM7 N_XI46/XI10/NET36_XI46/XI10/MM7_d
+ N_XI46/XI10/NET35_XI46/XI10/MM7_g N_VSS_XI46/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI10/MM8 N_XI46/XI10/NET35_XI46/XI10/MM8_d N_WL<89>_XI46/XI10/MM8_g
+ N_BLN<5>_XI46/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI10/MM5 N_XI46/XI10/NET34_XI46/XI10/MM5_d
+ N_XI46/XI10/NET33_XI46/XI10/MM5_g N_VDD_XI46/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI10/MM4 N_XI46/XI10/NET33_XI46/XI10/MM4_d
+ N_XI46/XI10/NET34_XI46/XI10/MM4_g N_VDD_XI46/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI10/MM10 N_XI46/XI10/NET35_XI46/XI10/MM10_d
+ N_XI46/XI10/NET36_XI46/XI10/MM10_g N_VDD_XI46/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI10/MM11 N_XI46/XI10/NET36_XI46/XI10/MM11_d
+ N_XI46/XI10/NET35_XI46/XI10/MM11_g N_VDD_XI46/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI11/MM2 N_XI46/XI11/NET34_XI46/XI11/MM2_d
+ N_XI46/XI11/NET33_XI46/XI11/MM2_g N_VSS_XI46/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI11/MM3 N_XI46/XI11/NET33_XI46/XI11/MM3_d N_WL<88>_XI46/XI11/MM3_g
+ N_BLN<4>_XI46/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI11/MM0 N_XI46/XI11/NET34_XI46/XI11/MM0_d N_WL<88>_XI46/XI11/MM0_g
+ N_BL<4>_XI46/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI11/MM1 N_XI46/XI11/NET33_XI46/XI11/MM1_d
+ N_XI46/XI11/NET34_XI46/XI11/MM1_g N_VSS_XI46/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI11/MM9 N_XI46/XI11/NET36_XI46/XI11/MM9_d N_WL<89>_XI46/XI11/MM9_g
+ N_BL<4>_XI46/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI11/MM6 N_XI46/XI11/NET35_XI46/XI11/MM6_d
+ N_XI46/XI11/NET36_XI46/XI11/MM6_g N_VSS_XI46/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI11/MM7 N_XI46/XI11/NET36_XI46/XI11/MM7_d
+ N_XI46/XI11/NET35_XI46/XI11/MM7_g N_VSS_XI46/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI11/MM8 N_XI46/XI11/NET35_XI46/XI11/MM8_d N_WL<89>_XI46/XI11/MM8_g
+ N_BLN<4>_XI46/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI11/MM5 N_XI46/XI11/NET34_XI46/XI11/MM5_d
+ N_XI46/XI11/NET33_XI46/XI11/MM5_g N_VDD_XI46/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI11/MM4 N_XI46/XI11/NET33_XI46/XI11/MM4_d
+ N_XI46/XI11/NET34_XI46/XI11/MM4_g N_VDD_XI46/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI11/MM10 N_XI46/XI11/NET35_XI46/XI11/MM10_d
+ N_XI46/XI11/NET36_XI46/XI11/MM10_g N_VDD_XI46/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI11/MM11 N_XI46/XI11/NET36_XI46/XI11/MM11_d
+ N_XI46/XI11/NET35_XI46/XI11/MM11_g N_VDD_XI46/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI12/MM2 N_XI46/XI12/NET34_XI46/XI12/MM2_d
+ N_XI46/XI12/NET33_XI46/XI12/MM2_g N_VSS_XI46/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI12/MM3 N_XI46/XI12/NET33_XI46/XI12/MM3_d N_WL<88>_XI46/XI12/MM3_g
+ N_BLN<3>_XI46/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI12/MM0 N_XI46/XI12/NET34_XI46/XI12/MM0_d N_WL<88>_XI46/XI12/MM0_g
+ N_BL<3>_XI46/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI12/MM1 N_XI46/XI12/NET33_XI46/XI12/MM1_d
+ N_XI46/XI12/NET34_XI46/XI12/MM1_g N_VSS_XI46/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI12/MM9 N_XI46/XI12/NET36_XI46/XI12/MM9_d N_WL<89>_XI46/XI12/MM9_g
+ N_BL<3>_XI46/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI12/MM6 N_XI46/XI12/NET35_XI46/XI12/MM6_d
+ N_XI46/XI12/NET36_XI46/XI12/MM6_g N_VSS_XI46/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI12/MM7 N_XI46/XI12/NET36_XI46/XI12/MM7_d
+ N_XI46/XI12/NET35_XI46/XI12/MM7_g N_VSS_XI46/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI12/MM8 N_XI46/XI12/NET35_XI46/XI12/MM8_d N_WL<89>_XI46/XI12/MM8_g
+ N_BLN<3>_XI46/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI12/MM5 N_XI46/XI12/NET34_XI46/XI12/MM5_d
+ N_XI46/XI12/NET33_XI46/XI12/MM5_g N_VDD_XI46/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI12/MM4 N_XI46/XI12/NET33_XI46/XI12/MM4_d
+ N_XI46/XI12/NET34_XI46/XI12/MM4_g N_VDD_XI46/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI12/MM10 N_XI46/XI12/NET35_XI46/XI12/MM10_d
+ N_XI46/XI12/NET36_XI46/XI12/MM10_g N_VDD_XI46/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI12/MM11 N_XI46/XI12/NET36_XI46/XI12/MM11_d
+ N_XI46/XI12/NET35_XI46/XI12/MM11_g N_VDD_XI46/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI13/MM2 N_XI46/XI13/NET34_XI46/XI13/MM2_d
+ N_XI46/XI13/NET33_XI46/XI13/MM2_g N_VSS_XI46/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI13/MM3 N_XI46/XI13/NET33_XI46/XI13/MM3_d N_WL<88>_XI46/XI13/MM3_g
+ N_BLN<2>_XI46/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI13/MM0 N_XI46/XI13/NET34_XI46/XI13/MM0_d N_WL<88>_XI46/XI13/MM0_g
+ N_BL<2>_XI46/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI13/MM1 N_XI46/XI13/NET33_XI46/XI13/MM1_d
+ N_XI46/XI13/NET34_XI46/XI13/MM1_g N_VSS_XI46/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI13/MM9 N_XI46/XI13/NET36_XI46/XI13/MM9_d N_WL<89>_XI46/XI13/MM9_g
+ N_BL<2>_XI46/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI13/MM6 N_XI46/XI13/NET35_XI46/XI13/MM6_d
+ N_XI46/XI13/NET36_XI46/XI13/MM6_g N_VSS_XI46/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI13/MM7 N_XI46/XI13/NET36_XI46/XI13/MM7_d
+ N_XI46/XI13/NET35_XI46/XI13/MM7_g N_VSS_XI46/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI13/MM8 N_XI46/XI13/NET35_XI46/XI13/MM8_d N_WL<89>_XI46/XI13/MM8_g
+ N_BLN<2>_XI46/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI13/MM5 N_XI46/XI13/NET34_XI46/XI13/MM5_d
+ N_XI46/XI13/NET33_XI46/XI13/MM5_g N_VDD_XI46/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI13/MM4 N_XI46/XI13/NET33_XI46/XI13/MM4_d
+ N_XI46/XI13/NET34_XI46/XI13/MM4_g N_VDD_XI46/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI13/MM10 N_XI46/XI13/NET35_XI46/XI13/MM10_d
+ N_XI46/XI13/NET36_XI46/XI13/MM10_g N_VDD_XI46/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI13/MM11 N_XI46/XI13/NET36_XI46/XI13/MM11_d
+ N_XI46/XI13/NET35_XI46/XI13/MM11_g N_VDD_XI46/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI14/MM2 N_XI46/XI14/NET34_XI46/XI14/MM2_d
+ N_XI46/XI14/NET33_XI46/XI14/MM2_g N_VSS_XI46/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI14/MM3 N_XI46/XI14/NET33_XI46/XI14/MM3_d N_WL<88>_XI46/XI14/MM3_g
+ N_BLN<1>_XI46/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI14/MM0 N_XI46/XI14/NET34_XI46/XI14/MM0_d N_WL<88>_XI46/XI14/MM0_g
+ N_BL<1>_XI46/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI14/MM1 N_XI46/XI14/NET33_XI46/XI14/MM1_d
+ N_XI46/XI14/NET34_XI46/XI14/MM1_g N_VSS_XI46/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI14/MM9 N_XI46/XI14/NET36_XI46/XI14/MM9_d N_WL<89>_XI46/XI14/MM9_g
+ N_BL<1>_XI46/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI14/MM6 N_XI46/XI14/NET35_XI46/XI14/MM6_d
+ N_XI46/XI14/NET36_XI46/XI14/MM6_g N_VSS_XI46/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI14/MM7 N_XI46/XI14/NET36_XI46/XI14/MM7_d
+ N_XI46/XI14/NET35_XI46/XI14/MM7_g N_VSS_XI46/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI14/MM8 N_XI46/XI14/NET35_XI46/XI14/MM8_d N_WL<89>_XI46/XI14/MM8_g
+ N_BLN<1>_XI46/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI14/MM5 N_XI46/XI14/NET34_XI46/XI14/MM5_d
+ N_XI46/XI14/NET33_XI46/XI14/MM5_g N_VDD_XI46/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI14/MM4 N_XI46/XI14/NET33_XI46/XI14/MM4_d
+ N_XI46/XI14/NET34_XI46/XI14/MM4_g N_VDD_XI46/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI14/MM10 N_XI46/XI14/NET35_XI46/XI14/MM10_d
+ N_XI46/XI14/NET36_XI46/XI14/MM10_g N_VDD_XI46/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI14/MM11 N_XI46/XI14/NET36_XI46/XI14/MM11_d
+ N_XI46/XI14/NET35_XI46/XI14/MM11_g N_VDD_XI46/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI15/MM2 N_XI46/XI15/NET34_XI46/XI15/MM2_d
+ N_XI46/XI15/NET33_XI46/XI15/MM2_g N_VSS_XI46/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI15/MM3 N_XI46/XI15/NET33_XI46/XI15/MM3_d N_WL<88>_XI46/XI15/MM3_g
+ N_BLN<0>_XI46/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI15/MM0 N_XI46/XI15/NET34_XI46/XI15/MM0_d N_WL<88>_XI46/XI15/MM0_g
+ N_BL<0>_XI46/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI15/MM1 N_XI46/XI15/NET33_XI46/XI15/MM1_d
+ N_XI46/XI15/NET34_XI46/XI15/MM1_g N_VSS_XI46/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI15/MM9 N_XI46/XI15/NET36_XI46/XI15/MM9_d N_WL<89>_XI46/XI15/MM9_g
+ N_BL<0>_XI46/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI15/MM6 N_XI46/XI15/NET35_XI46/XI15/MM6_d
+ N_XI46/XI15/NET36_XI46/XI15/MM6_g N_VSS_XI46/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI15/MM7 N_XI46/XI15/NET36_XI46/XI15/MM7_d
+ N_XI46/XI15/NET35_XI46/XI15/MM7_g N_VSS_XI46/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI46/XI15/MM8 N_XI46/XI15/NET35_XI46/XI15/MM8_d N_WL<89>_XI46/XI15/MM8_g
+ N_BLN<0>_XI46/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI46/XI15/MM5 N_XI46/XI15/NET34_XI46/XI15/MM5_d
+ N_XI46/XI15/NET33_XI46/XI15/MM5_g N_VDD_XI46/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI15/MM4 N_XI46/XI15/NET33_XI46/XI15/MM4_d
+ N_XI46/XI15/NET34_XI46/XI15/MM4_g N_VDD_XI46/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI15/MM10 N_XI46/XI15/NET35_XI46/XI15/MM10_d
+ N_XI46/XI15/NET36_XI46/XI15/MM10_g N_VDD_XI46/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI46/XI15/MM11 N_XI46/XI15/NET36_XI46/XI15/MM11_d
+ N_XI46/XI15/NET35_XI46/XI15/MM11_g N_VDD_XI46/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI0/MM2 N_XI47/XI0/NET34_XI47/XI0/MM2_d N_XI47/XI0/NET33_XI47/XI0/MM2_g
+ N_VSS_XI47/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI0/MM3 N_XI47/XI0/NET33_XI47/XI0/MM3_d N_WL<90>_XI47/XI0/MM3_g
+ N_BLN<15>_XI47/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI0/MM0 N_XI47/XI0/NET34_XI47/XI0/MM0_d N_WL<90>_XI47/XI0/MM0_g
+ N_BL<15>_XI47/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI0/MM1 N_XI47/XI0/NET33_XI47/XI0/MM1_d N_XI47/XI0/NET34_XI47/XI0/MM1_g
+ N_VSS_XI47/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI0/MM9 N_XI47/XI0/NET36_XI47/XI0/MM9_d N_WL<91>_XI47/XI0/MM9_g
+ N_BL<15>_XI47/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI0/MM6 N_XI47/XI0/NET35_XI47/XI0/MM6_d N_XI47/XI0/NET36_XI47/XI0/MM6_g
+ N_VSS_XI47/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI0/MM7 N_XI47/XI0/NET36_XI47/XI0/MM7_d N_XI47/XI0/NET35_XI47/XI0/MM7_g
+ N_VSS_XI47/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI0/MM8 N_XI47/XI0/NET35_XI47/XI0/MM8_d N_WL<91>_XI47/XI0/MM8_g
+ N_BLN<15>_XI47/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI0/MM5 N_XI47/XI0/NET34_XI47/XI0/MM5_d N_XI47/XI0/NET33_XI47/XI0/MM5_g
+ N_VDD_XI47/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI0/MM4 N_XI47/XI0/NET33_XI47/XI0/MM4_d N_XI47/XI0/NET34_XI47/XI0/MM4_g
+ N_VDD_XI47/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI0/MM10 N_XI47/XI0/NET35_XI47/XI0/MM10_d N_XI47/XI0/NET36_XI47/XI0/MM10_g
+ N_VDD_XI47/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI0/MM11 N_XI47/XI0/NET36_XI47/XI0/MM11_d N_XI47/XI0/NET35_XI47/XI0/MM11_g
+ N_VDD_XI47/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI1/MM2 N_XI47/XI1/NET34_XI47/XI1/MM2_d N_XI47/XI1/NET33_XI47/XI1/MM2_g
+ N_VSS_XI47/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI1/MM3 N_XI47/XI1/NET33_XI47/XI1/MM3_d N_WL<90>_XI47/XI1/MM3_g
+ N_BLN<14>_XI47/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI1/MM0 N_XI47/XI1/NET34_XI47/XI1/MM0_d N_WL<90>_XI47/XI1/MM0_g
+ N_BL<14>_XI47/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI1/MM1 N_XI47/XI1/NET33_XI47/XI1/MM1_d N_XI47/XI1/NET34_XI47/XI1/MM1_g
+ N_VSS_XI47/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI1/MM9 N_XI47/XI1/NET36_XI47/XI1/MM9_d N_WL<91>_XI47/XI1/MM9_g
+ N_BL<14>_XI47/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI1/MM6 N_XI47/XI1/NET35_XI47/XI1/MM6_d N_XI47/XI1/NET36_XI47/XI1/MM6_g
+ N_VSS_XI47/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI1/MM7 N_XI47/XI1/NET36_XI47/XI1/MM7_d N_XI47/XI1/NET35_XI47/XI1/MM7_g
+ N_VSS_XI47/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI1/MM8 N_XI47/XI1/NET35_XI47/XI1/MM8_d N_WL<91>_XI47/XI1/MM8_g
+ N_BLN<14>_XI47/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI1/MM5 N_XI47/XI1/NET34_XI47/XI1/MM5_d N_XI47/XI1/NET33_XI47/XI1/MM5_g
+ N_VDD_XI47/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI1/MM4 N_XI47/XI1/NET33_XI47/XI1/MM4_d N_XI47/XI1/NET34_XI47/XI1/MM4_g
+ N_VDD_XI47/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI1/MM10 N_XI47/XI1/NET35_XI47/XI1/MM10_d N_XI47/XI1/NET36_XI47/XI1/MM10_g
+ N_VDD_XI47/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI1/MM11 N_XI47/XI1/NET36_XI47/XI1/MM11_d N_XI47/XI1/NET35_XI47/XI1/MM11_g
+ N_VDD_XI47/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI2/MM2 N_XI47/XI2/NET34_XI47/XI2/MM2_d N_XI47/XI2/NET33_XI47/XI2/MM2_g
+ N_VSS_XI47/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI2/MM3 N_XI47/XI2/NET33_XI47/XI2/MM3_d N_WL<90>_XI47/XI2/MM3_g
+ N_BLN<13>_XI47/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI2/MM0 N_XI47/XI2/NET34_XI47/XI2/MM0_d N_WL<90>_XI47/XI2/MM0_g
+ N_BL<13>_XI47/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI2/MM1 N_XI47/XI2/NET33_XI47/XI2/MM1_d N_XI47/XI2/NET34_XI47/XI2/MM1_g
+ N_VSS_XI47/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI2/MM9 N_XI47/XI2/NET36_XI47/XI2/MM9_d N_WL<91>_XI47/XI2/MM9_g
+ N_BL<13>_XI47/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI2/MM6 N_XI47/XI2/NET35_XI47/XI2/MM6_d N_XI47/XI2/NET36_XI47/XI2/MM6_g
+ N_VSS_XI47/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI2/MM7 N_XI47/XI2/NET36_XI47/XI2/MM7_d N_XI47/XI2/NET35_XI47/XI2/MM7_g
+ N_VSS_XI47/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI2/MM8 N_XI47/XI2/NET35_XI47/XI2/MM8_d N_WL<91>_XI47/XI2/MM8_g
+ N_BLN<13>_XI47/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI2/MM5 N_XI47/XI2/NET34_XI47/XI2/MM5_d N_XI47/XI2/NET33_XI47/XI2/MM5_g
+ N_VDD_XI47/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI2/MM4 N_XI47/XI2/NET33_XI47/XI2/MM4_d N_XI47/XI2/NET34_XI47/XI2/MM4_g
+ N_VDD_XI47/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI2/MM10 N_XI47/XI2/NET35_XI47/XI2/MM10_d N_XI47/XI2/NET36_XI47/XI2/MM10_g
+ N_VDD_XI47/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI2/MM11 N_XI47/XI2/NET36_XI47/XI2/MM11_d N_XI47/XI2/NET35_XI47/XI2/MM11_g
+ N_VDD_XI47/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI3/MM2 N_XI47/XI3/NET34_XI47/XI3/MM2_d N_XI47/XI3/NET33_XI47/XI3/MM2_g
+ N_VSS_XI47/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI3/MM3 N_XI47/XI3/NET33_XI47/XI3/MM3_d N_WL<90>_XI47/XI3/MM3_g
+ N_BLN<12>_XI47/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI3/MM0 N_XI47/XI3/NET34_XI47/XI3/MM0_d N_WL<90>_XI47/XI3/MM0_g
+ N_BL<12>_XI47/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI3/MM1 N_XI47/XI3/NET33_XI47/XI3/MM1_d N_XI47/XI3/NET34_XI47/XI3/MM1_g
+ N_VSS_XI47/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI3/MM9 N_XI47/XI3/NET36_XI47/XI3/MM9_d N_WL<91>_XI47/XI3/MM9_g
+ N_BL<12>_XI47/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI3/MM6 N_XI47/XI3/NET35_XI47/XI3/MM6_d N_XI47/XI3/NET36_XI47/XI3/MM6_g
+ N_VSS_XI47/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI3/MM7 N_XI47/XI3/NET36_XI47/XI3/MM7_d N_XI47/XI3/NET35_XI47/XI3/MM7_g
+ N_VSS_XI47/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI3/MM8 N_XI47/XI3/NET35_XI47/XI3/MM8_d N_WL<91>_XI47/XI3/MM8_g
+ N_BLN<12>_XI47/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI3/MM5 N_XI47/XI3/NET34_XI47/XI3/MM5_d N_XI47/XI3/NET33_XI47/XI3/MM5_g
+ N_VDD_XI47/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI3/MM4 N_XI47/XI3/NET33_XI47/XI3/MM4_d N_XI47/XI3/NET34_XI47/XI3/MM4_g
+ N_VDD_XI47/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI3/MM10 N_XI47/XI3/NET35_XI47/XI3/MM10_d N_XI47/XI3/NET36_XI47/XI3/MM10_g
+ N_VDD_XI47/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI3/MM11 N_XI47/XI3/NET36_XI47/XI3/MM11_d N_XI47/XI3/NET35_XI47/XI3/MM11_g
+ N_VDD_XI47/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI4/MM2 N_XI47/XI4/NET34_XI47/XI4/MM2_d N_XI47/XI4/NET33_XI47/XI4/MM2_g
+ N_VSS_XI47/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI4/MM3 N_XI47/XI4/NET33_XI47/XI4/MM3_d N_WL<90>_XI47/XI4/MM3_g
+ N_BLN<11>_XI47/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI4/MM0 N_XI47/XI4/NET34_XI47/XI4/MM0_d N_WL<90>_XI47/XI4/MM0_g
+ N_BL<11>_XI47/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI4/MM1 N_XI47/XI4/NET33_XI47/XI4/MM1_d N_XI47/XI4/NET34_XI47/XI4/MM1_g
+ N_VSS_XI47/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI4/MM9 N_XI47/XI4/NET36_XI47/XI4/MM9_d N_WL<91>_XI47/XI4/MM9_g
+ N_BL<11>_XI47/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI4/MM6 N_XI47/XI4/NET35_XI47/XI4/MM6_d N_XI47/XI4/NET36_XI47/XI4/MM6_g
+ N_VSS_XI47/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI4/MM7 N_XI47/XI4/NET36_XI47/XI4/MM7_d N_XI47/XI4/NET35_XI47/XI4/MM7_g
+ N_VSS_XI47/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI4/MM8 N_XI47/XI4/NET35_XI47/XI4/MM8_d N_WL<91>_XI47/XI4/MM8_g
+ N_BLN<11>_XI47/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI4/MM5 N_XI47/XI4/NET34_XI47/XI4/MM5_d N_XI47/XI4/NET33_XI47/XI4/MM5_g
+ N_VDD_XI47/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI4/MM4 N_XI47/XI4/NET33_XI47/XI4/MM4_d N_XI47/XI4/NET34_XI47/XI4/MM4_g
+ N_VDD_XI47/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI4/MM10 N_XI47/XI4/NET35_XI47/XI4/MM10_d N_XI47/XI4/NET36_XI47/XI4/MM10_g
+ N_VDD_XI47/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI4/MM11 N_XI47/XI4/NET36_XI47/XI4/MM11_d N_XI47/XI4/NET35_XI47/XI4/MM11_g
+ N_VDD_XI47/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI5/MM2 N_XI47/XI5/NET34_XI47/XI5/MM2_d N_XI47/XI5/NET33_XI47/XI5/MM2_g
+ N_VSS_XI47/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI5/MM3 N_XI47/XI5/NET33_XI47/XI5/MM3_d N_WL<90>_XI47/XI5/MM3_g
+ N_BLN<10>_XI47/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI5/MM0 N_XI47/XI5/NET34_XI47/XI5/MM0_d N_WL<90>_XI47/XI5/MM0_g
+ N_BL<10>_XI47/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI5/MM1 N_XI47/XI5/NET33_XI47/XI5/MM1_d N_XI47/XI5/NET34_XI47/XI5/MM1_g
+ N_VSS_XI47/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI5/MM9 N_XI47/XI5/NET36_XI47/XI5/MM9_d N_WL<91>_XI47/XI5/MM9_g
+ N_BL<10>_XI47/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI5/MM6 N_XI47/XI5/NET35_XI47/XI5/MM6_d N_XI47/XI5/NET36_XI47/XI5/MM6_g
+ N_VSS_XI47/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI5/MM7 N_XI47/XI5/NET36_XI47/XI5/MM7_d N_XI47/XI5/NET35_XI47/XI5/MM7_g
+ N_VSS_XI47/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI5/MM8 N_XI47/XI5/NET35_XI47/XI5/MM8_d N_WL<91>_XI47/XI5/MM8_g
+ N_BLN<10>_XI47/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI5/MM5 N_XI47/XI5/NET34_XI47/XI5/MM5_d N_XI47/XI5/NET33_XI47/XI5/MM5_g
+ N_VDD_XI47/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI5/MM4 N_XI47/XI5/NET33_XI47/XI5/MM4_d N_XI47/XI5/NET34_XI47/XI5/MM4_g
+ N_VDD_XI47/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI5/MM10 N_XI47/XI5/NET35_XI47/XI5/MM10_d N_XI47/XI5/NET36_XI47/XI5/MM10_g
+ N_VDD_XI47/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI5/MM11 N_XI47/XI5/NET36_XI47/XI5/MM11_d N_XI47/XI5/NET35_XI47/XI5/MM11_g
+ N_VDD_XI47/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI6/MM2 N_XI47/XI6/NET34_XI47/XI6/MM2_d N_XI47/XI6/NET33_XI47/XI6/MM2_g
+ N_VSS_XI47/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM3 N_XI47/XI6/NET33_XI47/XI6/MM3_d N_WL<90>_XI47/XI6/MM3_g
+ N_BLN<9>_XI47/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM0 N_XI47/XI6/NET34_XI47/XI6/MM0_d N_WL<90>_XI47/XI6/MM0_g
+ N_BL<9>_XI47/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM1 N_XI47/XI6/NET33_XI47/XI6/MM1_d N_XI47/XI6/NET34_XI47/XI6/MM1_g
+ N_VSS_XI47/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM9 N_XI47/XI6/NET36_XI47/XI6/MM9_d N_WL<91>_XI47/XI6/MM9_g
+ N_BL<9>_XI47/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM6 N_XI47/XI6/NET35_XI47/XI6/MM6_d N_XI47/XI6/NET36_XI47/XI6/MM6_g
+ N_VSS_XI47/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM7 N_XI47/XI6/NET36_XI47/XI6/MM7_d N_XI47/XI6/NET35_XI47/XI6/MM7_g
+ N_VSS_XI47/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM8 N_XI47/XI6/NET35_XI47/XI6/MM8_d N_WL<91>_XI47/XI6/MM8_g
+ N_BLN<9>_XI47/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI6/MM5 N_XI47/XI6/NET34_XI47/XI6/MM5_d N_XI47/XI6/NET33_XI47/XI6/MM5_g
+ N_VDD_XI47/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI6/MM4 N_XI47/XI6/NET33_XI47/XI6/MM4_d N_XI47/XI6/NET34_XI47/XI6/MM4_g
+ N_VDD_XI47/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI6/MM10 N_XI47/XI6/NET35_XI47/XI6/MM10_d N_XI47/XI6/NET36_XI47/XI6/MM10_g
+ N_VDD_XI47/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI6/MM11 N_XI47/XI6/NET36_XI47/XI6/MM11_d N_XI47/XI6/NET35_XI47/XI6/MM11_g
+ N_VDD_XI47/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI7/MM2 N_XI47/XI7/NET34_XI47/XI7/MM2_d N_XI47/XI7/NET33_XI47/XI7/MM2_g
+ N_VSS_XI47/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM3 N_XI47/XI7/NET33_XI47/XI7/MM3_d N_WL<90>_XI47/XI7/MM3_g
+ N_BLN<8>_XI47/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM0 N_XI47/XI7/NET34_XI47/XI7/MM0_d N_WL<90>_XI47/XI7/MM0_g
+ N_BL<8>_XI47/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM1 N_XI47/XI7/NET33_XI47/XI7/MM1_d N_XI47/XI7/NET34_XI47/XI7/MM1_g
+ N_VSS_XI47/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM9 N_XI47/XI7/NET36_XI47/XI7/MM9_d N_WL<91>_XI47/XI7/MM9_g
+ N_BL<8>_XI47/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM6 N_XI47/XI7/NET35_XI47/XI7/MM6_d N_XI47/XI7/NET36_XI47/XI7/MM6_g
+ N_VSS_XI47/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM7 N_XI47/XI7/NET36_XI47/XI7/MM7_d N_XI47/XI7/NET35_XI47/XI7/MM7_g
+ N_VSS_XI47/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM8 N_XI47/XI7/NET35_XI47/XI7/MM8_d N_WL<91>_XI47/XI7/MM8_g
+ N_BLN<8>_XI47/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI7/MM5 N_XI47/XI7/NET34_XI47/XI7/MM5_d N_XI47/XI7/NET33_XI47/XI7/MM5_g
+ N_VDD_XI47/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI7/MM4 N_XI47/XI7/NET33_XI47/XI7/MM4_d N_XI47/XI7/NET34_XI47/XI7/MM4_g
+ N_VDD_XI47/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI7/MM10 N_XI47/XI7/NET35_XI47/XI7/MM10_d N_XI47/XI7/NET36_XI47/XI7/MM10_g
+ N_VDD_XI47/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI7/MM11 N_XI47/XI7/NET36_XI47/XI7/MM11_d N_XI47/XI7/NET35_XI47/XI7/MM11_g
+ N_VDD_XI47/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI8/MM2 N_XI47/XI8/NET34_XI47/XI8/MM2_d N_XI47/XI8/NET33_XI47/XI8/MM2_g
+ N_VSS_XI47/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM3 N_XI47/XI8/NET33_XI47/XI8/MM3_d N_WL<90>_XI47/XI8/MM3_g
+ N_BLN<7>_XI47/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM0 N_XI47/XI8/NET34_XI47/XI8/MM0_d N_WL<90>_XI47/XI8/MM0_g
+ N_BL<7>_XI47/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM1 N_XI47/XI8/NET33_XI47/XI8/MM1_d N_XI47/XI8/NET34_XI47/XI8/MM1_g
+ N_VSS_XI47/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM9 N_XI47/XI8/NET36_XI47/XI8/MM9_d N_WL<91>_XI47/XI8/MM9_g
+ N_BL<7>_XI47/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM6 N_XI47/XI8/NET35_XI47/XI8/MM6_d N_XI47/XI8/NET36_XI47/XI8/MM6_g
+ N_VSS_XI47/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM7 N_XI47/XI8/NET36_XI47/XI8/MM7_d N_XI47/XI8/NET35_XI47/XI8/MM7_g
+ N_VSS_XI47/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM8 N_XI47/XI8/NET35_XI47/XI8/MM8_d N_WL<91>_XI47/XI8/MM8_g
+ N_BLN<7>_XI47/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI8/MM5 N_XI47/XI8/NET34_XI47/XI8/MM5_d N_XI47/XI8/NET33_XI47/XI8/MM5_g
+ N_VDD_XI47/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI8/MM4 N_XI47/XI8/NET33_XI47/XI8/MM4_d N_XI47/XI8/NET34_XI47/XI8/MM4_g
+ N_VDD_XI47/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI8/MM10 N_XI47/XI8/NET35_XI47/XI8/MM10_d N_XI47/XI8/NET36_XI47/XI8/MM10_g
+ N_VDD_XI47/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI8/MM11 N_XI47/XI8/NET36_XI47/XI8/MM11_d N_XI47/XI8/NET35_XI47/XI8/MM11_g
+ N_VDD_XI47/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI9/MM2 N_XI47/XI9/NET34_XI47/XI9/MM2_d N_XI47/XI9/NET33_XI47/XI9/MM2_g
+ N_VSS_XI47/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM3 N_XI47/XI9/NET33_XI47/XI9/MM3_d N_WL<90>_XI47/XI9/MM3_g
+ N_BLN<6>_XI47/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM0 N_XI47/XI9/NET34_XI47/XI9/MM0_d N_WL<90>_XI47/XI9/MM0_g
+ N_BL<6>_XI47/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM1 N_XI47/XI9/NET33_XI47/XI9/MM1_d N_XI47/XI9/NET34_XI47/XI9/MM1_g
+ N_VSS_XI47/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM9 N_XI47/XI9/NET36_XI47/XI9/MM9_d N_WL<91>_XI47/XI9/MM9_g
+ N_BL<6>_XI47/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM6 N_XI47/XI9/NET35_XI47/XI9/MM6_d N_XI47/XI9/NET36_XI47/XI9/MM6_g
+ N_VSS_XI47/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM7 N_XI47/XI9/NET36_XI47/XI9/MM7_d N_XI47/XI9/NET35_XI47/XI9/MM7_g
+ N_VSS_XI47/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM8 N_XI47/XI9/NET35_XI47/XI9/MM8_d N_WL<91>_XI47/XI9/MM8_g
+ N_BLN<6>_XI47/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI9/MM5 N_XI47/XI9/NET34_XI47/XI9/MM5_d N_XI47/XI9/NET33_XI47/XI9/MM5_g
+ N_VDD_XI47/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI9/MM4 N_XI47/XI9/NET33_XI47/XI9/MM4_d N_XI47/XI9/NET34_XI47/XI9/MM4_g
+ N_VDD_XI47/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI9/MM10 N_XI47/XI9/NET35_XI47/XI9/MM10_d N_XI47/XI9/NET36_XI47/XI9/MM10_g
+ N_VDD_XI47/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI9/MM11 N_XI47/XI9/NET36_XI47/XI9/MM11_d N_XI47/XI9/NET35_XI47/XI9/MM11_g
+ N_VDD_XI47/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI10/MM2 N_XI47/XI10/NET34_XI47/XI10/MM2_d
+ N_XI47/XI10/NET33_XI47/XI10/MM2_g N_VSS_XI47/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI10/MM3 N_XI47/XI10/NET33_XI47/XI10/MM3_d N_WL<90>_XI47/XI10/MM3_g
+ N_BLN<5>_XI47/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI10/MM0 N_XI47/XI10/NET34_XI47/XI10/MM0_d N_WL<90>_XI47/XI10/MM0_g
+ N_BL<5>_XI47/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI10/MM1 N_XI47/XI10/NET33_XI47/XI10/MM1_d
+ N_XI47/XI10/NET34_XI47/XI10/MM1_g N_VSS_XI47/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI10/MM9 N_XI47/XI10/NET36_XI47/XI10/MM9_d N_WL<91>_XI47/XI10/MM9_g
+ N_BL<5>_XI47/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI10/MM6 N_XI47/XI10/NET35_XI47/XI10/MM6_d
+ N_XI47/XI10/NET36_XI47/XI10/MM6_g N_VSS_XI47/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI10/MM7 N_XI47/XI10/NET36_XI47/XI10/MM7_d
+ N_XI47/XI10/NET35_XI47/XI10/MM7_g N_VSS_XI47/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI10/MM8 N_XI47/XI10/NET35_XI47/XI10/MM8_d N_WL<91>_XI47/XI10/MM8_g
+ N_BLN<5>_XI47/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI10/MM5 N_XI47/XI10/NET34_XI47/XI10/MM5_d
+ N_XI47/XI10/NET33_XI47/XI10/MM5_g N_VDD_XI47/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI10/MM4 N_XI47/XI10/NET33_XI47/XI10/MM4_d
+ N_XI47/XI10/NET34_XI47/XI10/MM4_g N_VDD_XI47/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI10/MM10 N_XI47/XI10/NET35_XI47/XI10/MM10_d
+ N_XI47/XI10/NET36_XI47/XI10/MM10_g N_VDD_XI47/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI10/MM11 N_XI47/XI10/NET36_XI47/XI10/MM11_d
+ N_XI47/XI10/NET35_XI47/XI10/MM11_g N_VDD_XI47/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI11/MM2 N_XI47/XI11/NET34_XI47/XI11/MM2_d
+ N_XI47/XI11/NET33_XI47/XI11/MM2_g N_VSS_XI47/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI11/MM3 N_XI47/XI11/NET33_XI47/XI11/MM3_d N_WL<90>_XI47/XI11/MM3_g
+ N_BLN<4>_XI47/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI11/MM0 N_XI47/XI11/NET34_XI47/XI11/MM0_d N_WL<90>_XI47/XI11/MM0_g
+ N_BL<4>_XI47/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI11/MM1 N_XI47/XI11/NET33_XI47/XI11/MM1_d
+ N_XI47/XI11/NET34_XI47/XI11/MM1_g N_VSS_XI47/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI11/MM9 N_XI47/XI11/NET36_XI47/XI11/MM9_d N_WL<91>_XI47/XI11/MM9_g
+ N_BL<4>_XI47/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI11/MM6 N_XI47/XI11/NET35_XI47/XI11/MM6_d
+ N_XI47/XI11/NET36_XI47/XI11/MM6_g N_VSS_XI47/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI11/MM7 N_XI47/XI11/NET36_XI47/XI11/MM7_d
+ N_XI47/XI11/NET35_XI47/XI11/MM7_g N_VSS_XI47/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI11/MM8 N_XI47/XI11/NET35_XI47/XI11/MM8_d N_WL<91>_XI47/XI11/MM8_g
+ N_BLN<4>_XI47/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI11/MM5 N_XI47/XI11/NET34_XI47/XI11/MM5_d
+ N_XI47/XI11/NET33_XI47/XI11/MM5_g N_VDD_XI47/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI11/MM4 N_XI47/XI11/NET33_XI47/XI11/MM4_d
+ N_XI47/XI11/NET34_XI47/XI11/MM4_g N_VDD_XI47/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI11/MM10 N_XI47/XI11/NET35_XI47/XI11/MM10_d
+ N_XI47/XI11/NET36_XI47/XI11/MM10_g N_VDD_XI47/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI11/MM11 N_XI47/XI11/NET36_XI47/XI11/MM11_d
+ N_XI47/XI11/NET35_XI47/XI11/MM11_g N_VDD_XI47/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI12/MM2 N_XI47/XI12/NET34_XI47/XI12/MM2_d
+ N_XI47/XI12/NET33_XI47/XI12/MM2_g N_VSS_XI47/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI12/MM3 N_XI47/XI12/NET33_XI47/XI12/MM3_d N_WL<90>_XI47/XI12/MM3_g
+ N_BLN<3>_XI47/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI12/MM0 N_XI47/XI12/NET34_XI47/XI12/MM0_d N_WL<90>_XI47/XI12/MM0_g
+ N_BL<3>_XI47/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI12/MM1 N_XI47/XI12/NET33_XI47/XI12/MM1_d
+ N_XI47/XI12/NET34_XI47/XI12/MM1_g N_VSS_XI47/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI12/MM9 N_XI47/XI12/NET36_XI47/XI12/MM9_d N_WL<91>_XI47/XI12/MM9_g
+ N_BL<3>_XI47/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI12/MM6 N_XI47/XI12/NET35_XI47/XI12/MM6_d
+ N_XI47/XI12/NET36_XI47/XI12/MM6_g N_VSS_XI47/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI12/MM7 N_XI47/XI12/NET36_XI47/XI12/MM7_d
+ N_XI47/XI12/NET35_XI47/XI12/MM7_g N_VSS_XI47/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI12/MM8 N_XI47/XI12/NET35_XI47/XI12/MM8_d N_WL<91>_XI47/XI12/MM8_g
+ N_BLN<3>_XI47/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI12/MM5 N_XI47/XI12/NET34_XI47/XI12/MM5_d
+ N_XI47/XI12/NET33_XI47/XI12/MM5_g N_VDD_XI47/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI12/MM4 N_XI47/XI12/NET33_XI47/XI12/MM4_d
+ N_XI47/XI12/NET34_XI47/XI12/MM4_g N_VDD_XI47/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI12/MM10 N_XI47/XI12/NET35_XI47/XI12/MM10_d
+ N_XI47/XI12/NET36_XI47/XI12/MM10_g N_VDD_XI47/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI12/MM11 N_XI47/XI12/NET36_XI47/XI12/MM11_d
+ N_XI47/XI12/NET35_XI47/XI12/MM11_g N_VDD_XI47/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI13/MM2 N_XI47/XI13/NET34_XI47/XI13/MM2_d
+ N_XI47/XI13/NET33_XI47/XI13/MM2_g N_VSS_XI47/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI13/MM3 N_XI47/XI13/NET33_XI47/XI13/MM3_d N_WL<90>_XI47/XI13/MM3_g
+ N_BLN<2>_XI47/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI13/MM0 N_XI47/XI13/NET34_XI47/XI13/MM0_d N_WL<90>_XI47/XI13/MM0_g
+ N_BL<2>_XI47/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI13/MM1 N_XI47/XI13/NET33_XI47/XI13/MM1_d
+ N_XI47/XI13/NET34_XI47/XI13/MM1_g N_VSS_XI47/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI13/MM9 N_XI47/XI13/NET36_XI47/XI13/MM9_d N_WL<91>_XI47/XI13/MM9_g
+ N_BL<2>_XI47/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI13/MM6 N_XI47/XI13/NET35_XI47/XI13/MM6_d
+ N_XI47/XI13/NET36_XI47/XI13/MM6_g N_VSS_XI47/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI13/MM7 N_XI47/XI13/NET36_XI47/XI13/MM7_d
+ N_XI47/XI13/NET35_XI47/XI13/MM7_g N_VSS_XI47/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI13/MM8 N_XI47/XI13/NET35_XI47/XI13/MM8_d N_WL<91>_XI47/XI13/MM8_g
+ N_BLN<2>_XI47/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI13/MM5 N_XI47/XI13/NET34_XI47/XI13/MM5_d
+ N_XI47/XI13/NET33_XI47/XI13/MM5_g N_VDD_XI47/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI13/MM4 N_XI47/XI13/NET33_XI47/XI13/MM4_d
+ N_XI47/XI13/NET34_XI47/XI13/MM4_g N_VDD_XI47/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI13/MM10 N_XI47/XI13/NET35_XI47/XI13/MM10_d
+ N_XI47/XI13/NET36_XI47/XI13/MM10_g N_VDD_XI47/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI13/MM11 N_XI47/XI13/NET36_XI47/XI13/MM11_d
+ N_XI47/XI13/NET35_XI47/XI13/MM11_g N_VDD_XI47/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI14/MM2 N_XI47/XI14/NET34_XI47/XI14/MM2_d
+ N_XI47/XI14/NET33_XI47/XI14/MM2_g N_VSS_XI47/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI14/MM3 N_XI47/XI14/NET33_XI47/XI14/MM3_d N_WL<90>_XI47/XI14/MM3_g
+ N_BLN<1>_XI47/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI14/MM0 N_XI47/XI14/NET34_XI47/XI14/MM0_d N_WL<90>_XI47/XI14/MM0_g
+ N_BL<1>_XI47/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI14/MM1 N_XI47/XI14/NET33_XI47/XI14/MM1_d
+ N_XI47/XI14/NET34_XI47/XI14/MM1_g N_VSS_XI47/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI14/MM9 N_XI47/XI14/NET36_XI47/XI14/MM9_d N_WL<91>_XI47/XI14/MM9_g
+ N_BL<1>_XI47/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI14/MM6 N_XI47/XI14/NET35_XI47/XI14/MM6_d
+ N_XI47/XI14/NET36_XI47/XI14/MM6_g N_VSS_XI47/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI14/MM7 N_XI47/XI14/NET36_XI47/XI14/MM7_d
+ N_XI47/XI14/NET35_XI47/XI14/MM7_g N_VSS_XI47/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI14/MM8 N_XI47/XI14/NET35_XI47/XI14/MM8_d N_WL<91>_XI47/XI14/MM8_g
+ N_BLN<1>_XI47/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI14/MM5 N_XI47/XI14/NET34_XI47/XI14/MM5_d
+ N_XI47/XI14/NET33_XI47/XI14/MM5_g N_VDD_XI47/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI14/MM4 N_XI47/XI14/NET33_XI47/XI14/MM4_d
+ N_XI47/XI14/NET34_XI47/XI14/MM4_g N_VDD_XI47/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI14/MM10 N_XI47/XI14/NET35_XI47/XI14/MM10_d
+ N_XI47/XI14/NET36_XI47/XI14/MM10_g N_VDD_XI47/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI14/MM11 N_XI47/XI14/NET36_XI47/XI14/MM11_d
+ N_XI47/XI14/NET35_XI47/XI14/MM11_g N_VDD_XI47/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI15/MM2 N_XI47/XI15/NET34_XI47/XI15/MM2_d
+ N_XI47/XI15/NET33_XI47/XI15/MM2_g N_VSS_XI47/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI15/MM3 N_XI47/XI15/NET33_XI47/XI15/MM3_d N_WL<90>_XI47/XI15/MM3_g
+ N_BLN<0>_XI47/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI15/MM0 N_XI47/XI15/NET34_XI47/XI15/MM0_d N_WL<90>_XI47/XI15/MM0_g
+ N_BL<0>_XI47/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI15/MM1 N_XI47/XI15/NET33_XI47/XI15/MM1_d
+ N_XI47/XI15/NET34_XI47/XI15/MM1_g N_VSS_XI47/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI15/MM9 N_XI47/XI15/NET36_XI47/XI15/MM9_d N_WL<91>_XI47/XI15/MM9_g
+ N_BL<0>_XI47/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI15/MM6 N_XI47/XI15/NET35_XI47/XI15/MM6_d
+ N_XI47/XI15/NET36_XI47/XI15/MM6_g N_VSS_XI47/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI15/MM7 N_XI47/XI15/NET36_XI47/XI15/MM7_d
+ N_XI47/XI15/NET35_XI47/XI15/MM7_g N_VSS_XI47/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI47/XI15/MM8 N_XI47/XI15/NET35_XI47/XI15/MM8_d N_WL<91>_XI47/XI15/MM8_g
+ N_BLN<0>_XI47/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI47/XI15/MM5 N_XI47/XI15/NET34_XI47/XI15/MM5_d
+ N_XI47/XI15/NET33_XI47/XI15/MM5_g N_VDD_XI47/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI15/MM4 N_XI47/XI15/NET33_XI47/XI15/MM4_d
+ N_XI47/XI15/NET34_XI47/XI15/MM4_g N_VDD_XI47/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI15/MM10 N_XI47/XI15/NET35_XI47/XI15/MM10_d
+ N_XI47/XI15/NET36_XI47/XI15/MM10_g N_VDD_XI47/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI47/XI15/MM11 N_XI47/XI15/NET36_XI47/XI15/MM11_d
+ N_XI47/XI15/NET35_XI47/XI15/MM11_g N_VDD_XI47/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI0/MM2 N_XI48/XI0/NET34_XI48/XI0/MM2_d N_XI48/XI0/NET33_XI48/XI0/MM2_g
+ N_VSS_XI48/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI0/MM3 N_XI48/XI0/NET33_XI48/XI0/MM3_d N_WL<92>_XI48/XI0/MM3_g
+ N_BLN<15>_XI48/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI0/MM0 N_XI48/XI0/NET34_XI48/XI0/MM0_d N_WL<92>_XI48/XI0/MM0_g
+ N_BL<15>_XI48/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI0/MM1 N_XI48/XI0/NET33_XI48/XI0/MM1_d N_XI48/XI0/NET34_XI48/XI0/MM1_g
+ N_VSS_XI48/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI0/MM9 N_XI48/XI0/NET36_XI48/XI0/MM9_d N_WL<93>_XI48/XI0/MM9_g
+ N_BL<15>_XI48/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI0/MM6 N_XI48/XI0/NET35_XI48/XI0/MM6_d N_XI48/XI0/NET36_XI48/XI0/MM6_g
+ N_VSS_XI48/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI0/MM7 N_XI48/XI0/NET36_XI48/XI0/MM7_d N_XI48/XI0/NET35_XI48/XI0/MM7_g
+ N_VSS_XI48/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI0/MM8 N_XI48/XI0/NET35_XI48/XI0/MM8_d N_WL<93>_XI48/XI0/MM8_g
+ N_BLN<15>_XI48/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI0/MM5 N_XI48/XI0/NET34_XI48/XI0/MM5_d N_XI48/XI0/NET33_XI48/XI0/MM5_g
+ N_VDD_XI48/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI0/MM4 N_XI48/XI0/NET33_XI48/XI0/MM4_d N_XI48/XI0/NET34_XI48/XI0/MM4_g
+ N_VDD_XI48/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI0/MM10 N_XI48/XI0/NET35_XI48/XI0/MM10_d N_XI48/XI0/NET36_XI48/XI0/MM10_g
+ N_VDD_XI48/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI0/MM11 N_XI48/XI0/NET36_XI48/XI0/MM11_d N_XI48/XI0/NET35_XI48/XI0/MM11_g
+ N_VDD_XI48/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI1/MM2 N_XI48/XI1/NET34_XI48/XI1/MM2_d N_XI48/XI1/NET33_XI48/XI1/MM2_g
+ N_VSS_XI48/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI1/MM3 N_XI48/XI1/NET33_XI48/XI1/MM3_d N_WL<92>_XI48/XI1/MM3_g
+ N_BLN<14>_XI48/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI1/MM0 N_XI48/XI1/NET34_XI48/XI1/MM0_d N_WL<92>_XI48/XI1/MM0_g
+ N_BL<14>_XI48/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI1/MM1 N_XI48/XI1/NET33_XI48/XI1/MM1_d N_XI48/XI1/NET34_XI48/XI1/MM1_g
+ N_VSS_XI48/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI1/MM9 N_XI48/XI1/NET36_XI48/XI1/MM9_d N_WL<93>_XI48/XI1/MM9_g
+ N_BL<14>_XI48/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI1/MM6 N_XI48/XI1/NET35_XI48/XI1/MM6_d N_XI48/XI1/NET36_XI48/XI1/MM6_g
+ N_VSS_XI48/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI1/MM7 N_XI48/XI1/NET36_XI48/XI1/MM7_d N_XI48/XI1/NET35_XI48/XI1/MM7_g
+ N_VSS_XI48/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI1/MM8 N_XI48/XI1/NET35_XI48/XI1/MM8_d N_WL<93>_XI48/XI1/MM8_g
+ N_BLN<14>_XI48/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI1/MM5 N_XI48/XI1/NET34_XI48/XI1/MM5_d N_XI48/XI1/NET33_XI48/XI1/MM5_g
+ N_VDD_XI48/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI1/MM4 N_XI48/XI1/NET33_XI48/XI1/MM4_d N_XI48/XI1/NET34_XI48/XI1/MM4_g
+ N_VDD_XI48/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI1/MM10 N_XI48/XI1/NET35_XI48/XI1/MM10_d N_XI48/XI1/NET36_XI48/XI1/MM10_g
+ N_VDD_XI48/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI1/MM11 N_XI48/XI1/NET36_XI48/XI1/MM11_d N_XI48/XI1/NET35_XI48/XI1/MM11_g
+ N_VDD_XI48/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI2/MM2 N_XI48/XI2/NET34_XI48/XI2/MM2_d N_XI48/XI2/NET33_XI48/XI2/MM2_g
+ N_VSS_XI48/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI2/MM3 N_XI48/XI2/NET33_XI48/XI2/MM3_d N_WL<92>_XI48/XI2/MM3_g
+ N_BLN<13>_XI48/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI2/MM0 N_XI48/XI2/NET34_XI48/XI2/MM0_d N_WL<92>_XI48/XI2/MM0_g
+ N_BL<13>_XI48/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI2/MM1 N_XI48/XI2/NET33_XI48/XI2/MM1_d N_XI48/XI2/NET34_XI48/XI2/MM1_g
+ N_VSS_XI48/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI2/MM9 N_XI48/XI2/NET36_XI48/XI2/MM9_d N_WL<93>_XI48/XI2/MM9_g
+ N_BL<13>_XI48/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI2/MM6 N_XI48/XI2/NET35_XI48/XI2/MM6_d N_XI48/XI2/NET36_XI48/XI2/MM6_g
+ N_VSS_XI48/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI2/MM7 N_XI48/XI2/NET36_XI48/XI2/MM7_d N_XI48/XI2/NET35_XI48/XI2/MM7_g
+ N_VSS_XI48/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI2/MM8 N_XI48/XI2/NET35_XI48/XI2/MM8_d N_WL<93>_XI48/XI2/MM8_g
+ N_BLN<13>_XI48/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI2/MM5 N_XI48/XI2/NET34_XI48/XI2/MM5_d N_XI48/XI2/NET33_XI48/XI2/MM5_g
+ N_VDD_XI48/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI2/MM4 N_XI48/XI2/NET33_XI48/XI2/MM4_d N_XI48/XI2/NET34_XI48/XI2/MM4_g
+ N_VDD_XI48/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI2/MM10 N_XI48/XI2/NET35_XI48/XI2/MM10_d N_XI48/XI2/NET36_XI48/XI2/MM10_g
+ N_VDD_XI48/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI2/MM11 N_XI48/XI2/NET36_XI48/XI2/MM11_d N_XI48/XI2/NET35_XI48/XI2/MM11_g
+ N_VDD_XI48/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI3/MM2 N_XI48/XI3/NET34_XI48/XI3/MM2_d N_XI48/XI3/NET33_XI48/XI3/MM2_g
+ N_VSS_XI48/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI3/MM3 N_XI48/XI3/NET33_XI48/XI3/MM3_d N_WL<92>_XI48/XI3/MM3_g
+ N_BLN<12>_XI48/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI3/MM0 N_XI48/XI3/NET34_XI48/XI3/MM0_d N_WL<92>_XI48/XI3/MM0_g
+ N_BL<12>_XI48/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI3/MM1 N_XI48/XI3/NET33_XI48/XI3/MM1_d N_XI48/XI3/NET34_XI48/XI3/MM1_g
+ N_VSS_XI48/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI3/MM9 N_XI48/XI3/NET36_XI48/XI3/MM9_d N_WL<93>_XI48/XI3/MM9_g
+ N_BL<12>_XI48/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI3/MM6 N_XI48/XI3/NET35_XI48/XI3/MM6_d N_XI48/XI3/NET36_XI48/XI3/MM6_g
+ N_VSS_XI48/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI3/MM7 N_XI48/XI3/NET36_XI48/XI3/MM7_d N_XI48/XI3/NET35_XI48/XI3/MM7_g
+ N_VSS_XI48/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI3/MM8 N_XI48/XI3/NET35_XI48/XI3/MM8_d N_WL<93>_XI48/XI3/MM8_g
+ N_BLN<12>_XI48/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI3/MM5 N_XI48/XI3/NET34_XI48/XI3/MM5_d N_XI48/XI3/NET33_XI48/XI3/MM5_g
+ N_VDD_XI48/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI3/MM4 N_XI48/XI3/NET33_XI48/XI3/MM4_d N_XI48/XI3/NET34_XI48/XI3/MM4_g
+ N_VDD_XI48/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI3/MM10 N_XI48/XI3/NET35_XI48/XI3/MM10_d N_XI48/XI3/NET36_XI48/XI3/MM10_g
+ N_VDD_XI48/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI3/MM11 N_XI48/XI3/NET36_XI48/XI3/MM11_d N_XI48/XI3/NET35_XI48/XI3/MM11_g
+ N_VDD_XI48/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI4/MM2 N_XI48/XI4/NET34_XI48/XI4/MM2_d N_XI48/XI4/NET33_XI48/XI4/MM2_g
+ N_VSS_XI48/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI4/MM3 N_XI48/XI4/NET33_XI48/XI4/MM3_d N_WL<92>_XI48/XI4/MM3_g
+ N_BLN<11>_XI48/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI4/MM0 N_XI48/XI4/NET34_XI48/XI4/MM0_d N_WL<92>_XI48/XI4/MM0_g
+ N_BL<11>_XI48/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI4/MM1 N_XI48/XI4/NET33_XI48/XI4/MM1_d N_XI48/XI4/NET34_XI48/XI4/MM1_g
+ N_VSS_XI48/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI4/MM9 N_XI48/XI4/NET36_XI48/XI4/MM9_d N_WL<93>_XI48/XI4/MM9_g
+ N_BL<11>_XI48/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI4/MM6 N_XI48/XI4/NET35_XI48/XI4/MM6_d N_XI48/XI4/NET36_XI48/XI4/MM6_g
+ N_VSS_XI48/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI4/MM7 N_XI48/XI4/NET36_XI48/XI4/MM7_d N_XI48/XI4/NET35_XI48/XI4/MM7_g
+ N_VSS_XI48/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI4/MM8 N_XI48/XI4/NET35_XI48/XI4/MM8_d N_WL<93>_XI48/XI4/MM8_g
+ N_BLN<11>_XI48/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI4/MM5 N_XI48/XI4/NET34_XI48/XI4/MM5_d N_XI48/XI4/NET33_XI48/XI4/MM5_g
+ N_VDD_XI48/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI4/MM4 N_XI48/XI4/NET33_XI48/XI4/MM4_d N_XI48/XI4/NET34_XI48/XI4/MM4_g
+ N_VDD_XI48/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI4/MM10 N_XI48/XI4/NET35_XI48/XI4/MM10_d N_XI48/XI4/NET36_XI48/XI4/MM10_g
+ N_VDD_XI48/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI4/MM11 N_XI48/XI4/NET36_XI48/XI4/MM11_d N_XI48/XI4/NET35_XI48/XI4/MM11_g
+ N_VDD_XI48/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI5/MM2 N_XI48/XI5/NET34_XI48/XI5/MM2_d N_XI48/XI5/NET33_XI48/XI5/MM2_g
+ N_VSS_XI48/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI5/MM3 N_XI48/XI5/NET33_XI48/XI5/MM3_d N_WL<92>_XI48/XI5/MM3_g
+ N_BLN<10>_XI48/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI5/MM0 N_XI48/XI5/NET34_XI48/XI5/MM0_d N_WL<92>_XI48/XI5/MM0_g
+ N_BL<10>_XI48/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI5/MM1 N_XI48/XI5/NET33_XI48/XI5/MM1_d N_XI48/XI5/NET34_XI48/XI5/MM1_g
+ N_VSS_XI48/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI5/MM9 N_XI48/XI5/NET36_XI48/XI5/MM9_d N_WL<93>_XI48/XI5/MM9_g
+ N_BL<10>_XI48/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI5/MM6 N_XI48/XI5/NET35_XI48/XI5/MM6_d N_XI48/XI5/NET36_XI48/XI5/MM6_g
+ N_VSS_XI48/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI5/MM7 N_XI48/XI5/NET36_XI48/XI5/MM7_d N_XI48/XI5/NET35_XI48/XI5/MM7_g
+ N_VSS_XI48/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI5/MM8 N_XI48/XI5/NET35_XI48/XI5/MM8_d N_WL<93>_XI48/XI5/MM8_g
+ N_BLN<10>_XI48/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI5/MM5 N_XI48/XI5/NET34_XI48/XI5/MM5_d N_XI48/XI5/NET33_XI48/XI5/MM5_g
+ N_VDD_XI48/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI5/MM4 N_XI48/XI5/NET33_XI48/XI5/MM4_d N_XI48/XI5/NET34_XI48/XI5/MM4_g
+ N_VDD_XI48/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI5/MM10 N_XI48/XI5/NET35_XI48/XI5/MM10_d N_XI48/XI5/NET36_XI48/XI5/MM10_g
+ N_VDD_XI48/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI5/MM11 N_XI48/XI5/NET36_XI48/XI5/MM11_d N_XI48/XI5/NET35_XI48/XI5/MM11_g
+ N_VDD_XI48/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI6/MM2 N_XI48/XI6/NET34_XI48/XI6/MM2_d N_XI48/XI6/NET33_XI48/XI6/MM2_g
+ N_VSS_XI48/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM3 N_XI48/XI6/NET33_XI48/XI6/MM3_d N_WL<92>_XI48/XI6/MM3_g
+ N_BLN<9>_XI48/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM0 N_XI48/XI6/NET34_XI48/XI6/MM0_d N_WL<92>_XI48/XI6/MM0_g
+ N_BL<9>_XI48/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM1 N_XI48/XI6/NET33_XI48/XI6/MM1_d N_XI48/XI6/NET34_XI48/XI6/MM1_g
+ N_VSS_XI48/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM9 N_XI48/XI6/NET36_XI48/XI6/MM9_d N_WL<93>_XI48/XI6/MM9_g
+ N_BL<9>_XI48/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM6 N_XI48/XI6/NET35_XI48/XI6/MM6_d N_XI48/XI6/NET36_XI48/XI6/MM6_g
+ N_VSS_XI48/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM7 N_XI48/XI6/NET36_XI48/XI6/MM7_d N_XI48/XI6/NET35_XI48/XI6/MM7_g
+ N_VSS_XI48/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM8 N_XI48/XI6/NET35_XI48/XI6/MM8_d N_WL<93>_XI48/XI6/MM8_g
+ N_BLN<9>_XI48/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI6/MM5 N_XI48/XI6/NET34_XI48/XI6/MM5_d N_XI48/XI6/NET33_XI48/XI6/MM5_g
+ N_VDD_XI48/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI6/MM4 N_XI48/XI6/NET33_XI48/XI6/MM4_d N_XI48/XI6/NET34_XI48/XI6/MM4_g
+ N_VDD_XI48/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI6/MM10 N_XI48/XI6/NET35_XI48/XI6/MM10_d N_XI48/XI6/NET36_XI48/XI6/MM10_g
+ N_VDD_XI48/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI6/MM11 N_XI48/XI6/NET36_XI48/XI6/MM11_d N_XI48/XI6/NET35_XI48/XI6/MM11_g
+ N_VDD_XI48/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI7/MM2 N_XI48/XI7/NET34_XI48/XI7/MM2_d N_XI48/XI7/NET33_XI48/XI7/MM2_g
+ N_VSS_XI48/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM3 N_XI48/XI7/NET33_XI48/XI7/MM3_d N_WL<92>_XI48/XI7/MM3_g
+ N_BLN<8>_XI48/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM0 N_XI48/XI7/NET34_XI48/XI7/MM0_d N_WL<92>_XI48/XI7/MM0_g
+ N_BL<8>_XI48/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM1 N_XI48/XI7/NET33_XI48/XI7/MM1_d N_XI48/XI7/NET34_XI48/XI7/MM1_g
+ N_VSS_XI48/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM9 N_XI48/XI7/NET36_XI48/XI7/MM9_d N_WL<93>_XI48/XI7/MM9_g
+ N_BL<8>_XI48/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM6 N_XI48/XI7/NET35_XI48/XI7/MM6_d N_XI48/XI7/NET36_XI48/XI7/MM6_g
+ N_VSS_XI48/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM7 N_XI48/XI7/NET36_XI48/XI7/MM7_d N_XI48/XI7/NET35_XI48/XI7/MM7_g
+ N_VSS_XI48/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM8 N_XI48/XI7/NET35_XI48/XI7/MM8_d N_WL<93>_XI48/XI7/MM8_g
+ N_BLN<8>_XI48/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI7/MM5 N_XI48/XI7/NET34_XI48/XI7/MM5_d N_XI48/XI7/NET33_XI48/XI7/MM5_g
+ N_VDD_XI48/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI7/MM4 N_XI48/XI7/NET33_XI48/XI7/MM4_d N_XI48/XI7/NET34_XI48/XI7/MM4_g
+ N_VDD_XI48/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI7/MM10 N_XI48/XI7/NET35_XI48/XI7/MM10_d N_XI48/XI7/NET36_XI48/XI7/MM10_g
+ N_VDD_XI48/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI7/MM11 N_XI48/XI7/NET36_XI48/XI7/MM11_d N_XI48/XI7/NET35_XI48/XI7/MM11_g
+ N_VDD_XI48/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI8/MM2 N_XI48/XI8/NET34_XI48/XI8/MM2_d N_XI48/XI8/NET33_XI48/XI8/MM2_g
+ N_VSS_XI48/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM3 N_XI48/XI8/NET33_XI48/XI8/MM3_d N_WL<92>_XI48/XI8/MM3_g
+ N_BLN<7>_XI48/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM0 N_XI48/XI8/NET34_XI48/XI8/MM0_d N_WL<92>_XI48/XI8/MM0_g
+ N_BL<7>_XI48/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM1 N_XI48/XI8/NET33_XI48/XI8/MM1_d N_XI48/XI8/NET34_XI48/XI8/MM1_g
+ N_VSS_XI48/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM9 N_XI48/XI8/NET36_XI48/XI8/MM9_d N_WL<93>_XI48/XI8/MM9_g
+ N_BL<7>_XI48/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM6 N_XI48/XI8/NET35_XI48/XI8/MM6_d N_XI48/XI8/NET36_XI48/XI8/MM6_g
+ N_VSS_XI48/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM7 N_XI48/XI8/NET36_XI48/XI8/MM7_d N_XI48/XI8/NET35_XI48/XI8/MM7_g
+ N_VSS_XI48/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM8 N_XI48/XI8/NET35_XI48/XI8/MM8_d N_WL<93>_XI48/XI8/MM8_g
+ N_BLN<7>_XI48/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI8/MM5 N_XI48/XI8/NET34_XI48/XI8/MM5_d N_XI48/XI8/NET33_XI48/XI8/MM5_g
+ N_VDD_XI48/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI8/MM4 N_XI48/XI8/NET33_XI48/XI8/MM4_d N_XI48/XI8/NET34_XI48/XI8/MM4_g
+ N_VDD_XI48/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI8/MM10 N_XI48/XI8/NET35_XI48/XI8/MM10_d N_XI48/XI8/NET36_XI48/XI8/MM10_g
+ N_VDD_XI48/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI8/MM11 N_XI48/XI8/NET36_XI48/XI8/MM11_d N_XI48/XI8/NET35_XI48/XI8/MM11_g
+ N_VDD_XI48/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI9/MM2 N_XI48/XI9/NET34_XI48/XI9/MM2_d N_XI48/XI9/NET33_XI48/XI9/MM2_g
+ N_VSS_XI48/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM3 N_XI48/XI9/NET33_XI48/XI9/MM3_d N_WL<92>_XI48/XI9/MM3_g
+ N_BLN<6>_XI48/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM0 N_XI48/XI9/NET34_XI48/XI9/MM0_d N_WL<92>_XI48/XI9/MM0_g
+ N_BL<6>_XI48/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM1 N_XI48/XI9/NET33_XI48/XI9/MM1_d N_XI48/XI9/NET34_XI48/XI9/MM1_g
+ N_VSS_XI48/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM9 N_XI48/XI9/NET36_XI48/XI9/MM9_d N_WL<93>_XI48/XI9/MM9_g
+ N_BL<6>_XI48/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM6 N_XI48/XI9/NET35_XI48/XI9/MM6_d N_XI48/XI9/NET36_XI48/XI9/MM6_g
+ N_VSS_XI48/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM7 N_XI48/XI9/NET36_XI48/XI9/MM7_d N_XI48/XI9/NET35_XI48/XI9/MM7_g
+ N_VSS_XI48/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM8 N_XI48/XI9/NET35_XI48/XI9/MM8_d N_WL<93>_XI48/XI9/MM8_g
+ N_BLN<6>_XI48/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI9/MM5 N_XI48/XI9/NET34_XI48/XI9/MM5_d N_XI48/XI9/NET33_XI48/XI9/MM5_g
+ N_VDD_XI48/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI9/MM4 N_XI48/XI9/NET33_XI48/XI9/MM4_d N_XI48/XI9/NET34_XI48/XI9/MM4_g
+ N_VDD_XI48/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI9/MM10 N_XI48/XI9/NET35_XI48/XI9/MM10_d N_XI48/XI9/NET36_XI48/XI9/MM10_g
+ N_VDD_XI48/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI9/MM11 N_XI48/XI9/NET36_XI48/XI9/MM11_d N_XI48/XI9/NET35_XI48/XI9/MM11_g
+ N_VDD_XI48/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI10/MM2 N_XI48/XI10/NET34_XI48/XI10/MM2_d
+ N_XI48/XI10/NET33_XI48/XI10/MM2_g N_VSS_XI48/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI10/MM3 N_XI48/XI10/NET33_XI48/XI10/MM3_d N_WL<92>_XI48/XI10/MM3_g
+ N_BLN<5>_XI48/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI10/MM0 N_XI48/XI10/NET34_XI48/XI10/MM0_d N_WL<92>_XI48/XI10/MM0_g
+ N_BL<5>_XI48/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI10/MM1 N_XI48/XI10/NET33_XI48/XI10/MM1_d
+ N_XI48/XI10/NET34_XI48/XI10/MM1_g N_VSS_XI48/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI10/MM9 N_XI48/XI10/NET36_XI48/XI10/MM9_d N_WL<93>_XI48/XI10/MM9_g
+ N_BL<5>_XI48/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI10/MM6 N_XI48/XI10/NET35_XI48/XI10/MM6_d
+ N_XI48/XI10/NET36_XI48/XI10/MM6_g N_VSS_XI48/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI10/MM7 N_XI48/XI10/NET36_XI48/XI10/MM7_d
+ N_XI48/XI10/NET35_XI48/XI10/MM7_g N_VSS_XI48/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI10/MM8 N_XI48/XI10/NET35_XI48/XI10/MM8_d N_WL<93>_XI48/XI10/MM8_g
+ N_BLN<5>_XI48/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI10/MM5 N_XI48/XI10/NET34_XI48/XI10/MM5_d
+ N_XI48/XI10/NET33_XI48/XI10/MM5_g N_VDD_XI48/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI10/MM4 N_XI48/XI10/NET33_XI48/XI10/MM4_d
+ N_XI48/XI10/NET34_XI48/XI10/MM4_g N_VDD_XI48/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI10/MM10 N_XI48/XI10/NET35_XI48/XI10/MM10_d
+ N_XI48/XI10/NET36_XI48/XI10/MM10_g N_VDD_XI48/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI10/MM11 N_XI48/XI10/NET36_XI48/XI10/MM11_d
+ N_XI48/XI10/NET35_XI48/XI10/MM11_g N_VDD_XI48/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI11/MM2 N_XI48/XI11/NET34_XI48/XI11/MM2_d
+ N_XI48/XI11/NET33_XI48/XI11/MM2_g N_VSS_XI48/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI11/MM3 N_XI48/XI11/NET33_XI48/XI11/MM3_d N_WL<92>_XI48/XI11/MM3_g
+ N_BLN<4>_XI48/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI11/MM0 N_XI48/XI11/NET34_XI48/XI11/MM0_d N_WL<92>_XI48/XI11/MM0_g
+ N_BL<4>_XI48/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI11/MM1 N_XI48/XI11/NET33_XI48/XI11/MM1_d
+ N_XI48/XI11/NET34_XI48/XI11/MM1_g N_VSS_XI48/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI11/MM9 N_XI48/XI11/NET36_XI48/XI11/MM9_d N_WL<93>_XI48/XI11/MM9_g
+ N_BL<4>_XI48/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI11/MM6 N_XI48/XI11/NET35_XI48/XI11/MM6_d
+ N_XI48/XI11/NET36_XI48/XI11/MM6_g N_VSS_XI48/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI11/MM7 N_XI48/XI11/NET36_XI48/XI11/MM7_d
+ N_XI48/XI11/NET35_XI48/XI11/MM7_g N_VSS_XI48/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI11/MM8 N_XI48/XI11/NET35_XI48/XI11/MM8_d N_WL<93>_XI48/XI11/MM8_g
+ N_BLN<4>_XI48/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI11/MM5 N_XI48/XI11/NET34_XI48/XI11/MM5_d
+ N_XI48/XI11/NET33_XI48/XI11/MM5_g N_VDD_XI48/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI11/MM4 N_XI48/XI11/NET33_XI48/XI11/MM4_d
+ N_XI48/XI11/NET34_XI48/XI11/MM4_g N_VDD_XI48/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI11/MM10 N_XI48/XI11/NET35_XI48/XI11/MM10_d
+ N_XI48/XI11/NET36_XI48/XI11/MM10_g N_VDD_XI48/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI11/MM11 N_XI48/XI11/NET36_XI48/XI11/MM11_d
+ N_XI48/XI11/NET35_XI48/XI11/MM11_g N_VDD_XI48/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI12/MM2 N_XI48/XI12/NET34_XI48/XI12/MM2_d
+ N_XI48/XI12/NET33_XI48/XI12/MM2_g N_VSS_XI48/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI12/MM3 N_XI48/XI12/NET33_XI48/XI12/MM3_d N_WL<92>_XI48/XI12/MM3_g
+ N_BLN<3>_XI48/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI12/MM0 N_XI48/XI12/NET34_XI48/XI12/MM0_d N_WL<92>_XI48/XI12/MM0_g
+ N_BL<3>_XI48/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI12/MM1 N_XI48/XI12/NET33_XI48/XI12/MM1_d
+ N_XI48/XI12/NET34_XI48/XI12/MM1_g N_VSS_XI48/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI12/MM9 N_XI48/XI12/NET36_XI48/XI12/MM9_d N_WL<93>_XI48/XI12/MM9_g
+ N_BL<3>_XI48/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI12/MM6 N_XI48/XI12/NET35_XI48/XI12/MM6_d
+ N_XI48/XI12/NET36_XI48/XI12/MM6_g N_VSS_XI48/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI12/MM7 N_XI48/XI12/NET36_XI48/XI12/MM7_d
+ N_XI48/XI12/NET35_XI48/XI12/MM7_g N_VSS_XI48/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI12/MM8 N_XI48/XI12/NET35_XI48/XI12/MM8_d N_WL<93>_XI48/XI12/MM8_g
+ N_BLN<3>_XI48/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI12/MM5 N_XI48/XI12/NET34_XI48/XI12/MM5_d
+ N_XI48/XI12/NET33_XI48/XI12/MM5_g N_VDD_XI48/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI12/MM4 N_XI48/XI12/NET33_XI48/XI12/MM4_d
+ N_XI48/XI12/NET34_XI48/XI12/MM4_g N_VDD_XI48/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI12/MM10 N_XI48/XI12/NET35_XI48/XI12/MM10_d
+ N_XI48/XI12/NET36_XI48/XI12/MM10_g N_VDD_XI48/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI12/MM11 N_XI48/XI12/NET36_XI48/XI12/MM11_d
+ N_XI48/XI12/NET35_XI48/XI12/MM11_g N_VDD_XI48/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI13/MM2 N_XI48/XI13/NET34_XI48/XI13/MM2_d
+ N_XI48/XI13/NET33_XI48/XI13/MM2_g N_VSS_XI48/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI13/MM3 N_XI48/XI13/NET33_XI48/XI13/MM3_d N_WL<92>_XI48/XI13/MM3_g
+ N_BLN<2>_XI48/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI13/MM0 N_XI48/XI13/NET34_XI48/XI13/MM0_d N_WL<92>_XI48/XI13/MM0_g
+ N_BL<2>_XI48/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI13/MM1 N_XI48/XI13/NET33_XI48/XI13/MM1_d
+ N_XI48/XI13/NET34_XI48/XI13/MM1_g N_VSS_XI48/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI13/MM9 N_XI48/XI13/NET36_XI48/XI13/MM9_d N_WL<93>_XI48/XI13/MM9_g
+ N_BL<2>_XI48/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI13/MM6 N_XI48/XI13/NET35_XI48/XI13/MM6_d
+ N_XI48/XI13/NET36_XI48/XI13/MM6_g N_VSS_XI48/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI13/MM7 N_XI48/XI13/NET36_XI48/XI13/MM7_d
+ N_XI48/XI13/NET35_XI48/XI13/MM7_g N_VSS_XI48/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI13/MM8 N_XI48/XI13/NET35_XI48/XI13/MM8_d N_WL<93>_XI48/XI13/MM8_g
+ N_BLN<2>_XI48/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI13/MM5 N_XI48/XI13/NET34_XI48/XI13/MM5_d
+ N_XI48/XI13/NET33_XI48/XI13/MM5_g N_VDD_XI48/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI13/MM4 N_XI48/XI13/NET33_XI48/XI13/MM4_d
+ N_XI48/XI13/NET34_XI48/XI13/MM4_g N_VDD_XI48/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI13/MM10 N_XI48/XI13/NET35_XI48/XI13/MM10_d
+ N_XI48/XI13/NET36_XI48/XI13/MM10_g N_VDD_XI48/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI13/MM11 N_XI48/XI13/NET36_XI48/XI13/MM11_d
+ N_XI48/XI13/NET35_XI48/XI13/MM11_g N_VDD_XI48/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI14/MM2 N_XI48/XI14/NET34_XI48/XI14/MM2_d
+ N_XI48/XI14/NET33_XI48/XI14/MM2_g N_VSS_XI48/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI14/MM3 N_XI48/XI14/NET33_XI48/XI14/MM3_d N_WL<92>_XI48/XI14/MM3_g
+ N_BLN<1>_XI48/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI14/MM0 N_XI48/XI14/NET34_XI48/XI14/MM0_d N_WL<92>_XI48/XI14/MM0_g
+ N_BL<1>_XI48/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI14/MM1 N_XI48/XI14/NET33_XI48/XI14/MM1_d
+ N_XI48/XI14/NET34_XI48/XI14/MM1_g N_VSS_XI48/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI14/MM9 N_XI48/XI14/NET36_XI48/XI14/MM9_d N_WL<93>_XI48/XI14/MM9_g
+ N_BL<1>_XI48/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI14/MM6 N_XI48/XI14/NET35_XI48/XI14/MM6_d
+ N_XI48/XI14/NET36_XI48/XI14/MM6_g N_VSS_XI48/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI14/MM7 N_XI48/XI14/NET36_XI48/XI14/MM7_d
+ N_XI48/XI14/NET35_XI48/XI14/MM7_g N_VSS_XI48/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI14/MM8 N_XI48/XI14/NET35_XI48/XI14/MM8_d N_WL<93>_XI48/XI14/MM8_g
+ N_BLN<1>_XI48/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI14/MM5 N_XI48/XI14/NET34_XI48/XI14/MM5_d
+ N_XI48/XI14/NET33_XI48/XI14/MM5_g N_VDD_XI48/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI14/MM4 N_XI48/XI14/NET33_XI48/XI14/MM4_d
+ N_XI48/XI14/NET34_XI48/XI14/MM4_g N_VDD_XI48/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI14/MM10 N_XI48/XI14/NET35_XI48/XI14/MM10_d
+ N_XI48/XI14/NET36_XI48/XI14/MM10_g N_VDD_XI48/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI14/MM11 N_XI48/XI14/NET36_XI48/XI14/MM11_d
+ N_XI48/XI14/NET35_XI48/XI14/MM11_g N_VDD_XI48/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI15/MM2 N_XI48/XI15/NET34_XI48/XI15/MM2_d
+ N_XI48/XI15/NET33_XI48/XI15/MM2_g N_VSS_XI48/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI15/MM3 N_XI48/XI15/NET33_XI48/XI15/MM3_d N_WL<92>_XI48/XI15/MM3_g
+ N_BLN<0>_XI48/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI15/MM0 N_XI48/XI15/NET34_XI48/XI15/MM0_d N_WL<92>_XI48/XI15/MM0_g
+ N_BL<0>_XI48/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI15/MM1 N_XI48/XI15/NET33_XI48/XI15/MM1_d
+ N_XI48/XI15/NET34_XI48/XI15/MM1_g N_VSS_XI48/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI15/MM9 N_XI48/XI15/NET36_XI48/XI15/MM9_d N_WL<93>_XI48/XI15/MM9_g
+ N_BL<0>_XI48/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI15/MM6 N_XI48/XI15/NET35_XI48/XI15/MM6_d
+ N_XI48/XI15/NET36_XI48/XI15/MM6_g N_VSS_XI48/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI15/MM7 N_XI48/XI15/NET36_XI48/XI15/MM7_d
+ N_XI48/XI15/NET35_XI48/XI15/MM7_g N_VSS_XI48/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI48/XI15/MM8 N_XI48/XI15/NET35_XI48/XI15/MM8_d N_WL<93>_XI48/XI15/MM8_g
+ N_BLN<0>_XI48/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI48/XI15/MM5 N_XI48/XI15/NET34_XI48/XI15/MM5_d
+ N_XI48/XI15/NET33_XI48/XI15/MM5_g N_VDD_XI48/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI15/MM4 N_XI48/XI15/NET33_XI48/XI15/MM4_d
+ N_XI48/XI15/NET34_XI48/XI15/MM4_g N_VDD_XI48/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI15/MM10 N_XI48/XI15/NET35_XI48/XI15/MM10_d
+ N_XI48/XI15/NET36_XI48/XI15/MM10_g N_VDD_XI48/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI48/XI15/MM11 N_XI48/XI15/NET36_XI48/XI15/MM11_d
+ N_XI48/XI15/NET35_XI48/XI15/MM11_g N_VDD_XI48/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI0/MM2 N_XI49/XI0/NET34_XI49/XI0/MM2_d N_XI49/XI0/NET33_XI49/XI0/MM2_g
+ N_VSS_XI49/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI0/MM3 N_XI49/XI0/NET33_XI49/XI0/MM3_d N_WL<94>_XI49/XI0/MM3_g
+ N_BLN<15>_XI49/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI0/MM0 N_XI49/XI0/NET34_XI49/XI0/MM0_d N_WL<94>_XI49/XI0/MM0_g
+ N_BL<15>_XI49/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI0/MM1 N_XI49/XI0/NET33_XI49/XI0/MM1_d N_XI49/XI0/NET34_XI49/XI0/MM1_g
+ N_VSS_XI49/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI0/MM9 N_XI49/XI0/NET36_XI49/XI0/MM9_d N_WL<95>_XI49/XI0/MM9_g
+ N_BL<15>_XI49/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI0/MM6 N_XI49/XI0/NET35_XI49/XI0/MM6_d N_XI49/XI0/NET36_XI49/XI0/MM6_g
+ N_VSS_XI49/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI0/MM7 N_XI49/XI0/NET36_XI49/XI0/MM7_d N_XI49/XI0/NET35_XI49/XI0/MM7_g
+ N_VSS_XI49/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI0/MM8 N_XI49/XI0/NET35_XI49/XI0/MM8_d N_WL<95>_XI49/XI0/MM8_g
+ N_BLN<15>_XI49/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI0/MM5 N_XI49/XI0/NET34_XI49/XI0/MM5_d N_XI49/XI0/NET33_XI49/XI0/MM5_g
+ N_VDD_XI49/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI0/MM4 N_XI49/XI0/NET33_XI49/XI0/MM4_d N_XI49/XI0/NET34_XI49/XI0/MM4_g
+ N_VDD_XI49/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI0/MM10 N_XI49/XI0/NET35_XI49/XI0/MM10_d N_XI49/XI0/NET36_XI49/XI0/MM10_g
+ N_VDD_XI49/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI0/MM11 N_XI49/XI0/NET36_XI49/XI0/MM11_d N_XI49/XI0/NET35_XI49/XI0/MM11_g
+ N_VDD_XI49/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI1/MM2 N_XI49/XI1/NET34_XI49/XI1/MM2_d N_XI49/XI1/NET33_XI49/XI1/MM2_g
+ N_VSS_XI49/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI1/MM3 N_XI49/XI1/NET33_XI49/XI1/MM3_d N_WL<94>_XI49/XI1/MM3_g
+ N_BLN<14>_XI49/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI1/MM0 N_XI49/XI1/NET34_XI49/XI1/MM0_d N_WL<94>_XI49/XI1/MM0_g
+ N_BL<14>_XI49/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI1/MM1 N_XI49/XI1/NET33_XI49/XI1/MM1_d N_XI49/XI1/NET34_XI49/XI1/MM1_g
+ N_VSS_XI49/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI1/MM9 N_XI49/XI1/NET36_XI49/XI1/MM9_d N_WL<95>_XI49/XI1/MM9_g
+ N_BL<14>_XI49/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI1/MM6 N_XI49/XI1/NET35_XI49/XI1/MM6_d N_XI49/XI1/NET36_XI49/XI1/MM6_g
+ N_VSS_XI49/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI1/MM7 N_XI49/XI1/NET36_XI49/XI1/MM7_d N_XI49/XI1/NET35_XI49/XI1/MM7_g
+ N_VSS_XI49/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI1/MM8 N_XI49/XI1/NET35_XI49/XI1/MM8_d N_WL<95>_XI49/XI1/MM8_g
+ N_BLN<14>_XI49/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI1/MM5 N_XI49/XI1/NET34_XI49/XI1/MM5_d N_XI49/XI1/NET33_XI49/XI1/MM5_g
+ N_VDD_XI49/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI1/MM4 N_XI49/XI1/NET33_XI49/XI1/MM4_d N_XI49/XI1/NET34_XI49/XI1/MM4_g
+ N_VDD_XI49/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI1/MM10 N_XI49/XI1/NET35_XI49/XI1/MM10_d N_XI49/XI1/NET36_XI49/XI1/MM10_g
+ N_VDD_XI49/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI1/MM11 N_XI49/XI1/NET36_XI49/XI1/MM11_d N_XI49/XI1/NET35_XI49/XI1/MM11_g
+ N_VDD_XI49/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI2/MM2 N_XI49/XI2/NET34_XI49/XI2/MM2_d N_XI49/XI2/NET33_XI49/XI2/MM2_g
+ N_VSS_XI49/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI2/MM3 N_XI49/XI2/NET33_XI49/XI2/MM3_d N_WL<94>_XI49/XI2/MM3_g
+ N_BLN<13>_XI49/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI2/MM0 N_XI49/XI2/NET34_XI49/XI2/MM0_d N_WL<94>_XI49/XI2/MM0_g
+ N_BL<13>_XI49/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI2/MM1 N_XI49/XI2/NET33_XI49/XI2/MM1_d N_XI49/XI2/NET34_XI49/XI2/MM1_g
+ N_VSS_XI49/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI2/MM9 N_XI49/XI2/NET36_XI49/XI2/MM9_d N_WL<95>_XI49/XI2/MM9_g
+ N_BL<13>_XI49/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI2/MM6 N_XI49/XI2/NET35_XI49/XI2/MM6_d N_XI49/XI2/NET36_XI49/XI2/MM6_g
+ N_VSS_XI49/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI2/MM7 N_XI49/XI2/NET36_XI49/XI2/MM7_d N_XI49/XI2/NET35_XI49/XI2/MM7_g
+ N_VSS_XI49/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI2/MM8 N_XI49/XI2/NET35_XI49/XI2/MM8_d N_WL<95>_XI49/XI2/MM8_g
+ N_BLN<13>_XI49/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI2/MM5 N_XI49/XI2/NET34_XI49/XI2/MM5_d N_XI49/XI2/NET33_XI49/XI2/MM5_g
+ N_VDD_XI49/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI2/MM4 N_XI49/XI2/NET33_XI49/XI2/MM4_d N_XI49/XI2/NET34_XI49/XI2/MM4_g
+ N_VDD_XI49/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI2/MM10 N_XI49/XI2/NET35_XI49/XI2/MM10_d N_XI49/XI2/NET36_XI49/XI2/MM10_g
+ N_VDD_XI49/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI2/MM11 N_XI49/XI2/NET36_XI49/XI2/MM11_d N_XI49/XI2/NET35_XI49/XI2/MM11_g
+ N_VDD_XI49/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI3/MM2 N_XI49/XI3/NET34_XI49/XI3/MM2_d N_XI49/XI3/NET33_XI49/XI3/MM2_g
+ N_VSS_XI49/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI3/MM3 N_XI49/XI3/NET33_XI49/XI3/MM3_d N_WL<94>_XI49/XI3/MM3_g
+ N_BLN<12>_XI49/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI3/MM0 N_XI49/XI3/NET34_XI49/XI3/MM0_d N_WL<94>_XI49/XI3/MM0_g
+ N_BL<12>_XI49/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI3/MM1 N_XI49/XI3/NET33_XI49/XI3/MM1_d N_XI49/XI3/NET34_XI49/XI3/MM1_g
+ N_VSS_XI49/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI3/MM9 N_XI49/XI3/NET36_XI49/XI3/MM9_d N_WL<95>_XI49/XI3/MM9_g
+ N_BL<12>_XI49/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI3/MM6 N_XI49/XI3/NET35_XI49/XI3/MM6_d N_XI49/XI3/NET36_XI49/XI3/MM6_g
+ N_VSS_XI49/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI3/MM7 N_XI49/XI3/NET36_XI49/XI3/MM7_d N_XI49/XI3/NET35_XI49/XI3/MM7_g
+ N_VSS_XI49/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI3/MM8 N_XI49/XI3/NET35_XI49/XI3/MM8_d N_WL<95>_XI49/XI3/MM8_g
+ N_BLN<12>_XI49/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI3/MM5 N_XI49/XI3/NET34_XI49/XI3/MM5_d N_XI49/XI3/NET33_XI49/XI3/MM5_g
+ N_VDD_XI49/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI3/MM4 N_XI49/XI3/NET33_XI49/XI3/MM4_d N_XI49/XI3/NET34_XI49/XI3/MM4_g
+ N_VDD_XI49/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI3/MM10 N_XI49/XI3/NET35_XI49/XI3/MM10_d N_XI49/XI3/NET36_XI49/XI3/MM10_g
+ N_VDD_XI49/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI3/MM11 N_XI49/XI3/NET36_XI49/XI3/MM11_d N_XI49/XI3/NET35_XI49/XI3/MM11_g
+ N_VDD_XI49/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI4/MM2 N_XI49/XI4/NET34_XI49/XI4/MM2_d N_XI49/XI4/NET33_XI49/XI4/MM2_g
+ N_VSS_XI49/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI4/MM3 N_XI49/XI4/NET33_XI49/XI4/MM3_d N_WL<94>_XI49/XI4/MM3_g
+ N_BLN<11>_XI49/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI4/MM0 N_XI49/XI4/NET34_XI49/XI4/MM0_d N_WL<94>_XI49/XI4/MM0_g
+ N_BL<11>_XI49/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI4/MM1 N_XI49/XI4/NET33_XI49/XI4/MM1_d N_XI49/XI4/NET34_XI49/XI4/MM1_g
+ N_VSS_XI49/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI4/MM9 N_XI49/XI4/NET36_XI49/XI4/MM9_d N_WL<95>_XI49/XI4/MM9_g
+ N_BL<11>_XI49/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI4/MM6 N_XI49/XI4/NET35_XI49/XI4/MM6_d N_XI49/XI4/NET36_XI49/XI4/MM6_g
+ N_VSS_XI49/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI4/MM7 N_XI49/XI4/NET36_XI49/XI4/MM7_d N_XI49/XI4/NET35_XI49/XI4/MM7_g
+ N_VSS_XI49/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI4/MM8 N_XI49/XI4/NET35_XI49/XI4/MM8_d N_WL<95>_XI49/XI4/MM8_g
+ N_BLN<11>_XI49/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI4/MM5 N_XI49/XI4/NET34_XI49/XI4/MM5_d N_XI49/XI4/NET33_XI49/XI4/MM5_g
+ N_VDD_XI49/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI4/MM4 N_XI49/XI4/NET33_XI49/XI4/MM4_d N_XI49/XI4/NET34_XI49/XI4/MM4_g
+ N_VDD_XI49/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI4/MM10 N_XI49/XI4/NET35_XI49/XI4/MM10_d N_XI49/XI4/NET36_XI49/XI4/MM10_g
+ N_VDD_XI49/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI4/MM11 N_XI49/XI4/NET36_XI49/XI4/MM11_d N_XI49/XI4/NET35_XI49/XI4/MM11_g
+ N_VDD_XI49/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI5/MM2 N_XI49/XI5/NET34_XI49/XI5/MM2_d N_XI49/XI5/NET33_XI49/XI5/MM2_g
+ N_VSS_XI49/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI5/MM3 N_XI49/XI5/NET33_XI49/XI5/MM3_d N_WL<94>_XI49/XI5/MM3_g
+ N_BLN<10>_XI49/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI5/MM0 N_XI49/XI5/NET34_XI49/XI5/MM0_d N_WL<94>_XI49/XI5/MM0_g
+ N_BL<10>_XI49/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI5/MM1 N_XI49/XI5/NET33_XI49/XI5/MM1_d N_XI49/XI5/NET34_XI49/XI5/MM1_g
+ N_VSS_XI49/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI5/MM9 N_XI49/XI5/NET36_XI49/XI5/MM9_d N_WL<95>_XI49/XI5/MM9_g
+ N_BL<10>_XI49/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI5/MM6 N_XI49/XI5/NET35_XI49/XI5/MM6_d N_XI49/XI5/NET36_XI49/XI5/MM6_g
+ N_VSS_XI49/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI5/MM7 N_XI49/XI5/NET36_XI49/XI5/MM7_d N_XI49/XI5/NET35_XI49/XI5/MM7_g
+ N_VSS_XI49/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI5/MM8 N_XI49/XI5/NET35_XI49/XI5/MM8_d N_WL<95>_XI49/XI5/MM8_g
+ N_BLN<10>_XI49/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI5/MM5 N_XI49/XI5/NET34_XI49/XI5/MM5_d N_XI49/XI5/NET33_XI49/XI5/MM5_g
+ N_VDD_XI49/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI5/MM4 N_XI49/XI5/NET33_XI49/XI5/MM4_d N_XI49/XI5/NET34_XI49/XI5/MM4_g
+ N_VDD_XI49/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI5/MM10 N_XI49/XI5/NET35_XI49/XI5/MM10_d N_XI49/XI5/NET36_XI49/XI5/MM10_g
+ N_VDD_XI49/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI5/MM11 N_XI49/XI5/NET36_XI49/XI5/MM11_d N_XI49/XI5/NET35_XI49/XI5/MM11_g
+ N_VDD_XI49/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI6/MM2 N_XI49/XI6/NET34_XI49/XI6/MM2_d N_XI49/XI6/NET33_XI49/XI6/MM2_g
+ N_VSS_XI49/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM3 N_XI49/XI6/NET33_XI49/XI6/MM3_d N_WL<94>_XI49/XI6/MM3_g
+ N_BLN<9>_XI49/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM0 N_XI49/XI6/NET34_XI49/XI6/MM0_d N_WL<94>_XI49/XI6/MM0_g
+ N_BL<9>_XI49/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM1 N_XI49/XI6/NET33_XI49/XI6/MM1_d N_XI49/XI6/NET34_XI49/XI6/MM1_g
+ N_VSS_XI49/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM9 N_XI49/XI6/NET36_XI49/XI6/MM9_d N_WL<95>_XI49/XI6/MM9_g
+ N_BL<9>_XI49/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM6 N_XI49/XI6/NET35_XI49/XI6/MM6_d N_XI49/XI6/NET36_XI49/XI6/MM6_g
+ N_VSS_XI49/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM7 N_XI49/XI6/NET36_XI49/XI6/MM7_d N_XI49/XI6/NET35_XI49/XI6/MM7_g
+ N_VSS_XI49/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM8 N_XI49/XI6/NET35_XI49/XI6/MM8_d N_WL<95>_XI49/XI6/MM8_g
+ N_BLN<9>_XI49/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI6/MM5 N_XI49/XI6/NET34_XI49/XI6/MM5_d N_XI49/XI6/NET33_XI49/XI6/MM5_g
+ N_VDD_XI49/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI6/MM4 N_XI49/XI6/NET33_XI49/XI6/MM4_d N_XI49/XI6/NET34_XI49/XI6/MM4_g
+ N_VDD_XI49/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI6/MM10 N_XI49/XI6/NET35_XI49/XI6/MM10_d N_XI49/XI6/NET36_XI49/XI6/MM10_g
+ N_VDD_XI49/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI6/MM11 N_XI49/XI6/NET36_XI49/XI6/MM11_d N_XI49/XI6/NET35_XI49/XI6/MM11_g
+ N_VDD_XI49/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI7/MM2 N_XI49/XI7/NET34_XI49/XI7/MM2_d N_XI49/XI7/NET33_XI49/XI7/MM2_g
+ N_VSS_XI49/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM3 N_XI49/XI7/NET33_XI49/XI7/MM3_d N_WL<94>_XI49/XI7/MM3_g
+ N_BLN<8>_XI49/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM0 N_XI49/XI7/NET34_XI49/XI7/MM0_d N_WL<94>_XI49/XI7/MM0_g
+ N_BL<8>_XI49/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM1 N_XI49/XI7/NET33_XI49/XI7/MM1_d N_XI49/XI7/NET34_XI49/XI7/MM1_g
+ N_VSS_XI49/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM9 N_XI49/XI7/NET36_XI49/XI7/MM9_d N_WL<95>_XI49/XI7/MM9_g
+ N_BL<8>_XI49/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM6 N_XI49/XI7/NET35_XI49/XI7/MM6_d N_XI49/XI7/NET36_XI49/XI7/MM6_g
+ N_VSS_XI49/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM7 N_XI49/XI7/NET36_XI49/XI7/MM7_d N_XI49/XI7/NET35_XI49/XI7/MM7_g
+ N_VSS_XI49/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM8 N_XI49/XI7/NET35_XI49/XI7/MM8_d N_WL<95>_XI49/XI7/MM8_g
+ N_BLN<8>_XI49/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI7/MM5 N_XI49/XI7/NET34_XI49/XI7/MM5_d N_XI49/XI7/NET33_XI49/XI7/MM5_g
+ N_VDD_XI49/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI7/MM4 N_XI49/XI7/NET33_XI49/XI7/MM4_d N_XI49/XI7/NET34_XI49/XI7/MM4_g
+ N_VDD_XI49/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI7/MM10 N_XI49/XI7/NET35_XI49/XI7/MM10_d N_XI49/XI7/NET36_XI49/XI7/MM10_g
+ N_VDD_XI49/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI7/MM11 N_XI49/XI7/NET36_XI49/XI7/MM11_d N_XI49/XI7/NET35_XI49/XI7/MM11_g
+ N_VDD_XI49/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI8/MM2 N_XI49/XI8/NET34_XI49/XI8/MM2_d N_XI49/XI8/NET33_XI49/XI8/MM2_g
+ N_VSS_XI49/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM3 N_XI49/XI8/NET33_XI49/XI8/MM3_d N_WL<94>_XI49/XI8/MM3_g
+ N_BLN<7>_XI49/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM0 N_XI49/XI8/NET34_XI49/XI8/MM0_d N_WL<94>_XI49/XI8/MM0_g
+ N_BL<7>_XI49/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM1 N_XI49/XI8/NET33_XI49/XI8/MM1_d N_XI49/XI8/NET34_XI49/XI8/MM1_g
+ N_VSS_XI49/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM9 N_XI49/XI8/NET36_XI49/XI8/MM9_d N_WL<95>_XI49/XI8/MM9_g
+ N_BL<7>_XI49/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM6 N_XI49/XI8/NET35_XI49/XI8/MM6_d N_XI49/XI8/NET36_XI49/XI8/MM6_g
+ N_VSS_XI49/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM7 N_XI49/XI8/NET36_XI49/XI8/MM7_d N_XI49/XI8/NET35_XI49/XI8/MM7_g
+ N_VSS_XI49/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM8 N_XI49/XI8/NET35_XI49/XI8/MM8_d N_WL<95>_XI49/XI8/MM8_g
+ N_BLN<7>_XI49/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI8/MM5 N_XI49/XI8/NET34_XI49/XI8/MM5_d N_XI49/XI8/NET33_XI49/XI8/MM5_g
+ N_VDD_XI49/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI8/MM4 N_XI49/XI8/NET33_XI49/XI8/MM4_d N_XI49/XI8/NET34_XI49/XI8/MM4_g
+ N_VDD_XI49/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI8/MM10 N_XI49/XI8/NET35_XI49/XI8/MM10_d N_XI49/XI8/NET36_XI49/XI8/MM10_g
+ N_VDD_XI49/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI8/MM11 N_XI49/XI8/NET36_XI49/XI8/MM11_d N_XI49/XI8/NET35_XI49/XI8/MM11_g
+ N_VDD_XI49/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI9/MM2 N_XI49/XI9/NET34_XI49/XI9/MM2_d N_XI49/XI9/NET33_XI49/XI9/MM2_g
+ N_VSS_XI49/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM3 N_XI49/XI9/NET33_XI49/XI9/MM3_d N_WL<94>_XI49/XI9/MM3_g
+ N_BLN<6>_XI49/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM0 N_XI49/XI9/NET34_XI49/XI9/MM0_d N_WL<94>_XI49/XI9/MM0_g
+ N_BL<6>_XI49/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM1 N_XI49/XI9/NET33_XI49/XI9/MM1_d N_XI49/XI9/NET34_XI49/XI9/MM1_g
+ N_VSS_XI49/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM9 N_XI49/XI9/NET36_XI49/XI9/MM9_d N_WL<95>_XI49/XI9/MM9_g
+ N_BL<6>_XI49/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM6 N_XI49/XI9/NET35_XI49/XI9/MM6_d N_XI49/XI9/NET36_XI49/XI9/MM6_g
+ N_VSS_XI49/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM7 N_XI49/XI9/NET36_XI49/XI9/MM7_d N_XI49/XI9/NET35_XI49/XI9/MM7_g
+ N_VSS_XI49/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM8 N_XI49/XI9/NET35_XI49/XI9/MM8_d N_WL<95>_XI49/XI9/MM8_g
+ N_BLN<6>_XI49/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI9/MM5 N_XI49/XI9/NET34_XI49/XI9/MM5_d N_XI49/XI9/NET33_XI49/XI9/MM5_g
+ N_VDD_XI49/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI9/MM4 N_XI49/XI9/NET33_XI49/XI9/MM4_d N_XI49/XI9/NET34_XI49/XI9/MM4_g
+ N_VDD_XI49/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI9/MM10 N_XI49/XI9/NET35_XI49/XI9/MM10_d N_XI49/XI9/NET36_XI49/XI9/MM10_g
+ N_VDD_XI49/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI9/MM11 N_XI49/XI9/NET36_XI49/XI9/MM11_d N_XI49/XI9/NET35_XI49/XI9/MM11_g
+ N_VDD_XI49/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI10/MM2 N_XI49/XI10/NET34_XI49/XI10/MM2_d
+ N_XI49/XI10/NET33_XI49/XI10/MM2_g N_VSS_XI49/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI10/MM3 N_XI49/XI10/NET33_XI49/XI10/MM3_d N_WL<94>_XI49/XI10/MM3_g
+ N_BLN<5>_XI49/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI10/MM0 N_XI49/XI10/NET34_XI49/XI10/MM0_d N_WL<94>_XI49/XI10/MM0_g
+ N_BL<5>_XI49/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI10/MM1 N_XI49/XI10/NET33_XI49/XI10/MM1_d
+ N_XI49/XI10/NET34_XI49/XI10/MM1_g N_VSS_XI49/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI10/MM9 N_XI49/XI10/NET36_XI49/XI10/MM9_d N_WL<95>_XI49/XI10/MM9_g
+ N_BL<5>_XI49/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI10/MM6 N_XI49/XI10/NET35_XI49/XI10/MM6_d
+ N_XI49/XI10/NET36_XI49/XI10/MM6_g N_VSS_XI49/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI10/MM7 N_XI49/XI10/NET36_XI49/XI10/MM7_d
+ N_XI49/XI10/NET35_XI49/XI10/MM7_g N_VSS_XI49/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI10/MM8 N_XI49/XI10/NET35_XI49/XI10/MM8_d N_WL<95>_XI49/XI10/MM8_g
+ N_BLN<5>_XI49/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI10/MM5 N_XI49/XI10/NET34_XI49/XI10/MM5_d
+ N_XI49/XI10/NET33_XI49/XI10/MM5_g N_VDD_XI49/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI10/MM4 N_XI49/XI10/NET33_XI49/XI10/MM4_d
+ N_XI49/XI10/NET34_XI49/XI10/MM4_g N_VDD_XI49/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI10/MM10 N_XI49/XI10/NET35_XI49/XI10/MM10_d
+ N_XI49/XI10/NET36_XI49/XI10/MM10_g N_VDD_XI49/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI10/MM11 N_XI49/XI10/NET36_XI49/XI10/MM11_d
+ N_XI49/XI10/NET35_XI49/XI10/MM11_g N_VDD_XI49/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI11/MM2 N_XI49/XI11/NET34_XI49/XI11/MM2_d
+ N_XI49/XI11/NET33_XI49/XI11/MM2_g N_VSS_XI49/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI11/MM3 N_XI49/XI11/NET33_XI49/XI11/MM3_d N_WL<94>_XI49/XI11/MM3_g
+ N_BLN<4>_XI49/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI11/MM0 N_XI49/XI11/NET34_XI49/XI11/MM0_d N_WL<94>_XI49/XI11/MM0_g
+ N_BL<4>_XI49/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI11/MM1 N_XI49/XI11/NET33_XI49/XI11/MM1_d
+ N_XI49/XI11/NET34_XI49/XI11/MM1_g N_VSS_XI49/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI11/MM9 N_XI49/XI11/NET36_XI49/XI11/MM9_d N_WL<95>_XI49/XI11/MM9_g
+ N_BL<4>_XI49/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI11/MM6 N_XI49/XI11/NET35_XI49/XI11/MM6_d
+ N_XI49/XI11/NET36_XI49/XI11/MM6_g N_VSS_XI49/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI11/MM7 N_XI49/XI11/NET36_XI49/XI11/MM7_d
+ N_XI49/XI11/NET35_XI49/XI11/MM7_g N_VSS_XI49/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI11/MM8 N_XI49/XI11/NET35_XI49/XI11/MM8_d N_WL<95>_XI49/XI11/MM8_g
+ N_BLN<4>_XI49/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI11/MM5 N_XI49/XI11/NET34_XI49/XI11/MM5_d
+ N_XI49/XI11/NET33_XI49/XI11/MM5_g N_VDD_XI49/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI11/MM4 N_XI49/XI11/NET33_XI49/XI11/MM4_d
+ N_XI49/XI11/NET34_XI49/XI11/MM4_g N_VDD_XI49/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI11/MM10 N_XI49/XI11/NET35_XI49/XI11/MM10_d
+ N_XI49/XI11/NET36_XI49/XI11/MM10_g N_VDD_XI49/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI11/MM11 N_XI49/XI11/NET36_XI49/XI11/MM11_d
+ N_XI49/XI11/NET35_XI49/XI11/MM11_g N_VDD_XI49/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI12/MM2 N_XI49/XI12/NET34_XI49/XI12/MM2_d
+ N_XI49/XI12/NET33_XI49/XI12/MM2_g N_VSS_XI49/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI12/MM3 N_XI49/XI12/NET33_XI49/XI12/MM3_d N_WL<94>_XI49/XI12/MM3_g
+ N_BLN<3>_XI49/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI12/MM0 N_XI49/XI12/NET34_XI49/XI12/MM0_d N_WL<94>_XI49/XI12/MM0_g
+ N_BL<3>_XI49/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI12/MM1 N_XI49/XI12/NET33_XI49/XI12/MM1_d
+ N_XI49/XI12/NET34_XI49/XI12/MM1_g N_VSS_XI49/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI12/MM9 N_XI49/XI12/NET36_XI49/XI12/MM9_d N_WL<95>_XI49/XI12/MM9_g
+ N_BL<3>_XI49/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI12/MM6 N_XI49/XI12/NET35_XI49/XI12/MM6_d
+ N_XI49/XI12/NET36_XI49/XI12/MM6_g N_VSS_XI49/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI12/MM7 N_XI49/XI12/NET36_XI49/XI12/MM7_d
+ N_XI49/XI12/NET35_XI49/XI12/MM7_g N_VSS_XI49/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI12/MM8 N_XI49/XI12/NET35_XI49/XI12/MM8_d N_WL<95>_XI49/XI12/MM8_g
+ N_BLN<3>_XI49/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI12/MM5 N_XI49/XI12/NET34_XI49/XI12/MM5_d
+ N_XI49/XI12/NET33_XI49/XI12/MM5_g N_VDD_XI49/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI12/MM4 N_XI49/XI12/NET33_XI49/XI12/MM4_d
+ N_XI49/XI12/NET34_XI49/XI12/MM4_g N_VDD_XI49/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI12/MM10 N_XI49/XI12/NET35_XI49/XI12/MM10_d
+ N_XI49/XI12/NET36_XI49/XI12/MM10_g N_VDD_XI49/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI12/MM11 N_XI49/XI12/NET36_XI49/XI12/MM11_d
+ N_XI49/XI12/NET35_XI49/XI12/MM11_g N_VDD_XI49/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI13/MM2 N_XI49/XI13/NET34_XI49/XI13/MM2_d
+ N_XI49/XI13/NET33_XI49/XI13/MM2_g N_VSS_XI49/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI13/MM3 N_XI49/XI13/NET33_XI49/XI13/MM3_d N_WL<94>_XI49/XI13/MM3_g
+ N_BLN<2>_XI49/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI13/MM0 N_XI49/XI13/NET34_XI49/XI13/MM0_d N_WL<94>_XI49/XI13/MM0_g
+ N_BL<2>_XI49/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI13/MM1 N_XI49/XI13/NET33_XI49/XI13/MM1_d
+ N_XI49/XI13/NET34_XI49/XI13/MM1_g N_VSS_XI49/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI13/MM9 N_XI49/XI13/NET36_XI49/XI13/MM9_d N_WL<95>_XI49/XI13/MM9_g
+ N_BL<2>_XI49/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI13/MM6 N_XI49/XI13/NET35_XI49/XI13/MM6_d
+ N_XI49/XI13/NET36_XI49/XI13/MM6_g N_VSS_XI49/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI13/MM7 N_XI49/XI13/NET36_XI49/XI13/MM7_d
+ N_XI49/XI13/NET35_XI49/XI13/MM7_g N_VSS_XI49/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI13/MM8 N_XI49/XI13/NET35_XI49/XI13/MM8_d N_WL<95>_XI49/XI13/MM8_g
+ N_BLN<2>_XI49/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI13/MM5 N_XI49/XI13/NET34_XI49/XI13/MM5_d
+ N_XI49/XI13/NET33_XI49/XI13/MM5_g N_VDD_XI49/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI13/MM4 N_XI49/XI13/NET33_XI49/XI13/MM4_d
+ N_XI49/XI13/NET34_XI49/XI13/MM4_g N_VDD_XI49/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI13/MM10 N_XI49/XI13/NET35_XI49/XI13/MM10_d
+ N_XI49/XI13/NET36_XI49/XI13/MM10_g N_VDD_XI49/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI13/MM11 N_XI49/XI13/NET36_XI49/XI13/MM11_d
+ N_XI49/XI13/NET35_XI49/XI13/MM11_g N_VDD_XI49/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI14/MM2 N_XI49/XI14/NET34_XI49/XI14/MM2_d
+ N_XI49/XI14/NET33_XI49/XI14/MM2_g N_VSS_XI49/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI14/MM3 N_XI49/XI14/NET33_XI49/XI14/MM3_d N_WL<94>_XI49/XI14/MM3_g
+ N_BLN<1>_XI49/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI14/MM0 N_XI49/XI14/NET34_XI49/XI14/MM0_d N_WL<94>_XI49/XI14/MM0_g
+ N_BL<1>_XI49/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI14/MM1 N_XI49/XI14/NET33_XI49/XI14/MM1_d
+ N_XI49/XI14/NET34_XI49/XI14/MM1_g N_VSS_XI49/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI14/MM9 N_XI49/XI14/NET36_XI49/XI14/MM9_d N_WL<95>_XI49/XI14/MM9_g
+ N_BL<1>_XI49/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI14/MM6 N_XI49/XI14/NET35_XI49/XI14/MM6_d
+ N_XI49/XI14/NET36_XI49/XI14/MM6_g N_VSS_XI49/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI14/MM7 N_XI49/XI14/NET36_XI49/XI14/MM7_d
+ N_XI49/XI14/NET35_XI49/XI14/MM7_g N_VSS_XI49/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI14/MM8 N_XI49/XI14/NET35_XI49/XI14/MM8_d N_WL<95>_XI49/XI14/MM8_g
+ N_BLN<1>_XI49/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI14/MM5 N_XI49/XI14/NET34_XI49/XI14/MM5_d
+ N_XI49/XI14/NET33_XI49/XI14/MM5_g N_VDD_XI49/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI14/MM4 N_XI49/XI14/NET33_XI49/XI14/MM4_d
+ N_XI49/XI14/NET34_XI49/XI14/MM4_g N_VDD_XI49/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI14/MM10 N_XI49/XI14/NET35_XI49/XI14/MM10_d
+ N_XI49/XI14/NET36_XI49/XI14/MM10_g N_VDD_XI49/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI14/MM11 N_XI49/XI14/NET36_XI49/XI14/MM11_d
+ N_XI49/XI14/NET35_XI49/XI14/MM11_g N_VDD_XI49/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI15/MM2 N_XI49/XI15/NET34_XI49/XI15/MM2_d
+ N_XI49/XI15/NET33_XI49/XI15/MM2_g N_VSS_XI49/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI15/MM3 N_XI49/XI15/NET33_XI49/XI15/MM3_d N_WL<94>_XI49/XI15/MM3_g
+ N_BLN<0>_XI49/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI15/MM0 N_XI49/XI15/NET34_XI49/XI15/MM0_d N_WL<94>_XI49/XI15/MM0_g
+ N_BL<0>_XI49/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI15/MM1 N_XI49/XI15/NET33_XI49/XI15/MM1_d
+ N_XI49/XI15/NET34_XI49/XI15/MM1_g N_VSS_XI49/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI15/MM9 N_XI49/XI15/NET36_XI49/XI15/MM9_d N_WL<95>_XI49/XI15/MM9_g
+ N_BL<0>_XI49/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI15/MM6 N_XI49/XI15/NET35_XI49/XI15/MM6_d
+ N_XI49/XI15/NET36_XI49/XI15/MM6_g N_VSS_XI49/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI15/MM7 N_XI49/XI15/NET36_XI49/XI15/MM7_d
+ N_XI49/XI15/NET35_XI49/XI15/MM7_g N_VSS_XI49/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI49/XI15/MM8 N_XI49/XI15/NET35_XI49/XI15/MM8_d N_WL<95>_XI49/XI15/MM8_g
+ N_BLN<0>_XI49/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI49/XI15/MM5 N_XI49/XI15/NET34_XI49/XI15/MM5_d
+ N_XI49/XI15/NET33_XI49/XI15/MM5_g N_VDD_XI49/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI15/MM4 N_XI49/XI15/NET33_XI49/XI15/MM4_d
+ N_XI49/XI15/NET34_XI49/XI15/MM4_g N_VDD_XI49/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI15/MM10 N_XI49/XI15/NET35_XI49/XI15/MM10_d
+ N_XI49/XI15/NET36_XI49/XI15/MM10_g N_VDD_XI49/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI49/XI15/MM11 N_XI49/XI15/NET36_XI49/XI15/MM11_d
+ N_XI49/XI15/NET35_XI49/XI15/MM11_g N_VDD_XI49/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI0/MM2 N_XI50/XI0/NET34_XI50/XI0/MM2_d N_XI50/XI0/NET33_XI50/XI0/MM2_g
+ N_VSS_XI50/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI0/MM3 N_XI50/XI0/NET33_XI50/XI0/MM3_d N_WL<96>_XI50/XI0/MM3_g
+ N_BLN<15>_XI50/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI0/MM0 N_XI50/XI0/NET34_XI50/XI0/MM0_d N_WL<96>_XI50/XI0/MM0_g
+ N_BL<15>_XI50/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI0/MM1 N_XI50/XI0/NET33_XI50/XI0/MM1_d N_XI50/XI0/NET34_XI50/XI0/MM1_g
+ N_VSS_XI50/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI0/MM9 N_XI50/XI0/NET36_XI50/XI0/MM9_d N_WL<97>_XI50/XI0/MM9_g
+ N_BL<15>_XI50/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI0/MM6 N_XI50/XI0/NET35_XI50/XI0/MM6_d N_XI50/XI0/NET36_XI50/XI0/MM6_g
+ N_VSS_XI50/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI0/MM7 N_XI50/XI0/NET36_XI50/XI0/MM7_d N_XI50/XI0/NET35_XI50/XI0/MM7_g
+ N_VSS_XI50/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI0/MM8 N_XI50/XI0/NET35_XI50/XI0/MM8_d N_WL<97>_XI50/XI0/MM8_g
+ N_BLN<15>_XI50/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI0/MM5 N_XI50/XI0/NET34_XI50/XI0/MM5_d N_XI50/XI0/NET33_XI50/XI0/MM5_g
+ N_VDD_XI50/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI0/MM4 N_XI50/XI0/NET33_XI50/XI0/MM4_d N_XI50/XI0/NET34_XI50/XI0/MM4_g
+ N_VDD_XI50/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI0/MM10 N_XI50/XI0/NET35_XI50/XI0/MM10_d N_XI50/XI0/NET36_XI50/XI0/MM10_g
+ N_VDD_XI50/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI0/MM11 N_XI50/XI0/NET36_XI50/XI0/MM11_d N_XI50/XI0/NET35_XI50/XI0/MM11_g
+ N_VDD_XI50/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI1/MM2 N_XI50/XI1/NET34_XI50/XI1/MM2_d N_XI50/XI1/NET33_XI50/XI1/MM2_g
+ N_VSS_XI50/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI1/MM3 N_XI50/XI1/NET33_XI50/XI1/MM3_d N_WL<96>_XI50/XI1/MM3_g
+ N_BLN<14>_XI50/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI1/MM0 N_XI50/XI1/NET34_XI50/XI1/MM0_d N_WL<96>_XI50/XI1/MM0_g
+ N_BL<14>_XI50/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI1/MM1 N_XI50/XI1/NET33_XI50/XI1/MM1_d N_XI50/XI1/NET34_XI50/XI1/MM1_g
+ N_VSS_XI50/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI1/MM9 N_XI50/XI1/NET36_XI50/XI1/MM9_d N_WL<97>_XI50/XI1/MM9_g
+ N_BL<14>_XI50/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI1/MM6 N_XI50/XI1/NET35_XI50/XI1/MM6_d N_XI50/XI1/NET36_XI50/XI1/MM6_g
+ N_VSS_XI50/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI1/MM7 N_XI50/XI1/NET36_XI50/XI1/MM7_d N_XI50/XI1/NET35_XI50/XI1/MM7_g
+ N_VSS_XI50/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI1/MM8 N_XI50/XI1/NET35_XI50/XI1/MM8_d N_WL<97>_XI50/XI1/MM8_g
+ N_BLN<14>_XI50/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI1/MM5 N_XI50/XI1/NET34_XI50/XI1/MM5_d N_XI50/XI1/NET33_XI50/XI1/MM5_g
+ N_VDD_XI50/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI1/MM4 N_XI50/XI1/NET33_XI50/XI1/MM4_d N_XI50/XI1/NET34_XI50/XI1/MM4_g
+ N_VDD_XI50/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI1/MM10 N_XI50/XI1/NET35_XI50/XI1/MM10_d N_XI50/XI1/NET36_XI50/XI1/MM10_g
+ N_VDD_XI50/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI1/MM11 N_XI50/XI1/NET36_XI50/XI1/MM11_d N_XI50/XI1/NET35_XI50/XI1/MM11_g
+ N_VDD_XI50/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI2/MM2 N_XI50/XI2/NET34_XI50/XI2/MM2_d N_XI50/XI2/NET33_XI50/XI2/MM2_g
+ N_VSS_XI50/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI2/MM3 N_XI50/XI2/NET33_XI50/XI2/MM3_d N_WL<96>_XI50/XI2/MM3_g
+ N_BLN<13>_XI50/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI2/MM0 N_XI50/XI2/NET34_XI50/XI2/MM0_d N_WL<96>_XI50/XI2/MM0_g
+ N_BL<13>_XI50/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI2/MM1 N_XI50/XI2/NET33_XI50/XI2/MM1_d N_XI50/XI2/NET34_XI50/XI2/MM1_g
+ N_VSS_XI50/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI2/MM9 N_XI50/XI2/NET36_XI50/XI2/MM9_d N_WL<97>_XI50/XI2/MM9_g
+ N_BL<13>_XI50/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI2/MM6 N_XI50/XI2/NET35_XI50/XI2/MM6_d N_XI50/XI2/NET36_XI50/XI2/MM6_g
+ N_VSS_XI50/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI2/MM7 N_XI50/XI2/NET36_XI50/XI2/MM7_d N_XI50/XI2/NET35_XI50/XI2/MM7_g
+ N_VSS_XI50/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI2/MM8 N_XI50/XI2/NET35_XI50/XI2/MM8_d N_WL<97>_XI50/XI2/MM8_g
+ N_BLN<13>_XI50/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI2/MM5 N_XI50/XI2/NET34_XI50/XI2/MM5_d N_XI50/XI2/NET33_XI50/XI2/MM5_g
+ N_VDD_XI50/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI2/MM4 N_XI50/XI2/NET33_XI50/XI2/MM4_d N_XI50/XI2/NET34_XI50/XI2/MM4_g
+ N_VDD_XI50/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI2/MM10 N_XI50/XI2/NET35_XI50/XI2/MM10_d N_XI50/XI2/NET36_XI50/XI2/MM10_g
+ N_VDD_XI50/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI2/MM11 N_XI50/XI2/NET36_XI50/XI2/MM11_d N_XI50/XI2/NET35_XI50/XI2/MM11_g
+ N_VDD_XI50/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI3/MM2 N_XI50/XI3/NET34_XI50/XI3/MM2_d N_XI50/XI3/NET33_XI50/XI3/MM2_g
+ N_VSS_XI50/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI3/MM3 N_XI50/XI3/NET33_XI50/XI3/MM3_d N_WL<96>_XI50/XI3/MM3_g
+ N_BLN<12>_XI50/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI3/MM0 N_XI50/XI3/NET34_XI50/XI3/MM0_d N_WL<96>_XI50/XI3/MM0_g
+ N_BL<12>_XI50/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI3/MM1 N_XI50/XI3/NET33_XI50/XI3/MM1_d N_XI50/XI3/NET34_XI50/XI3/MM1_g
+ N_VSS_XI50/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI3/MM9 N_XI50/XI3/NET36_XI50/XI3/MM9_d N_WL<97>_XI50/XI3/MM9_g
+ N_BL<12>_XI50/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI3/MM6 N_XI50/XI3/NET35_XI50/XI3/MM6_d N_XI50/XI3/NET36_XI50/XI3/MM6_g
+ N_VSS_XI50/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI3/MM7 N_XI50/XI3/NET36_XI50/XI3/MM7_d N_XI50/XI3/NET35_XI50/XI3/MM7_g
+ N_VSS_XI50/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI3/MM8 N_XI50/XI3/NET35_XI50/XI3/MM8_d N_WL<97>_XI50/XI3/MM8_g
+ N_BLN<12>_XI50/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI3/MM5 N_XI50/XI3/NET34_XI50/XI3/MM5_d N_XI50/XI3/NET33_XI50/XI3/MM5_g
+ N_VDD_XI50/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI3/MM4 N_XI50/XI3/NET33_XI50/XI3/MM4_d N_XI50/XI3/NET34_XI50/XI3/MM4_g
+ N_VDD_XI50/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI3/MM10 N_XI50/XI3/NET35_XI50/XI3/MM10_d N_XI50/XI3/NET36_XI50/XI3/MM10_g
+ N_VDD_XI50/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI3/MM11 N_XI50/XI3/NET36_XI50/XI3/MM11_d N_XI50/XI3/NET35_XI50/XI3/MM11_g
+ N_VDD_XI50/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI4/MM2 N_XI50/XI4/NET34_XI50/XI4/MM2_d N_XI50/XI4/NET33_XI50/XI4/MM2_g
+ N_VSS_XI50/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI4/MM3 N_XI50/XI4/NET33_XI50/XI4/MM3_d N_WL<96>_XI50/XI4/MM3_g
+ N_BLN<11>_XI50/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI4/MM0 N_XI50/XI4/NET34_XI50/XI4/MM0_d N_WL<96>_XI50/XI4/MM0_g
+ N_BL<11>_XI50/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI4/MM1 N_XI50/XI4/NET33_XI50/XI4/MM1_d N_XI50/XI4/NET34_XI50/XI4/MM1_g
+ N_VSS_XI50/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI4/MM9 N_XI50/XI4/NET36_XI50/XI4/MM9_d N_WL<97>_XI50/XI4/MM9_g
+ N_BL<11>_XI50/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI4/MM6 N_XI50/XI4/NET35_XI50/XI4/MM6_d N_XI50/XI4/NET36_XI50/XI4/MM6_g
+ N_VSS_XI50/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI4/MM7 N_XI50/XI4/NET36_XI50/XI4/MM7_d N_XI50/XI4/NET35_XI50/XI4/MM7_g
+ N_VSS_XI50/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI4/MM8 N_XI50/XI4/NET35_XI50/XI4/MM8_d N_WL<97>_XI50/XI4/MM8_g
+ N_BLN<11>_XI50/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI4/MM5 N_XI50/XI4/NET34_XI50/XI4/MM5_d N_XI50/XI4/NET33_XI50/XI4/MM5_g
+ N_VDD_XI50/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI4/MM4 N_XI50/XI4/NET33_XI50/XI4/MM4_d N_XI50/XI4/NET34_XI50/XI4/MM4_g
+ N_VDD_XI50/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI4/MM10 N_XI50/XI4/NET35_XI50/XI4/MM10_d N_XI50/XI4/NET36_XI50/XI4/MM10_g
+ N_VDD_XI50/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI4/MM11 N_XI50/XI4/NET36_XI50/XI4/MM11_d N_XI50/XI4/NET35_XI50/XI4/MM11_g
+ N_VDD_XI50/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI5/MM2 N_XI50/XI5/NET34_XI50/XI5/MM2_d N_XI50/XI5/NET33_XI50/XI5/MM2_g
+ N_VSS_XI50/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI5/MM3 N_XI50/XI5/NET33_XI50/XI5/MM3_d N_WL<96>_XI50/XI5/MM3_g
+ N_BLN<10>_XI50/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI5/MM0 N_XI50/XI5/NET34_XI50/XI5/MM0_d N_WL<96>_XI50/XI5/MM0_g
+ N_BL<10>_XI50/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI5/MM1 N_XI50/XI5/NET33_XI50/XI5/MM1_d N_XI50/XI5/NET34_XI50/XI5/MM1_g
+ N_VSS_XI50/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI5/MM9 N_XI50/XI5/NET36_XI50/XI5/MM9_d N_WL<97>_XI50/XI5/MM9_g
+ N_BL<10>_XI50/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI5/MM6 N_XI50/XI5/NET35_XI50/XI5/MM6_d N_XI50/XI5/NET36_XI50/XI5/MM6_g
+ N_VSS_XI50/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI5/MM7 N_XI50/XI5/NET36_XI50/XI5/MM7_d N_XI50/XI5/NET35_XI50/XI5/MM7_g
+ N_VSS_XI50/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI5/MM8 N_XI50/XI5/NET35_XI50/XI5/MM8_d N_WL<97>_XI50/XI5/MM8_g
+ N_BLN<10>_XI50/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI5/MM5 N_XI50/XI5/NET34_XI50/XI5/MM5_d N_XI50/XI5/NET33_XI50/XI5/MM5_g
+ N_VDD_XI50/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI5/MM4 N_XI50/XI5/NET33_XI50/XI5/MM4_d N_XI50/XI5/NET34_XI50/XI5/MM4_g
+ N_VDD_XI50/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI5/MM10 N_XI50/XI5/NET35_XI50/XI5/MM10_d N_XI50/XI5/NET36_XI50/XI5/MM10_g
+ N_VDD_XI50/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI5/MM11 N_XI50/XI5/NET36_XI50/XI5/MM11_d N_XI50/XI5/NET35_XI50/XI5/MM11_g
+ N_VDD_XI50/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI6/MM2 N_XI50/XI6/NET34_XI50/XI6/MM2_d N_XI50/XI6/NET33_XI50/XI6/MM2_g
+ N_VSS_XI50/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM3 N_XI50/XI6/NET33_XI50/XI6/MM3_d N_WL<96>_XI50/XI6/MM3_g
+ N_BLN<9>_XI50/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM0 N_XI50/XI6/NET34_XI50/XI6/MM0_d N_WL<96>_XI50/XI6/MM0_g
+ N_BL<9>_XI50/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM1 N_XI50/XI6/NET33_XI50/XI6/MM1_d N_XI50/XI6/NET34_XI50/XI6/MM1_g
+ N_VSS_XI50/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM9 N_XI50/XI6/NET36_XI50/XI6/MM9_d N_WL<97>_XI50/XI6/MM9_g
+ N_BL<9>_XI50/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM6 N_XI50/XI6/NET35_XI50/XI6/MM6_d N_XI50/XI6/NET36_XI50/XI6/MM6_g
+ N_VSS_XI50/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM7 N_XI50/XI6/NET36_XI50/XI6/MM7_d N_XI50/XI6/NET35_XI50/XI6/MM7_g
+ N_VSS_XI50/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM8 N_XI50/XI6/NET35_XI50/XI6/MM8_d N_WL<97>_XI50/XI6/MM8_g
+ N_BLN<9>_XI50/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI6/MM5 N_XI50/XI6/NET34_XI50/XI6/MM5_d N_XI50/XI6/NET33_XI50/XI6/MM5_g
+ N_VDD_XI50/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI6/MM4 N_XI50/XI6/NET33_XI50/XI6/MM4_d N_XI50/XI6/NET34_XI50/XI6/MM4_g
+ N_VDD_XI50/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI6/MM10 N_XI50/XI6/NET35_XI50/XI6/MM10_d N_XI50/XI6/NET36_XI50/XI6/MM10_g
+ N_VDD_XI50/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI6/MM11 N_XI50/XI6/NET36_XI50/XI6/MM11_d N_XI50/XI6/NET35_XI50/XI6/MM11_g
+ N_VDD_XI50/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI7/MM2 N_XI50/XI7/NET34_XI50/XI7/MM2_d N_XI50/XI7/NET33_XI50/XI7/MM2_g
+ N_VSS_XI50/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM3 N_XI50/XI7/NET33_XI50/XI7/MM3_d N_WL<96>_XI50/XI7/MM3_g
+ N_BLN<8>_XI50/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM0 N_XI50/XI7/NET34_XI50/XI7/MM0_d N_WL<96>_XI50/XI7/MM0_g
+ N_BL<8>_XI50/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM1 N_XI50/XI7/NET33_XI50/XI7/MM1_d N_XI50/XI7/NET34_XI50/XI7/MM1_g
+ N_VSS_XI50/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM9 N_XI50/XI7/NET36_XI50/XI7/MM9_d N_WL<97>_XI50/XI7/MM9_g
+ N_BL<8>_XI50/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM6 N_XI50/XI7/NET35_XI50/XI7/MM6_d N_XI50/XI7/NET36_XI50/XI7/MM6_g
+ N_VSS_XI50/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM7 N_XI50/XI7/NET36_XI50/XI7/MM7_d N_XI50/XI7/NET35_XI50/XI7/MM7_g
+ N_VSS_XI50/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM8 N_XI50/XI7/NET35_XI50/XI7/MM8_d N_WL<97>_XI50/XI7/MM8_g
+ N_BLN<8>_XI50/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI7/MM5 N_XI50/XI7/NET34_XI50/XI7/MM5_d N_XI50/XI7/NET33_XI50/XI7/MM5_g
+ N_VDD_XI50/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI7/MM4 N_XI50/XI7/NET33_XI50/XI7/MM4_d N_XI50/XI7/NET34_XI50/XI7/MM4_g
+ N_VDD_XI50/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI7/MM10 N_XI50/XI7/NET35_XI50/XI7/MM10_d N_XI50/XI7/NET36_XI50/XI7/MM10_g
+ N_VDD_XI50/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI7/MM11 N_XI50/XI7/NET36_XI50/XI7/MM11_d N_XI50/XI7/NET35_XI50/XI7/MM11_g
+ N_VDD_XI50/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI8/MM2 N_XI50/XI8/NET34_XI50/XI8/MM2_d N_XI50/XI8/NET33_XI50/XI8/MM2_g
+ N_VSS_XI50/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM3 N_XI50/XI8/NET33_XI50/XI8/MM3_d N_WL<96>_XI50/XI8/MM3_g
+ N_BLN<7>_XI50/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM0 N_XI50/XI8/NET34_XI50/XI8/MM0_d N_WL<96>_XI50/XI8/MM0_g
+ N_BL<7>_XI50/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM1 N_XI50/XI8/NET33_XI50/XI8/MM1_d N_XI50/XI8/NET34_XI50/XI8/MM1_g
+ N_VSS_XI50/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM9 N_XI50/XI8/NET36_XI50/XI8/MM9_d N_WL<97>_XI50/XI8/MM9_g
+ N_BL<7>_XI50/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM6 N_XI50/XI8/NET35_XI50/XI8/MM6_d N_XI50/XI8/NET36_XI50/XI8/MM6_g
+ N_VSS_XI50/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM7 N_XI50/XI8/NET36_XI50/XI8/MM7_d N_XI50/XI8/NET35_XI50/XI8/MM7_g
+ N_VSS_XI50/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM8 N_XI50/XI8/NET35_XI50/XI8/MM8_d N_WL<97>_XI50/XI8/MM8_g
+ N_BLN<7>_XI50/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI8/MM5 N_XI50/XI8/NET34_XI50/XI8/MM5_d N_XI50/XI8/NET33_XI50/XI8/MM5_g
+ N_VDD_XI50/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI8/MM4 N_XI50/XI8/NET33_XI50/XI8/MM4_d N_XI50/XI8/NET34_XI50/XI8/MM4_g
+ N_VDD_XI50/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI8/MM10 N_XI50/XI8/NET35_XI50/XI8/MM10_d N_XI50/XI8/NET36_XI50/XI8/MM10_g
+ N_VDD_XI50/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI8/MM11 N_XI50/XI8/NET36_XI50/XI8/MM11_d N_XI50/XI8/NET35_XI50/XI8/MM11_g
+ N_VDD_XI50/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI9/MM2 N_XI50/XI9/NET34_XI50/XI9/MM2_d N_XI50/XI9/NET33_XI50/XI9/MM2_g
+ N_VSS_XI50/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM3 N_XI50/XI9/NET33_XI50/XI9/MM3_d N_WL<96>_XI50/XI9/MM3_g
+ N_BLN<6>_XI50/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM0 N_XI50/XI9/NET34_XI50/XI9/MM0_d N_WL<96>_XI50/XI9/MM0_g
+ N_BL<6>_XI50/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM1 N_XI50/XI9/NET33_XI50/XI9/MM1_d N_XI50/XI9/NET34_XI50/XI9/MM1_g
+ N_VSS_XI50/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM9 N_XI50/XI9/NET36_XI50/XI9/MM9_d N_WL<97>_XI50/XI9/MM9_g
+ N_BL<6>_XI50/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM6 N_XI50/XI9/NET35_XI50/XI9/MM6_d N_XI50/XI9/NET36_XI50/XI9/MM6_g
+ N_VSS_XI50/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM7 N_XI50/XI9/NET36_XI50/XI9/MM7_d N_XI50/XI9/NET35_XI50/XI9/MM7_g
+ N_VSS_XI50/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM8 N_XI50/XI9/NET35_XI50/XI9/MM8_d N_WL<97>_XI50/XI9/MM8_g
+ N_BLN<6>_XI50/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI9/MM5 N_XI50/XI9/NET34_XI50/XI9/MM5_d N_XI50/XI9/NET33_XI50/XI9/MM5_g
+ N_VDD_XI50/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI9/MM4 N_XI50/XI9/NET33_XI50/XI9/MM4_d N_XI50/XI9/NET34_XI50/XI9/MM4_g
+ N_VDD_XI50/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI9/MM10 N_XI50/XI9/NET35_XI50/XI9/MM10_d N_XI50/XI9/NET36_XI50/XI9/MM10_g
+ N_VDD_XI50/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI9/MM11 N_XI50/XI9/NET36_XI50/XI9/MM11_d N_XI50/XI9/NET35_XI50/XI9/MM11_g
+ N_VDD_XI50/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI10/MM2 N_XI50/XI10/NET34_XI50/XI10/MM2_d
+ N_XI50/XI10/NET33_XI50/XI10/MM2_g N_VSS_XI50/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI10/MM3 N_XI50/XI10/NET33_XI50/XI10/MM3_d N_WL<96>_XI50/XI10/MM3_g
+ N_BLN<5>_XI50/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI10/MM0 N_XI50/XI10/NET34_XI50/XI10/MM0_d N_WL<96>_XI50/XI10/MM0_g
+ N_BL<5>_XI50/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI10/MM1 N_XI50/XI10/NET33_XI50/XI10/MM1_d
+ N_XI50/XI10/NET34_XI50/XI10/MM1_g N_VSS_XI50/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI10/MM9 N_XI50/XI10/NET36_XI50/XI10/MM9_d N_WL<97>_XI50/XI10/MM9_g
+ N_BL<5>_XI50/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI10/MM6 N_XI50/XI10/NET35_XI50/XI10/MM6_d
+ N_XI50/XI10/NET36_XI50/XI10/MM6_g N_VSS_XI50/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI10/MM7 N_XI50/XI10/NET36_XI50/XI10/MM7_d
+ N_XI50/XI10/NET35_XI50/XI10/MM7_g N_VSS_XI50/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI10/MM8 N_XI50/XI10/NET35_XI50/XI10/MM8_d N_WL<97>_XI50/XI10/MM8_g
+ N_BLN<5>_XI50/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI10/MM5 N_XI50/XI10/NET34_XI50/XI10/MM5_d
+ N_XI50/XI10/NET33_XI50/XI10/MM5_g N_VDD_XI50/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI10/MM4 N_XI50/XI10/NET33_XI50/XI10/MM4_d
+ N_XI50/XI10/NET34_XI50/XI10/MM4_g N_VDD_XI50/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI10/MM10 N_XI50/XI10/NET35_XI50/XI10/MM10_d
+ N_XI50/XI10/NET36_XI50/XI10/MM10_g N_VDD_XI50/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI10/MM11 N_XI50/XI10/NET36_XI50/XI10/MM11_d
+ N_XI50/XI10/NET35_XI50/XI10/MM11_g N_VDD_XI50/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI11/MM2 N_XI50/XI11/NET34_XI50/XI11/MM2_d
+ N_XI50/XI11/NET33_XI50/XI11/MM2_g N_VSS_XI50/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI11/MM3 N_XI50/XI11/NET33_XI50/XI11/MM3_d N_WL<96>_XI50/XI11/MM3_g
+ N_BLN<4>_XI50/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI11/MM0 N_XI50/XI11/NET34_XI50/XI11/MM0_d N_WL<96>_XI50/XI11/MM0_g
+ N_BL<4>_XI50/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI11/MM1 N_XI50/XI11/NET33_XI50/XI11/MM1_d
+ N_XI50/XI11/NET34_XI50/XI11/MM1_g N_VSS_XI50/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI11/MM9 N_XI50/XI11/NET36_XI50/XI11/MM9_d N_WL<97>_XI50/XI11/MM9_g
+ N_BL<4>_XI50/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI11/MM6 N_XI50/XI11/NET35_XI50/XI11/MM6_d
+ N_XI50/XI11/NET36_XI50/XI11/MM6_g N_VSS_XI50/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI11/MM7 N_XI50/XI11/NET36_XI50/XI11/MM7_d
+ N_XI50/XI11/NET35_XI50/XI11/MM7_g N_VSS_XI50/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI11/MM8 N_XI50/XI11/NET35_XI50/XI11/MM8_d N_WL<97>_XI50/XI11/MM8_g
+ N_BLN<4>_XI50/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI11/MM5 N_XI50/XI11/NET34_XI50/XI11/MM5_d
+ N_XI50/XI11/NET33_XI50/XI11/MM5_g N_VDD_XI50/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI11/MM4 N_XI50/XI11/NET33_XI50/XI11/MM4_d
+ N_XI50/XI11/NET34_XI50/XI11/MM4_g N_VDD_XI50/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI11/MM10 N_XI50/XI11/NET35_XI50/XI11/MM10_d
+ N_XI50/XI11/NET36_XI50/XI11/MM10_g N_VDD_XI50/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI11/MM11 N_XI50/XI11/NET36_XI50/XI11/MM11_d
+ N_XI50/XI11/NET35_XI50/XI11/MM11_g N_VDD_XI50/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI12/MM2 N_XI50/XI12/NET34_XI50/XI12/MM2_d
+ N_XI50/XI12/NET33_XI50/XI12/MM2_g N_VSS_XI50/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI12/MM3 N_XI50/XI12/NET33_XI50/XI12/MM3_d N_WL<96>_XI50/XI12/MM3_g
+ N_BLN<3>_XI50/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI12/MM0 N_XI50/XI12/NET34_XI50/XI12/MM0_d N_WL<96>_XI50/XI12/MM0_g
+ N_BL<3>_XI50/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI12/MM1 N_XI50/XI12/NET33_XI50/XI12/MM1_d
+ N_XI50/XI12/NET34_XI50/XI12/MM1_g N_VSS_XI50/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI12/MM9 N_XI50/XI12/NET36_XI50/XI12/MM9_d N_WL<97>_XI50/XI12/MM9_g
+ N_BL<3>_XI50/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI12/MM6 N_XI50/XI12/NET35_XI50/XI12/MM6_d
+ N_XI50/XI12/NET36_XI50/XI12/MM6_g N_VSS_XI50/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI12/MM7 N_XI50/XI12/NET36_XI50/XI12/MM7_d
+ N_XI50/XI12/NET35_XI50/XI12/MM7_g N_VSS_XI50/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI12/MM8 N_XI50/XI12/NET35_XI50/XI12/MM8_d N_WL<97>_XI50/XI12/MM8_g
+ N_BLN<3>_XI50/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI12/MM5 N_XI50/XI12/NET34_XI50/XI12/MM5_d
+ N_XI50/XI12/NET33_XI50/XI12/MM5_g N_VDD_XI50/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI12/MM4 N_XI50/XI12/NET33_XI50/XI12/MM4_d
+ N_XI50/XI12/NET34_XI50/XI12/MM4_g N_VDD_XI50/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI12/MM10 N_XI50/XI12/NET35_XI50/XI12/MM10_d
+ N_XI50/XI12/NET36_XI50/XI12/MM10_g N_VDD_XI50/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI12/MM11 N_XI50/XI12/NET36_XI50/XI12/MM11_d
+ N_XI50/XI12/NET35_XI50/XI12/MM11_g N_VDD_XI50/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI13/MM2 N_XI50/XI13/NET34_XI50/XI13/MM2_d
+ N_XI50/XI13/NET33_XI50/XI13/MM2_g N_VSS_XI50/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI13/MM3 N_XI50/XI13/NET33_XI50/XI13/MM3_d N_WL<96>_XI50/XI13/MM3_g
+ N_BLN<2>_XI50/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI13/MM0 N_XI50/XI13/NET34_XI50/XI13/MM0_d N_WL<96>_XI50/XI13/MM0_g
+ N_BL<2>_XI50/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI13/MM1 N_XI50/XI13/NET33_XI50/XI13/MM1_d
+ N_XI50/XI13/NET34_XI50/XI13/MM1_g N_VSS_XI50/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI13/MM9 N_XI50/XI13/NET36_XI50/XI13/MM9_d N_WL<97>_XI50/XI13/MM9_g
+ N_BL<2>_XI50/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI13/MM6 N_XI50/XI13/NET35_XI50/XI13/MM6_d
+ N_XI50/XI13/NET36_XI50/XI13/MM6_g N_VSS_XI50/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI13/MM7 N_XI50/XI13/NET36_XI50/XI13/MM7_d
+ N_XI50/XI13/NET35_XI50/XI13/MM7_g N_VSS_XI50/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI13/MM8 N_XI50/XI13/NET35_XI50/XI13/MM8_d N_WL<97>_XI50/XI13/MM8_g
+ N_BLN<2>_XI50/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI13/MM5 N_XI50/XI13/NET34_XI50/XI13/MM5_d
+ N_XI50/XI13/NET33_XI50/XI13/MM5_g N_VDD_XI50/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI13/MM4 N_XI50/XI13/NET33_XI50/XI13/MM4_d
+ N_XI50/XI13/NET34_XI50/XI13/MM4_g N_VDD_XI50/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI13/MM10 N_XI50/XI13/NET35_XI50/XI13/MM10_d
+ N_XI50/XI13/NET36_XI50/XI13/MM10_g N_VDD_XI50/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI13/MM11 N_XI50/XI13/NET36_XI50/XI13/MM11_d
+ N_XI50/XI13/NET35_XI50/XI13/MM11_g N_VDD_XI50/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI14/MM2 N_XI50/XI14/NET34_XI50/XI14/MM2_d
+ N_XI50/XI14/NET33_XI50/XI14/MM2_g N_VSS_XI50/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI14/MM3 N_XI50/XI14/NET33_XI50/XI14/MM3_d N_WL<96>_XI50/XI14/MM3_g
+ N_BLN<1>_XI50/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI14/MM0 N_XI50/XI14/NET34_XI50/XI14/MM0_d N_WL<96>_XI50/XI14/MM0_g
+ N_BL<1>_XI50/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI14/MM1 N_XI50/XI14/NET33_XI50/XI14/MM1_d
+ N_XI50/XI14/NET34_XI50/XI14/MM1_g N_VSS_XI50/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI14/MM9 N_XI50/XI14/NET36_XI50/XI14/MM9_d N_WL<97>_XI50/XI14/MM9_g
+ N_BL<1>_XI50/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI14/MM6 N_XI50/XI14/NET35_XI50/XI14/MM6_d
+ N_XI50/XI14/NET36_XI50/XI14/MM6_g N_VSS_XI50/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI14/MM7 N_XI50/XI14/NET36_XI50/XI14/MM7_d
+ N_XI50/XI14/NET35_XI50/XI14/MM7_g N_VSS_XI50/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI14/MM8 N_XI50/XI14/NET35_XI50/XI14/MM8_d N_WL<97>_XI50/XI14/MM8_g
+ N_BLN<1>_XI50/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI14/MM5 N_XI50/XI14/NET34_XI50/XI14/MM5_d
+ N_XI50/XI14/NET33_XI50/XI14/MM5_g N_VDD_XI50/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI14/MM4 N_XI50/XI14/NET33_XI50/XI14/MM4_d
+ N_XI50/XI14/NET34_XI50/XI14/MM4_g N_VDD_XI50/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI14/MM10 N_XI50/XI14/NET35_XI50/XI14/MM10_d
+ N_XI50/XI14/NET36_XI50/XI14/MM10_g N_VDD_XI50/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI14/MM11 N_XI50/XI14/NET36_XI50/XI14/MM11_d
+ N_XI50/XI14/NET35_XI50/XI14/MM11_g N_VDD_XI50/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI15/MM2 N_XI50/XI15/NET34_XI50/XI15/MM2_d
+ N_XI50/XI15/NET33_XI50/XI15/MM2_g N_VSS_XI50/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI15/MM3 N_XI50/XI15/NET33_XI50/XI15/MM3_d N_WL<96>_XI50/XI15/MM3_g
+ N_BLN<0>_XI50/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI15/MM0 N_XI50/XI15/NET34_XI50/XI15/MM0_d N_WL<96>_XI50/XI15/MM0_g
+ N_BL<0>_XI50/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI15/MM1 N_XI50/XI15/NET33_XI50/XI15/MM1_d
+ N_XI50/XI15/NET34_XI50/XI15/MM1_g N_VSS_XI50/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI15/MM9 N_XI50/XI15/NET36_XI50/XI15/MM9_d N_WL<97>_XI50/XI15/MM9_g
+ N_BL<0>_XI50/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI15/MM6 N_XI50/XI15/NET35_XI50/XI15/MM6_d
+ N_XI50/XI15/NET36_XI50/XI15/MM6_g N_VSS_XI50/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI15/MM7 N_XI50/XI15/NET36_XI50/XI15/MM7_d
+ N_XI50/XI15/NET35_XI50/XI15/MM7_g N_VSS_XI50/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI50/XI15/MM8 N_XI50/XI15/NET35_XI50/XI15/MM8_d N_WL<97>_XI50/XI15/MM8_g
+ N_BLN<0>_XI50/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI50/XI15/MM5 N_XI50/XI15/NET34_XI50/XI15/MM5_d
+ N_XI50/XI15/NET33_XI50/XI15/MM5_g N_VDD_XI50/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI15/MM4 N_XI50/XI15/NET33_XI50/XI15/MM4_d
+ N_XI50/XI15/NET34_XI50/XI15/MM4_g N_VDD_XI50/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI15/MM10 N_XI50/XI15/NET35_XI50/XI15/MM10_d
+ N_XI50/XI15/NET36_XI50/XI15/MM10_g N_VDD_XI50/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI50/XI15/MM11 N_XI50/XI15/NET36_XI50/XI15/MM11_d
+ N_XI50/XI15/NET35_XI50/XI15/MM11_g N_VDD_XI50/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI0/MM2 N_XI51/XI0/NET34_XI51/XI0/MM2_d N_XI51/XI0/NET33_XI51/XI0/MM2_g
+ N_VSS_XI51/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI0/MM3 N_XI51/XI0/NET33_XI51/XI0/MM3_d N_WL<98>_XI51/XI0/MM3_g
+ N_BLN<15>_XI51/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI0/MM0 N_XI51/XI0/NET34_XI51/XI0/MM0_d N_WL<98>_XI51/XI0/MM0_g
+ N_BL<15>_XI51/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI0/MM1 N_XI51/XI0/NET33_XI51/XI0/MM1_d N_XI51/XI0/NET34_XI51/XI0/MM1_g
+ N_VSS_XI51/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI0/MM9 N_XI51/XI0/NET36_XI51/XI0/MM9_d N_WL<99>_XI51/XI0/MM9_g
+ N_BL<15>_XI51/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI0/MM6 N_XI51/XI0/NET35_XI51/XI0/MM6_d N_XI51/XI0/NET36_XI51/XI0/MM6_g
+ N_VSS_XI51/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI0/MM7 N_XI51/XI0/NET36_XI51/XI0/MM7_d N_XI51/XI0/NET35_XI51/XI0/MM7_g
+ N_VSS_XI51/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI0/MM8 N_XI51/XI0/NET35_XI51/XI0/MM8_d N_WL<99>_XI51/XI0/MM8_g
+ N_BLN<15>_XI51/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI0/MM5 N_XI51/XI0/NET34_XI51/XI0/MM5_d N_XI51/XI0/NET33_XI51/XI0/MM5_g
+ N_VDD_XI51/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI0/MM4 N_XI51/XI0/NET33_XI51/XI0/MM4_d N_XI51/XI0/NET34_XI51/XI0/MM4_g
+ N_VDD_XI51/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI0/MM10 N_XI51/XI0/NET35_XI51/XI0/MM10_d N_XI51/XI0/NET36_XI51/XI0/MM10_g
+ N_VDD_XI51/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI0/MM11 N_XI51/XI0/NET36_XI51/XI0/MM11_d N_XI51/XI0/NET35_XI51/XI0/MM11_g
+ N_VDD_XI51/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI1/MM2 N_XI51/XI1/NET34_XI51/XI1/MM2_d N_XI51/XI1/NET33_XI51/XI1/MM2_g
+ N_VSS_XI51/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI1/MM3 N_XI51/XI1/NET33_XI51/XI1/MM3_d N_WL<98>_XI51/XI1/MM3_g
+ N_BLN<14>_XI51/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI1/MM0 N_XI51/XI1/NET34_XI51/XI1/MM0_d N_WL<98>_XI51/XI1/MM0_g
+ N_BL<14>_XI51/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI1/MM1 N_XI51/XI1/NET33_XI51/XI1/MM1_d N_XI51/XI1/NET34_XI51/XI1/MM1_g
+ N_VSS_XI51/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI1/MM9 N_XI51/XI1/NET36_XI51/XI1/MM9_d N_WL<99>_XI51/XI1/MM9_g
+ N_BL<14>_XI51/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI1/MM6 N_XI51/XI1/NET35_XI51/XI1/MM6_d N_XI51/XI1/NET36_XI51/XI1/MM6_g
+ N_VSS_XI51/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI1/MM7 N_XI51/XI1/NET36_XI51/XI1/MM7_d N_XI51/XI1/NET35_XI51/XI1/MM7_g
+ N_VSS_XI51/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI1/MM8 N_XI51/XI1/NET35_XI51/XI1/MM8_d N_WL<99>_XI51/XI1/MM8_g
+ N_BLN<14>_XI51/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI1/MM5 N_XI51/XI1/NET34_XI51/XI1/MM5_d N_XI51/XI1/NET33_XI51/XI1/MM5_g
+ N_VDD_XI51/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI1/MM4 N_XI51/XI1/NET33_XI51/XI1/MM4_d N_XI51/XI1/NET34_XI51/XI1/MM4_g
+ N_VDD_XI51/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI1/MM10 N_XI51/XI1/NET35_XI51/XI1/MM10_d N_XI51/XI1/NET36_XI51/XI1/MM10_g
+ N_VDD_XI51/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI1/MM11 N_XI51/XI1/NET36_XI51/XI1/MM11_d N_XI51/XI1/NET35_XI51/XI1/MM11_g
+ N_VDD_XI51/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI2/MM2 N_XI51/XI2/NET34_XI51/XI2/MM2_d N_XI51/XI2/NET33_XI51/XI2/MM2_g
+ N_VSS_XI51/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI2/MM3 N_XI51/XI2/NET33_XI51/XI2/MM3_d N_WL<98>_XI51/XI2/MM3_g
+ N_BLN<13>_XI51/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI2/MM0 N_XI51/XI2/NET34_XI51/XI2/MM0_d N_WL<98>_XI51/XI2/MM0_g
+ N_BL<13>_XI51/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI2/MM1 N_XI51/XI2/NET33_XI51/XI2/MM1_d N_XI51/XI2/NET34_XI51/XI2/MM1_g
+ N_VSS_XI51/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI2/MM9 N_XI51/XI2/NET36_XI51/XI2/MM9_d N_WL<99>_XI51/XI2/MM9_g
+ N_BL<13>_XI51/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI2/MM6 N_XI51/XI2/NET35_XI51/XI2/MM6_d N_XI51/XI2/NET36_XI51/XI2/MM6_g
+ N_VSS_XI51/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI2/MM7 N_XI51/XI2/NET36_XI51/XI2/MM7_d N_XI51/XI2/NET35_XI51/XI2/MM7_g
+ N_VSS_XI51/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI2/MM8 N_XI51/XI2/NET35_XI51/XI2/MM8_d N_WL<99>_XI51/XI2/MM8_g
+ N_BLN<13>_XI51/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI2/MM5 N_XI51/XI2/NET34_XI51/XI2/MM5_d N_XI51/XI2/NET33_XI51/XI2/MM5_g
+ N_VDD_XI51/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI2/MM4 N_XI51/XI2/NET33_XI51/XI2/MM4_d N_XI51/XI2/NET34_XI51/XI2/MM4_g
+ N_VDD_XI51/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI2/MM10 N_XI51/XI2/NET35_XI51/XI2/MM10_d N_XI51/XI2/NET36_XI51/XI2/MM10_g
+ N_VDD_XI51/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI2/MM11 N_XI51/XI2/NET36_XI51/XI2/MM11_d N_XI51/XI2/NET35_XI51/XI2/MM11_g
+ N_VDD_XI51/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI3/MM2 N_XI51/XI3/NET34_XI51/XI3/MM2_d N_XI51/XI3/NET33_XI51/XI3/MM2_g
+ N_VSS_XI51/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI3/MM3 N_XI51/XI3/NET33_XI51/XI3/MM3_d N_WL<98>_XI51/XI3/MM3_g
+ N_BLN<12>_XI51/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI3/MM0 N_XI51/XI3/NET34_XI51/XI3/MM0_d N_WL<98>_XI51/XI3/MM0_g
+ N_BL<12>_XI51/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI3/MM1 N_XI51/XI3/NET33_XI51/XI3/MM1_d N_XI51/XI3/NET34_XI51/XI3/MM1_g
+ N_VSS_XI51/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI3/MM9 N_XI51/XI3/NET36_XI51/XI3/MM9_d N_WL<99>_XI51/XI3/MM9_g
+ N_BL<12>_XI51/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI3/MM6 N_XI51/XI3/NET35_XI51/XI3/MM6_d N_XI51/XI3/NET36_XI51/XI3/MM6_g
+ N_VSS_XI51/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI3/MM7 N_XI51/XI3/NET36_XI51/XI3/MM7_d N_XI51/XI3/NET35_XI51/XI3/MM7_g
+ N_VSS_XI51/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI3/MM8 N_XI51/XI3/NET35_XI51/XI3/MM8_d N_WL<99>_XI51/XI3/MM8_g
+ N_BLN<12>_XI51/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI3/MM5 N_XI51/XI3/NET34_XI51/XI3/MM5_d N_XI51/XI3/NET33_XI51/XI3/MM5_g
+ N_VDD_XI51/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI3/MM4 N_XI51/XI3/NET33_XI51/XI3/MM4_d N_XI51/XI3/NET34_XI51/XI3/MM4_g
+ N_VDD_XI51/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI3/MM10 N_XI51/XI3/NET35_XI51/XI3/MM10_d N_XI51/XI3/NET36_XI51/XI3/MM10_g
+ N_VDD_XI51/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI3/MM11 N_XI51/XI3/NET36_XI51/XI3/MM11_d N_XI51/XI3/NET35_XI51/XI3/MM11_g
+ N_VDD_XI51/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI4/MM2 N_XI51/XI4/NET34_XI51/XI4/MM2_d N_XI51/XI4/NET33_XI51/XI4/MM2_g
+ N_VSS_XI51/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI4/MM3 N_XI51/XI4/NET33_XI51/XI4/MM3_d N_WL<98>_XI51/XI4/MM3_g
+ N_BLN<11>_XI51/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI4/MM0 N_XI51/XI4/NET34_XI51/XI4/MM0_d N_WL<98>_XI51/XI4/MM0_g
+ N_BL<11>_XI51/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI4/MM1 N_XI51/XI4/NET33_XI51/XI4/MM1_d N_XI51/XI4/NET34_XI51/XI4/MM1_g
+ N_VSS_XI51/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI4/MM9 N_XI51/XI4/NET36_XI51/XI4/MM9_d N_WL<99>_XI51/XI4/MM9_g
+ N_BL<11>_XI51/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI4/MM6 N_XI51/XI4/NET35_XI51/XI4/MM6_d N_XI51/XI4/NET36_XI51/XI4/MM6_g
+ N_VSS_XI51/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI4/MM7 N_XI51/XI4/NET36_XI51/XI4/MM7_d N_XI51/XI4/NET35_XI51/XI4/MM7_g
+ N_VSS_XI51/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI4/MM8 N_XI51/XI4/NET35_XI51/XI4/MM8_d N_WL<99>_XI51/XI4/MM8_g
+ N_BLN<11>_XI51/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI4/MM5 N_XI51/XI4/NET34_XI51/XI4/MM5_d N_XI51/XI4/NET33_XI51/XI4/MM5_g
+ N_VDD_XI51/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI4/MM4 N_XI51/XI4/NET33_XI51/XI4/MM4_d N_XI51/XI4/NET34_XI51/XI4/MM4_g
+ N_VDD_XI51/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI4/MM10 N_XI51/XI4/NET35_XI51/XI4/MM10_d N_XI51/XI4/NET36_XI51/XI4/MM10_g
+ N_VDD_XI51/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI4/MM11 N_XI51/XI4/NET36_XI51/XI4/MM11_d N_XI51/XI4/NET35_XI51/XI4/MM11_g
+ N_VDD_XI51/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI5/MM2 N_XI51/XI5/NET34_XI51/XI5/MM2_d N_XI51/XI5/NET33_XI51/XI5/MM2_g
+ N_VSS_XI51/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI5/MM3 N_XI51/XI5/NET33_XI51/XI5/MM3_d N_WL<98>_XI51/XI5/MM3_g
+ N_BLN<10>_XI51/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI5/MM0 N_XI51/XI5/NET34_XI51/XI5/MM0_d N_WL<98>_XI51/XI5/MM0_g
+ N_BL<10>_XI51/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI5/MM1 N_XI51/XI5/NET33_XI51/XI5/MM1_d N_XI51/XI5/NET34_XI51/XI5/MM1_g
+ N_VSS_XI51/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI5/MM9 N_XI51/XI5/NET36_XI51/XI5/MM9_d N_WL<99>_XI51/XI5/MM9_g
+ N_BL<10>_XI51/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI5/MM6 N_XI51/XI5/NET35_XI51/XI5/MM6_d N_XI51/XI5/NET36_XI51/XI5/MM6_g
+ N_VSS_XI51/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI5/MM7 N_XI51/XI5/NET36_XI51/XI5/MM7_d N_XI51/XI5/NET35_XI51/XI5/MM7_g
+ N_VSS_XI51/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI5/MM8 N_XI51/XI5/NET35_XI51/XI5/MM8_d N_WL<99>_XI51/XI5/MM8_g
+ N_BLN<10>_XI51/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI5/MM5 N_XI51/XI5/NET34_XI51/XI5/MM5_d N_XI51/XI5/NET33_XI51/XI5/MM5_g
+ N_VDD_XI51/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI5/MM4 N_XI51/XI5/NET33_XI51/XI5/MM4_d N_XI51/XI5/NET34_XI51/XI5/MM4_g
+ N_VDD_XI51/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI5/MM10 N_XI51/XI5/NET35_XI51/XI5/MM10_d N_XI51/XI5/NET36_XI51/XI5/MM10_g
+ N_VDD_XI51/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI5/MM11 N_XI51/XI5/NET36_XI51/XI5/MM11_d N_XI51/XI5/NET35_XI51/XI5/MM11_g
+ N_VDD_XI51/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI6/MM2 N_XI51/XI6/NET34_XI51/XI6/MM2_d N_XI51/XI6/NET33_XI51/XI6/MM2_g
+ N_VSS_XI51/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM3 N_XI51/XI6/NET33_XI51/XI6/MM3_d N_WL<98>_XI51/XI6/MM3_g
+ N_BLN<9>_XI51/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM0 N_XI51/XI6/NET34_XI51/XI6/MM0_d N_WL<98>_XI51/XI6/MM0_g
+ N_BL<9>_XI51/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM1 N_XI51/XI6/NET33_XI51/XI6/MM1_d N_XI51/XI6/NET34_XI51/XI6/MM1_g
+ N_VSS_XI51/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM9 N_XI51/XI6/NET36_XI51/XI6/MM9_d N_WL<99>_XI51/XI6/MM9_g
+ N_BL<9>_XI51/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM6 N_XI51/XI6/NET35_XI51/XI6/MM6_d N_XI51/XI6/NET36_XI51/XI6/MM6_g
+ N_VSS_XI51/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM7 N_XI51/XI6/NET36_XI51/XI6/MM7_d N_XI51/XI6/NET35_XI51/XI6/MM7_g
+ N_VSS_XI51/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM8 N_XI51/XI6/NET35_XI51/XI6/MM8_d N_WL<99>_XI51/XI6/MM8_g
+ N_BLN<9>_XI51/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI6/MM5 N_XI51/XI6/NET34_XI51/XI6/MM5_d N_XI51/XI6/NET33_XI51/XI6/MM5_g
+ N_VDD_XI51/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI6/MM4 N_XI51/XI6/NET33_XI51/XI6/MM4_d N_XI51/XI6/NET34_XI51/XI6/MM4_g
+ N_VDD_XI51/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI6/MM10 N_XI51/XI6/NET35_XI51/XI6/MM10_d N_XI51/XI6/NET36_XI51/XI6/MM10_g
+ N_VDD_XI51/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI6/MM11 N_XI51/XI6/NET36_XI51/XI6/MM11_d N_XI51/XI6/NET35_XI51/XI6/MM11_g
+ N_VDD_XI51/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI7/MM2 N_XI51/XI7/NET34_XI51/XI7/MM2_d N_XI51/XI7/NET33_XI51/XI7/MM2_g
+ N_VSS_XI51/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM3 N_XI51/XI7/NET33_XI51/XI7/MM3_d N_WL<98>_XI51/XI7/MM3_g
+ N_BLN<8>_XI51/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM0 N_XI51/XI7/NET34_XI51/XI7/MM0_d N_WL<98>_XI51/XI7/MM0_g
+ N_BL<8>_XI51/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM1 N_XI51/XI7/NET33_XI51/XI7/MM1_d N_XI51/XI7/NET34_XI51/XI7/MM1_g
+ N_VSS_XI51/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM9 N_XI51/XI7/NET36_XI51/XI7/MM9_d N_WL<99>_XI51/XI7/MM9_g
+ N_BL<8>_XI51/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM6 N_XI51/XI7/NET35_XI51/XI7/MM6_d N_XI51/XI7/NET36_XI51/XI7/MM6_g
+ N_VSS_XI51/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM7 N_XI51/XI7/NET36_XI51/XI7/MM7_d N_XI51/XI7/NET35_XI51/XI7/MM7_g
+ N_VSS_XI51/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM8 N_XI51/XI7/NET35_XI51/XI7/MM8_d N_WL<99>_XI51/XI7/MM8_g
+ N_BLN<8>_XI51/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI7/MM5 N_XI51/XI7/NET34_XI51/XI7/MM5_d N_XI51/XI7/NET33_XI51/XI7/MM5_g
+ N_VDD_XI51/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI7/MM4 N_XI51/XI7/NET33_XI51/XI7/MM4_d N_XI51/XI7/NET34_XI51/XI7/MM4_g
+ N_VDD_XI51/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI7/MM10 N_XI51/XI7/NET35_XI51/XI7/MM10_d N_XI51/XI7/NET36_XI51/XI7/MM10_g
+ N_VDD_XI51/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI7/MM11 N_XI51/XI7/NET36_XI51/XI7/MM11_d N_XI51/XI7/NET35_XI51/XI7/MM11_g
+ N_VDD_XI51/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI8/MM2 N_XI51/XI8/NET34_XI51/XI8/MM2_d N_XI51/XI8/NET33_XI51/XI8/MM2_g
+ N_VSS_XI51/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM3 N_XI51/XI8/NET33_XI51/XI8/MM3_d N_WL<98>_XI51/XI8/MM3_g
+ N_BLN<7>_XI51/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM0 N_XI51/XI8/NET34_XI51/XI8/MM0_d N_WL<98>_XI51/XI8/MM0_g
+ N_BL<7>_XI51/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM1 N_XI51/XI8/NET33_XI51/XI8/MM1_d N_XI51/XI8/NET34_XI51/XI8/MM1_g
+ N_VSS_XI51/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM9 N_XI51/XI8/NET36_XI51/XI8/MM9_d N_WL<99>_XI51/XI8/MM9_g
+ N_BL<7>_XI51/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM6 N_XI51/XI8/NET35_XI51/XI8/MM6_d N_XI51/XI8/NET36_XI51/XI8/MM6_g
+ N_VSS_XI51/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM7 N_XI51/XI8/NET36_XI51/XI8/MM7_d N_XI51/XI8/NET35_XI51/XI8/MM7_g
+ N_VSS_XI51/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM8 N_XI51/XI8/NET35_XI51/XI8/MM8_d N_WL<99>_XI51/XI8/MM8_g
+ N_BLN<7>_XI51/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI8/MM5 N_XI51/XI8/NET34_XI51/XI8/MM5_d N_XI51/XI8/NET33_XI51/XI8/MM5_g
+ N_VDD_XI51/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI8/MM4 N_XI51/XI8/NET33_XI51/XI8/MM4_d N_XI51/XI8/NET34_XI51/XI8/MM4_g
+ N_VDD_XI51/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI8/MM10 N_XI51/XI8/NET35_XI51/XI8/MM10_d N_XI51/XI8/NET36_XI51/XI8/MM10_g
+ N_VDD_XI51/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI8/MM11 N_XI51/XI8/NET36_XI51/XI8/MM11_d N_XI51/XI8/NET35_XI51/XI8/MM11_g
+ N_VDD_XI51/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI9/MM2 N_XI51/XI9/NET34_XI51/XI9/MM2_d N_XI51/XI9/NET33_XI51/XI9/MM2_g
+ N_VSS_XI51/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM3 N_XI51/XI9/NET33_XI51/XI9/MM3_d N_WL<98>_XI51/XI9/MM3_g
+ N_BLN<6>_XI51/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM0 N_XI51/XI9/NET34_XI51/XI9/MM0_d N_WL<98>_XI51/XI9/MM0_g
+ N_BL<6>_XI51/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM1 N_XI51/XI9/NET33_XI51/XI9/MM1_d N_XI51/XI9/NET34_XI51/XI9/MM1_g
+ N_VSS_XI51/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM9 N_XI51/XI9/NET36_XI51/XI9/MM9_d N_WL<99>_XI51/XI9/MM9_g
+ N_BL<6>_XI51/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM6 N_XI51/XI9/NET35_XI51/XI9/MM6_d N_XI51/XI9/NET36_XI51/XI9/MM6_g
+ N_VSS_XI51/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM7 N_XI51/XI9/NET36_XI51/XI9/MM7_d N_XI51/XI9/NET35_XI51/XI9/MM7_g
+ N_VSS_XI51/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM8 N_XI51/XI9/NET35_XI51/XI9/MM8_d N_WL<99>_XI51/XI9/MM8_g
+ N_BLN<6>_XI51/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI9/MM5 N_XI51/XI9/NET34_XI51/XI9/MM5_d N_XI51/XI9/NET33_XI51/XI9/MM5_g
+ N_VDD_XI51/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI9/MM4 N_XI51/XI9/NET33_XI51/XI9/MM4_d N_XI51/XI9/NET34_XI51/XI9/MM4_g
+ N_VDD_XI51/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI9/MM10 N_XI51/XI9/NET35_XI51/XI9/MM10_d N_XI51/XI9/NET36_XI51/XI9/MM10_g
+ N_VDD_XI51/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI9/MM11 N_XI51/XI9/NET36_XI51/XI9/MM11_d N_XI51/XI9/NET35_XI51/XI9/MM11_g
+ N_VDD_XI51/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI10/MM2 N_XI51/XI10/NET34_XI51/XI10/MM2_d
+ N_XI51/XI10/NET33_XI51/XI10/MM2_g N_VSS_XI51/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI10/MM3 N_XI51/XI10/NET33_XI51/XI10/MM3_d N_WL<98>_XI51/XI10/MM3_g
+ N_BLN<5>_XI51/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI10/MM0 N_XI51/XI10/NET34_XI51/XI10/MM0_d N_WL<98>_XI51/XI10/MM0_g
+ N_BL<5>_XI51/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI10/MM1 N_XI51/XI10/NET33_XI51/XI10/MM1_d
+ N_XI51/XI10/NET34_XI51/XI10/MM1_g N_VSS_XI51/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI10/MM9 N_XI51/XI10/NET36_XI51/XI10/MM9_d N_WL<99>_XI51/XI10/MM9_g
+ N_BL<5>_XI51/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI10/MM6 N_XI51/XI10/NET35_XI51/XI10/MM6_d
+ N_XI51/XI10/NET36_XI51/XI10/MM6_g N_VSS_XI51/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI10/MM7 N_XI51/XI10/NET36_XI51/XI10/MM7_d
+ N_XI51/XI10/NET35_XI51/XI10/MM7_g N_VSS_XI51/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI10/MM8 N_XI51/XI10/NET35_XI51/XI10/MM8_d N_WL<99>_XI51/XI10/MM8_g
+ N_BLN<5>_XI51/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI10/MM5 N_XI51/XI10/NET34_XI51/XI10/MM5_d
+ N_XI51/XI10/NET33_XI51/XI10/MM5_g N_VDD_XI51/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI10/MM4 N_XI51/XI10/NET33_XI51/XI10/MM4_d
+ N_XI51/XI10/NET34_XI51/XI10/MM4_g N_VDD_XI51/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI10/MM10 N_XI51/XI10/NET35_XI51/XI10/MM10_d
+ N_XI51/XI10/NET36_XI51/XI10/MM10_g N_VDD_XI51/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI10/MM11 N_XI51/XI10/NET36_XI51/XI10/MM11_d
+ N_XI51/XI10/NET35_XI51/XI10/MM11_g N_VDD_XI51/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI11/MM2 N_XI51/XI11/NET34_XI51/XI11/MM2_d
+ N_XI51/XI11/NET33_XI51/XI11/MM2_g N_VSS_XI51/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI11/MM3 N_XI51/XI11/NET33_XI51/XI11/MM3_d N_WL<98>_XI51/XI11/MM3_g
+ N_BLN<4>_XI51/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI11/MM0 N_XI51/XI11/NET34_XI51/XI11/MM0_d N_WL<98>_XI51/XI11/MM0_g
+ N_BL<4>_XI51/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI11/MM1 N_XI51/XI11/NET33_XI51/XI11/MM1_d
+ N_XI51/XI11/NET34_XI51/XI11/MM1_g N_VSS_XI51/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI11/MM9 N_XI51/XI11/NET36_XI51/XI11/MM9_d N_WL<99>_XI51/XI11/MM9_g
+ N_BL<4>_XI51/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI11/MM6 N_XI51/XI11/NET35_XI51/XI11/MM6_d
+ N_XI51/XI11/NET36_XI51/XI11/MM6_g N_VSS_XI51/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI11/MM7 N_XI51/XI11/NET36_XI51/XI11/MM7_d
+ N_XI51/XI11/NET35_XI51/XI11/MM7_g N_VSS_XI51/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI11/MM8 N_XI51/XI11/NET35_XI51/XI11/MM8_d N_WL<99>_XI51/XI11/MM8_g
+ N_BLN<4>_XI51/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI11/MM5 N_XI51/XI11/NET34_XI51/XI11/MM5_d
+ N_XI51/XI11/NET33_XI51/XI11/MM5_g N_VDD_XI51/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI11/MM4 N_XI51/XI11/NET33_XI51/XI11/MM4_d
+ N_XI51/XI11/NET34_XI51/XI11/MM4_g N_VDD_XI51/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI11/MM10 N_XI51/XI11/NET35_XI51/XI11/MM10_d
+ N_XI51/XI11/NET36_XI51/XI11/MM10_g N_VDD_XI51/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI11/MM11 N_XI51/XI11/NET36_XI51/XI11/MM11_d
+ N_XI51/XI11/NET35_XI51/XI11/MM11_g N_VDD_XI51/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI12/MM2 N_XI51/XI12/NET34_XI51/XI12/MM2_d
+ N_XI51/XI12/NET33_XI51/XI12/MM2_g N_VSS_XI51/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI12/MM3 N_XI51/XI12/NET33_XI51/XI12/MM3_d N_WL<98>_XI51/XI12/MM3_g
+ N_BLN<3>_XI51/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI12/MM0 N_XI51/XI12/NET34_XI51/XI12/MM0_d N_WL<98>_XI51/XI12/MM0_g
+ N_BL<3>_XI51/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI12/MM1 N_XI51/XI12/NET33_XI51/XI12/MM1_d
+ N_XI51/XI12/NET34_XI51/XI12/MM1_g N_VSS_XI51/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI12/MM9 N_XI51/XI12/NET36_XI51/XI12/MM9_d N_WL<99>_XI51/XI12/MM9_g
+ N_BL<3>_XI51/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI12/MM6 N_XI51/XI12/NET35_XI51/XI12/MM6_d
+ N_XI51/XI12/NET36_XI51/XI12/MM6_g N_VSS_XI51/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI12/MM7 N_XI51/XI12/NET36_XI51/XI12/MM7_d
+ N_XI51/XI12/NET35_XI51/XI12/MM7_g N_VSS_XI51/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI12/MM8 N_XI51/XI12/NET35_XI51/XI12/MM8_d N_WL<99>_XI51/XI12/MM8_g
+ N_BLN<3>_XI51/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI12/MM5 N_XI51/XI12/NET34_XI51/XI12/MM5_d
+ N_XI51/XI12/NET33_XI51/XI12/MM5_g N_VDD_XI51/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI12/MM4 N_XI51/XI12/NET33_XI51/XI12/MM4_d
+ N_XI51/XI12/NET34_XI51/XI12/MM4_g N_VDD_XI51/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI12/MM10 N_XI51/XI12/NET35_XI51/XI12/MM10_d
+ N_XI51/XI12/NET36_XI51/XI12/MM10_g N_VDD_XI51/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI12/MM11 N_XI51/XI12/NET36_XI51/XI12/MM11_d
+ N_XI51/XI12/NET35_XI51/XI12/MM11_g N_VDD_XI51/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI13/MM2 N_XI51/XI13/NET34_XI51/XI13/MM2_d
+ N_XI51/XI13/NET33_XI51/XI13/MM2_g N_VSS_XI51/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI13/MM3 N_XI51/XI13/NET33_XI51/XI13/MM3_d N_WL<98>_XI51/XI13/MM3_g
+ N_BLN<2>_XI51/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI13/MM0 N_XI51/XI13/NET34_XI51/XI13/MM0_d N_WL<98>_XI51/XI13/MM0_g
+ N_BL<2>_XI51/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI13/MM1 N_XI51/XI13/NET33_XI51/XI13/MM1_d
+ N_XI51/XI13/NET34_XI51/XI13/MM1_g N_VSS_XI51/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI13/MM9 N_XI51/XI13/NET36_XI51/XI13/MM9_d N_WL<99>_XI51/XI13/MM9_g
+ N_BL<2>_XI51/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI13/MM6 N_XI51/XI13/NET35_XI51/XI13/MM6_d
+ N_XI51/XI13/NET36_XI51/XI13/MM6_g N_VSS_XI51/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI13/MM7 N_XI51/XI13/NET36_XI51/XI13/MM7_d
+ N_XI51/XI13/NET35_XI51/XI13/MM7_g N_VSS_XI51/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI13/MM8 N_XI51/XI13/NET35_XI51/XI13/MM8_d N_WL<99>_XI51/XI13/MM8_g
+ N_BLN<2>_XI51/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI13/MM5 N_XI51/XI13/NET34_XI51/XI13/MM5_d
+ N_XI51/XI13/NET33_XI51/XI13/MM5_g N_VDD_XI51/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI13/MM4 N_XI51/XI13/NET33_XI51/XI13/MM4_d
+ N_XI51/XI13/NET34_XI51/XI13/MM4_g N_VDD_XI51/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI13/MM10 N_XI51/XI13/NET35_XI51/XI13/MM10_d
+ N_XI51/XI13/NET36_XI51/XI13/MM10_g N_VDD_XI51/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI13/MM11 N_XI51/XI13/NET36_XI51/XI13/MM11_d
+ N_XI51/XI13/NET35_XI51/XI13/MM11_g N_VDD_XI51/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI14/MM2 N_XI51/XI14/NET34_XI51/XI14/MM2_d
+ N_XI51/XI14/NET33_XI51/XI14/MM2_g N_VSS_XI51/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI14/MM3 N_XI51/XI14/NET33_XI51/XI14/MM3_d N_WL<98>_XI51/XI14/MM3_g
+ N_BLN<1>_XI51/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI14/MM0 N_XI51/XI14/NET34_XI51/XI14/MM0_d N_WL<98>_XI51/XI14/MM0_g
+ N_BL<1>_XI51/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI14/MM1 N_XI51/XI14/NET33_XI51/XI14/MM1_d
+ N_XI51/XI14/NET34_XI51/XI14/MM1_g N_VSS_XI51/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI14/MM9 N_XI51/XI14/NET36_XI51/XI14/MM9_d N_WL<99>_XI51/XI14/MM9_g
+ N_BL<1>_XI51/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI14/MM6 N_XI51/XI14/NET35_XI51/XI14/MM6_d
+ N_XI51/XI14/NET36_XI51/XI14/MM6_g N_VSS_XI51/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI14/MM7 N_XI51/XI14/NET36_XI51/XI14/MM7_d
+ N_XI51/XI14/NET35_XI51/XI14/MM7_g N_VSS_XI51/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI14/MM8 N_XI51/XI14/NET35_XI51/XI14/MM8_d N_WL<99>_XI51/XI14/MM8_g
+ N_BLN<1>_XI51/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI14/MM5 N_XI51/XI14/NET34_XI51/XI14/MM5_d
+ N_XI51/XI14/NET33_XI51/XI14/MM5_g N_VDD_XI51/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI14/MM4 N_XI51/XI14/NET33_XI51/XI14/MM4_d
+ N_XI51/XI14/NET34_XI51/XI14/MM4_g N_VDD_XI51/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI14/MM10 N_XI51/XI14/NET35_XI51/XI14/MM10_d
+ N_XI51/XI14/NET36_XI51/XI14/MM10_g N_VDD_XI51/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI14/MM11 N_XI51/XI14/NET36_XI51/XI14/MM11_d
+ N_XI51/XI14/NET35_XI51/XI14/MM11_g N_VDD_XI51/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI15/MM2 N_XI51/XI15/NET34_XI51/XI15/MM2_d
+ N_XI51/XI15/NET33_XI51/XI15/MM2_g N_VSS_XI51/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI15/MM3 N_XI51/XI15/NET33_XI51/XI15/MM3_d N_WL<98>_XI51/XI15/MM3_g
+ N_BLN<0>_XI51/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI15/MM0 N_XI51/XI15/NET34_XI51/XI15/MM0_d N_WL<98>_XI51/XI15/MM0_g
+ N_BL<0>_XI51/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI15/MM1 N_XI51/XI15/NET33_XI51/XI15/MM1_d
+ N_XI51/XI15/NET34_XI51/XI15/MM1_g N_VSS_XI51/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI15/MM9 N_XI51/XI15/NET36_XI51/XI15/MM9_d N_WL<99>_XI51/XI15/MM9_g
+ N_BL<0>_XI51/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI15/MM6 N_XI51/XI15/NET35_XI51/XI15/MM6_d
+ N_XI51/XI15/NET36_XI51/XI15/MM6_g N_VSS_XI51/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI15/MM7 N_XI51/XI15/NET36_XI51/XI15/MM7_d
+ N_XI51/XI15/NET35_XI51/XI15/MM7_g N_VSS_XI51/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI51/XI15/MM8 N_XI51/XI15/NET35_XI51/XI15/MM8_d N_WL<99>_XI51/XI15/MM8_g
+ N_BLN<0>_XI51/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI51/XI15/MM5 N_XI51/XI15/NET34_XI51/XI15/MM5_d
+ N_XI51/XI15/NET33_XI51/XI15/MM5_g N_VDD_XI51/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI15/MM4 N_XI51/XI15/NET33_XI51/XI15/MM4_d
+ N_XI51/XI15/NET34_XI51/XI15/MM4_g N_VDD_XI51/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI15/MM10 N_XI51/XI15/NET35_XI51/XI15/MM10_d
+ N_XI51/XI15/NET36_XI51/XI15/MM10_g N_VDD_XI51/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI51/XI15/MM11 N_XI51/XI15/NET36_XI51/XI15/MM11_d
+ N_XI51/XI15/NET35_XI51/XI15/MM11_g N_VDD_XI51/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI0/MM2 N_XI52/XI0/NET34_XI52/XI0/MM2_d N_XI52/XI0/NET33_XI52/XI0/MM2_g
+ N_VSS_XI52/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI0/MM3 N_XI52/XI0/NET33_XI52/XI0/MM3_d N_WL<100>_XI52/XI0/MM3_g
+ N_BLN<15>_XI52/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI0/MM0 N_XI52/XI0/NET34_XI52/XI0/MM0_d N_WL<100>_XI52/XI0/MM0_g
+ N_BL<15>_XI52/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI0/MM1 N_XI52/XI0/NET33_XI52/XI0/MM1_d N_XI52/XI0/NET34_XI52/XI0/MM1_g
+ N_VSS_XI52/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI0/MM9 N_XI52/XI0/NET36_XI52/XI0/MM9_d N_WL<101>_XI52/XI0/MM9_g
+ N_BL<15>_XI52/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI0/MM6 N_XI52/XI0/NET35_XI52/XI0/MM6_d N_XI52/XI0/NET36_XI52/XI0/MM6_g
+ N_VSS_XI52/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI0/MM7 N_XI52/XI0/NET36_XI52/XI0/MM7_d N_XI52/XI0/NET35_XI52/XI0/MM7_g
+ N_VSS_XI52/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI0/MM8 N_XI52/XI0/NET35_XI52/XI0/MM8_d N_WL<101>_XI52/XI0/MM8_g
+ N_BLN<15>_XI52/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI0/MM5 N_XI52/XI0/NET34_XI52/XI0/MM5_d N_XI52/XI0/NET33_XI52/XI0/MM5_g
+ N_VDD_XI52/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI0/MM4 N_XI52/XI0/NET33_XI52/XI0/MM4_d N_XI52/XI0/NET34_XI52/XI0/MM4_g
+ N_VDD_XI52/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI0/MM10 N_XI52/XI0/NET35_XI52/XI0/MM10_d N_XI52/XI0/NET36_XI52/XI0/MM10_g
+ N_VDD_XI52/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI0/MM11 N_XI52/XI0/NET36_XI52/XI0/MM11_d N_XI52/XI0/NET35_XI52/XI0/MM11_g
+ N_VDD_XI52/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI1/MM2 N_XI52/XI1/NET34_XI52/XI1/MM2_d N_XI52/XI1/NET33_XI52/XI1/MM2_g
+ N_VSS_XI52/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI1/MM3 N_XI52/XI1/NET33_XI52/XI1/MM3_d N_WL<100>_XI52/XI1/MM3_g
+ N_BLN<14>_XI52/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI1/MM0 N_XI52/XI1/NET34_XI52/XI1/MM0_d N_WL<100>_XI52/XI1/MM0_g
+ N_BL<14>_XI52/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI1/MM1 N_XI52/XI1/NET33_XI52/XI1/MM1_d N_XI52/XI1/NET34_XI52/XI1/MM1_g
+ N_VSS_XI52/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI1/MM9 N_XI52/XI1/NET36_XI52/XI1/MM9_d N_WL<101>_XI52/XI1/MM9_g
+ N_BL<14>_XI52/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI1/MM6 N_XI52/XI1/NET35_XI52/XI1/MM6_d N_XI52/XI1/NET36_XI52/XI1/MM6_g
+ N_VSS_XI52/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI1/MM7 N_XI52/XI1/NET36_XI52/XI1/MM7_d N_XI52/XI1/NET35_XI52/XI1/MM7_g
+ N_VSS_XI52/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI1/MM8 N_XI52/XI1/NET35_XI52/XI1/MM8_d N_WL<101>_XI52/XI1/MM8_g
+ N_BLN<14>_XI52/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI1/MM5 N_XI52/XI1/NET34_XI52/XI1/MM5_d N_XI52/XI1/NET33_XI52/XI1/MM5_g
+ N_VDD_XI52/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI1/MM4 N_XI52/XI1/NET33_XI52/XI1/MM4_d N_XI52/XI1/NET34_XI52/XI1/MM4_g
+ N_VDD_XI52/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI1/MM10 N_XI52/XI1/NET35_XI52/XI1/MM10_d N_XI52/XI1/NET36_XI52/XI1/MM10_g
+ N_VDD_XI52/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI1/MM11 N_XI52/XI1/NET36_XI52/XI1/MM11_d N_XI52/XI1/NET35_XI52/XI1/MM11_g
+ N_VDD_XI52/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI2/MM2 N_XI52/XI2/NET34_XI52/XI2/MM2_d N_XI52/XI2/NET33_XI52/XI2/MM2_g
+ N_VSS_XI52/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI2/MM3 N_XI52/XI2/NET33_XI52/XI2/MM3_d N_WL<100>_XI52/XI2/MM3_g
+ N_BLN<13>_XI52/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI2/MM0 N_XI52/XI2/NET34_XI52/XI2/MM0_d N_WL<100>_XI52/XI2/MM0_g
+ N_BL<13>_XI52/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI2/MM1 N_XI52/XI2/NET33_XI52/XI2/MM1_d N_XI52/XI2/NET34_XI52/XI2/MM1_g
+ N_VSS_XI52/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI2/MM9 N_XI52/XI2/NET36_XI52/XI2/MM9_d N_WL<101>_XI52/XI2/MM9_g
+ N_BL<13>_XI52/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI2/MM6 N_XI52/XI2/NET35_XI52/XI2/MM6_d N_XI52/XI2/NET36_XI52/XI2/MM6_g
+ N_VSS_XI52/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI2/MM7 N_XI52/XI2/NET36_XI52/XI2/MM7_d N_XI52/XI2/NET35_XI52/XI2/MM7_g
+ N_VSS_XI52/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI2/MM8 N_XI52/XI2/NET35_XI52/XI2/MM8_d N_WL<101>_XI52/XI2/MM8_g
+ N_BLN<13>_XI52/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI2/MM5 N_XI52/XI2/NET34_XI52/XI2/MM5_d N_XI52/XI2/NET33_XI52/XI2/MM5_g
+ N_VDD_XI52/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI2/MM4 N_XI52/XI2/NET33_XI52/XI2/MM4_d N_XI52/XI2/NET34_XI52/XI2/MM4_g
+ N_VDD_XI52/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI2/MM10 N_XI52/XI2/NET35_XI52/XI2/MM10_d N_XI52/XI2/NET36_XI52/XI2/MM10_g
+ N_VDD_XI52/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI2/MM11 N_XI52/XI2/NET36_XI52/XI2/MM11_d N_XI52/XI2/NET35_XI52/XI2/MM11_g
+ N_VDD_XI52/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI3/MM2 N_XI52/XI3/NET34_XI52/XI3/MM2_d N_XI52/XI3/NET33_XI52/XI3/MM2_g
+ N_VSS_XI52/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI3/MM3 N_XI52/XI3/NET33_XI52/XI3/MM3_d N_WL<100>_XI52/XI3/MM3_g
+ N_BLN<12>_XI52/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI3/MM0 N_XI52/XI3/NET34_XI52/XI3/MM0_d N_WL<100>_XI52/XI3/MM0_g
+ N_BL<12>_XI52/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI3/MM1 N_XI52/XI3/NET33_XI52/XI3/MM1_d N_XI52/XI3/NET34_XI52/XI3/MM1_g
+ N_VSS_XI52/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI3/MM9 N_XI52/XI3/NET36_XI52/XI3/MM9_d N_WL<101>_XI52/XI3/MM9_g
+ N_BL<12>_XI52/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI3/MM6 N_XI52/XI3/NET35_XI52/XI3/MM6_d N_XI52/XI3/NET36_XI52/XI3/MM6_g
+ N_VSS_XI52/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI3/MM7 N_XI52/XI3/NET36_XI52/XI3/MM7_d N_XI52/XI3/NET35_XI52/XI3/MM7_g
+ N_VSS_XI52/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI3/MM8 N_XI52/XI3/NET35_XI52/XI3/MM8_d N_WL<101>_XI52/XI3/MM8_g
+ N_BLN<12>_XI52/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI3/MM5 N_XI52/XI3/NET34_XI52/XI3/MM5_d N_XI52/XI3/NET33_XI52/XI3/MM5_g
+ N_VDD_XI52/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI3/MM4 N_XI52/XI3/NET33_XI52/XI3/MM4_d N_XI52/XI3/NET34_XI52/XI3/MM4_g
+ N_VDD_XI52/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI3/MM10 N_XI52/XI3/NET35_XI52/XI3/MM10_d N_XI52/XI3/NET36_XI52/XI3/MM10_g
+ N_VDD_XI52/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI3/MM11 N_XI52/XI3/NET36_XI52/XI3/MM11_d N_XI52/XI3/NET35_XI52/XI3/MM11_g
+ N_VDD_XI52/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI4/MM2 N_XI52/XI4/NET34_XI52/XI4/MM2_d N_XI52/XI4/NET33_XI52/XI4/MM2_g
+ N_VSS_XI52/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI4/MM3 N_XI52/XI4/NET33_XI52/XI4/MM3_d N_WL<100>_XI52/XI4/MM3_g
+ N_BLN<11>_XI52/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI4/MM0 N_XI52/XI4/NET34_XI52/XI4/MM0_d N_WL<100>_XI52/XI4/MM0_g
+ N_BL<11>_XI52/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI4/MM1 N_XI52/XI4/NET33_XI52/XI4/MM1_d N_XI52/XI4/NET34_XI52/XI4/MM1_g
+ N_VSS_XI52/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI4/MM9 N_XI52/XI4/NET36_XI52/XI4/MM9_d N_WL<101>_XI52/XI4/MM9_g
+ N_BL<11>_XI52/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI4/MM6 N_XI52/XI4/NET35_XI52/XI4/MM6_d N_XI52/XI4/NET36_XI52/XI4/MM6_g
+ N_VSS_XI52/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI4/MM7 N_XI52/XI4/NET36_XI52/XI4/MM7_d N_XI52/XI4/NET35_XI52/XI4/MM7_g
+ N_VSS_XI52/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI4/MM8 N_XI52/XI4/NET35_XI52/XI4/MM8_d N_WL<101>_XI52/XI4/MM8_g
+ N_BLN<11>_XI52/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI4/MM5 N_XI52/XI4/NET34_XI52/XI4/MM5_d N_XI52/XI4/NET33_XI52/XI4/MM5_g
+ N_VDD_XI52/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI4/MM4 N_XI52/XI4/NET33_XI52/XI4/MM4_d N_XI52/XI4/NET34_XI52/XI4/MM4_g
+ N_VDD_XI52/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI4/MM10 N_XI52/XI4/NET35_XI52/XI4/MM10_d N_XI52/XI4/NET36_XI52/XI4/MM10_g
+ N_VDD_XI52/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI4/MM11 N_XI52/XI4/NET36_XI52/XI4/MM11_d N_XI52/XI4/NET35_XI52/XI4/MM11_g
+ N_VDD_XI52/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI5/MM2 N_XI52/XI5/NET34_XI52/XI5/MM2_d N_XI52/XI5/NET33_XI52/XI5/MM2_g
+ N_VSS_XI52/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI5/MM3 N_XI52/XI5/NET33_XI52/XI5/MM3_d N_WL<100>_XI52/XI5/MM3_g
+ N_BLN<10>_XI52/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI5/MM0 N_XI52/XI5/NET34_XI52/XI5/MM0_d N_WL<100>_XI52/XI5/MM0_g
+ N_BL<10>_XI52/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI5/MM1 N_XI52/XI5/NET33_XI52/XI5/MM1_d N_XI52/XI5/NET34_XI52/XI5/MM1_g
+ N_VSS_XI52/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI5/MM9 N_XI52/XI5/NET36_XI52/XI5/MM9_d N_WL<101>_XI52/XI5/MM9_g
+ N_BL<10>_XI52/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI5/MM6 N_XI52/XI5/NET35_XI52/XI5/MM6_d N_XI52/XI5/NET36_XI52/XI5/MM6_g
+ N_VSS_XI52/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI5/MM7 N_XI52/XI5/NET36_XI52/XI5/MM7_d N_XI52/XI5/NET35_XI52/XI5/MM7_g
+ N_VSS_XI52/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI5/MM8 N_XI52/XI5/NET35_XI52/XI5/MM8_d N_WL<101>_XI52/XI5/MM8_g
+ N_BLN<10>_XI52/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI5/MM5 N_XI52/XI5/NET34_XI52/XI5/MM5_d N_XI52/XI5/NET33_XI52/XI5/MM5_g
+ N_VDD_XI52/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI5/MM4 N_XI52/XI5/NET33_XI52/XI5/MM4_d N_XI52/XI5/NET34_XI52/XI5/MM4_g
+ N_VDD_XI52/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI5/MM10 N_XI52/XI5/NET35_XI52/XI5/MM10_d N_XI52/XI5/NET36_XI52/XI5/MM10_g
+ N_VDD_XI52/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI5/MM11 N_XI52/XI5/NET36_XI52/XI5/MM11_d N_XI52/XI5/NET35_XI52/XI5/MM11_g
+ N_VDD_XI52/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI6/MM2 N_XI52/XI6/NET34_XI52/XI6/MM2_d N_XI52/XI6/NET33_XI52/XI6/MM2_g
+ N_VSS_XI52/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM3 N_XI52/XI6/NET33_XI52/XI6/MM3_d N_WL<100>_XI52/XI6/MM3_g
+ N_BLN<9>_XI52/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM0 N_XI52/XI6/NET34_XI52/XI6/MM0_d N_WL<100>_XI52/XI6/MM0_g
+ N_BL<9>_XI52/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM1 N_XI52/XI6/NET33_XI52/XI6/MM1_d N_XI52/XI6/NET34_XI52/XI6/MM1_g
+ N_VSS_XI52/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM9 N_XI52/XI6/NET36_XI52/XI6/MM9_d N_WL<101>_XI52/XI6/MM9_g
+ N_BL<9>_XI52/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM6 N_XI52/XI6/NET35_XI52/XI6/MM6_d N_XI52/XI6/NET36_XI52/XI6/MM6_g
+ N_VSS_XI52/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM7 N_XI52/XI6/NET36_XI52/XI6/MM7_d N_XI52/XI6/NET35_XI52/XI6/MM7_g
+ N_VSS_XI52/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM8 N_XI52/XI6/NET35_XI52/XI6/MM8_d N_WL<101>_XI52/XI6/MM8_g
+ N_BLN<9>_XI52/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI6/MM5 N_XI52/XI6/NET34_XI52/XI6/MM5_d N_XI52/XI6/NET33_XI52/XI6/MM5_g
+ N_VDD_XI52/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI6/MM4 N_XI52/XI6/NET33_XI52/XI6/MM4_d N_XI52/XI6/NET34_XI52/XI6/MM4_g
+ N_VDD_XI52/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI6/MM10 N_XI52/XI6/NET35_XI52/XI6/MM10_d N_XI52/XI6/NET36_XI52/XI6/MM10_g
+ N_VDD_XI52/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI6/MM11 N_XI52/XI6/NET36_XI52/XI6/MM11_d N_XI52/XI6/NET35_XI52/XI6/MM11_g
+ N_VDD_XI52/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI7/MM2 N_XI52/XI7/NET34_XI52/XI7/MM2_d N_XI52/XI7/NET33_XI52/XI7/MM2_g
+ N_VSS_XI52/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM3 N_XI52/XI7/NET33_XI52/XI7/MM3_d N_WL<100>_XI52/XI7/MM3_g
+ N_BLN<8>_XI52/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM0 N_XI52/XI7/NET34_XI52/XI7/MM0_d N_WL<100>_XI52/XI7/MM0_g
+ N_BL<8>_XI52/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM1 N_XI52/XI7/NET33_XI52/XI7/MM1_d N_XI52/XI7/NET34_XI52/XI7/MM1_g
+ N_VSS_XI52/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM9 N_XI52/XI7/NET36_XI52/XI7/MM9_d N_WL<101>_XI52/XI7/MM9_g
+ N_BL<8>_XI52/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM6 N_XI52/XI7/NET35_XI52/XI7/MM6_d N_XI52/XI7/NET36_XI52/XI7/MM6_g
+ N_VSS_XI52/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM7 N_XI52/XI7/NET36_XI52/XI7/MM7_d N_XI52/XI7/NET35_XI52/XI7/MM7_g
+ N_VSS_XI52/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM8 N_XI52/XI7/NET35_XI52/XI7/MM8_d N_WL<101>_XI52/XI7/MM8_g
+ N_BLN<8>_XI52/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI7/MM5 N_XI52/XI7/NET34_XI52/XI7/MM5_d N_XI52/XI7/NET33_XI52/XI7/MM5_g
+ N_VDD_XI52/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI7/MM4 N_XI52/XI7/NET33_XI52/XI7/MM4_d N_XI52/XI7/NET34_XI52/XI7/MM4_g
+ N_VDD_XI52/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI7/MM10 N_XI52/XI7/NET35_XI52/XI7/MM10_d N_XI52/XI7/NET36_XI52/XI7/MM10_g
+ N_VDD_XI52/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI7/MM11 N_XI52/XI7/NET36_XI52/XI7/MM11_d N_XI52/XI7/NET35_XI52/XI7/MM11_g
+ N_VDD_XI52/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI8/MM2 N_XI52/XI8/NET34_XI52/XI8/MM2_d N_XI52/XI8/NET33_XI52/XI8/MM2_g
+ N_VSS_XI52/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM3 N_XI52/XI8/NET33_XI52/XI8/MM3_d N_WL<100>_XI52/XI8/MM3_g
+ N_BLN<7>_XI52/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM0 N_XI52/XI8/NET34_XI52/XI8/MM0_d N_WL<100>_XI52/XI8/MM0_g
+ N_BL<7>_XI52/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM1 N_XI52/XI8/NET33_XI52/XI8/MM1_d N_XI52/XI8/NET34_XI52/XI8/MM1_g
+ N_VSS_XI52/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM9 N_XI52/XI8/NET36_XI52/XI8/MM9_d N_WL<101>_XI52/XI8/MM9_g
+ N_BL<7>_XI52/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM6 N_XI52/XI8/NET35_XI52/XI8/MM6_d N_XI52/XI8/NET36_XI52/XI8/MM6_g
+ N_VSS_XI52/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM7 N_XI52/XI8/NET36_XI52/XI8/MM7_d N_XI52/XI8/NET35_XI52/XI8/MM7_g
+ N_VSS_XI52/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM8 N_XI52/XI8/NET35_XI52/XI8/MM8_d N_WL<101>_XI52/XI8/MM8_g
+ N_BLN<7>_XI52/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI8/MM5 N_XI52/XI8/NET34_XI52/XI8/MM5_d N_XI52/XI8/NET33_XI52/XI8/MM5_g
+ N_VDD_XI52/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI8/MM4 N_XI52/XI8/NET33_XI52/XI8/MM4_d N_XI52/XI8/NET34_XI52/XI8/MM4_g
+ N_VDD_XI52/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI8/MM10 N_XI52/XI8/NET35_XI52/XI8/MM10_d N_XI52/XI8/NET36_XI52/XI8/MM10_g
+ N_VDD_XI52/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI8/MM11 N_XI52/XI8/NET36_XI52/XI8/MM11_d N_XI52/XI8/NET35_XI52/XI8/MM11_g
+ N_VDD_XI52/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI9/MM2 N_XI52/XI9/NET34_XI52/XI9/MM2_d N_XI52/XI9/NET33_XI52/XI9/MM2_g
+ N_VSS_XI52/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM3 N_XI52/XI9/NET33_XI52/XI9/MM3_d N_WL<100>_XI52/XI9/MM3_g
+ N_BLN<6>_XI52/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM0 N_XI52/XI9/NET34_XI52/XI9/MM0_d N_WL<100>_XI52/XI9/MM0_g
+ N_BL<6>_XI52/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM1 N_XI52/XI9/NET33_XI52/XI9/MM1_d N_XI52/XI9/NET34_XI52/XI9/MM1_g
+ N_VSS_XI52/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM9 N_XI52/XI9/NET36_XI52/XI9/MM9_d N_WL<101>_XI52/XI9/MM9_g
+ N_BL<6>_XI52/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM6 N_XI52/XI9/NET35_XI52/XI9/MM6_d N_XI52/XI9/NET36_XI52/XI9/MM6_g
+ N_VSS_XI52/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM7 N_XI52/XI9/NET36_XI52/XI9/MM7_d N_XI52/XI9/NET35_XI52/XI9/MM7_g
+ N_VSS_XI52/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM8 N_XI52/XI9/NET35_XI52/XI9/MM8_d N_WL<101>_XI52/XI9/MM8_g
+ N_BLN<6>_XI52/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI9/MM5 N_XI52/XI9/NET34_XI52/XI9/MM5_d N_XI52/XI9/NET33_XI52/XI9/MM5_g
+ N_VDD_XI52/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI9/MM4 N_XI52/XI9/NET33_XI52/XI9/MM4_d N_XI52/XI9/NET34_XI52/XI9/MM4_g
+ N_VDD_XI52/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI9/MM10 N_XI52/XI9/NET35_XI52/XI9/MM10_d N_XI52/XI9/NET36_XI52/XI9/MM10_g
+ N_VDD_XI52/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI9/MM11 N_XI52/XI9/NET36_XI52/XI9/MM11_d N_XI52/XI9/NET35_XI52/XI9/MM11_g
+ N_VDD_XI52/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI10/MM2 N_XI52/XI10/NET34_XI52/XI10/MM2_d
+ N_XI52/XI10/NET33_XI52/XI10/MM2_g N_VSS_XI52/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI10/MM3 N_XI52/XI10/NET33_XI52/XI10/MM3_d N_WL<100>_XI52/XI10/MM3_g
+ N_BLN<5>_XI52/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI10/MM0 N_XI52/XI10/NET34_XI52/XI10/MM0_d N_WL<100>_XI52/XI10/MM0_g
+ N_BL<5>_XI52/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI10/MM1 N_XI52/XI10/NET33_XI52/XI10/MM1_d
+ N_XI52/XI10/NET34_XI52/XI10/MM1_g N_VSS_XI52/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI10/MM9 N_XI52/XI10/NET36_XI52/XI10/MM9_d N_WL<101>_XI52/XI10/MM9_g
+ N_BL<5>_XI52/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI10/MM6 N_XI52/XI10/NET35_XI52/XI10/MM6_d
+ N_XI52/XI10/NET36_XI52/XI10/MM6_g N_VSS_XI52/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI10/MM7 N_XI52/XI10/NET36_XI52/XI10/MM7_d
+ N_XI52/XI10/NET35_XI52/XI10/MM7_g N_VSS_XI52/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI10/MM8 N_XI52/XI10/NET35_XI52/XI10/MM8_d N_WL<101>_XI52/XI10/MM8_g
+ N_BLN<5>_XI52/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI10/MM5 N_XI52/XI10/NET34_XI52/XI10/MM5_d
+ N_XI52/XI10/NET33_XI52/XI10/MM5_g N_VDD_XI52/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI10/MM4 N_XI52/XI10/NET33_XI52/XI10/MM4_d
+ N_XI52/XI10/NET34_XI52/XI10/MM4_g N_VDD_XI52/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI10/MM10 N_XI52/XI10/NET35_XI52/XI10/MM10_d
+ N_XI52/XI10/NET36_XI52/XI10/MM10_g N_VDD_XI52/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI10/MM11 N_XI52/XI10/NET36_XI52/XI10/MM11_d
+ N_XI52/XI10/NET35_XI52/XI10/MM11_g N_VDD_XI52/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI11/MM2 N_XI52/XI11/NET34_XI52/XI11/MM2_d
+ N_XI52/XI11/NET33_XI52/XI11/MM2_g N_VSS_XI52/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI11/MM3 N_XI52/XI11/NET33_XI52/XI11/MM3_d N_WL<100>_XI52/XI11/MM3_g
+ N_BLN<4>_XI52/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI11/MM0 N_XI52/XI11/NET34_XI52/XI11/MM0_d N_WL<100>_XI52/XI11/MM0_g
+ N_BL<4>_XI52/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI11/MM1 N_XI52/XI11/NET33_XI52/XI11/MM1_d
+ N_XI52/XI11/NET34_XI52/XI11/MM1_g N_VSS_XI52/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI11/MM9 N_XI52/XI11/NET36_XI52/XI11/MM9_d N_WL<101>_XI52/XI11/MM9_g
+ N_BL<4>_XI52/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI11/MM6 N_XI52/XI11/NET35_XI52/XI11/MM6_d
+ N_XI52/XI11/NET36_XI52/XI11/MM6_g N_VSS_XI52/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI11/MM7 N_XI52/XI11/NET36_XI52/XI11/MM7_d
+ N_XI52/XI11/NET35_XI52/XI11/MM7_g N_VSS_XI52/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI11/MM8 N_XI52/XI11/NET35_XI52/XI11/MM8_d N_WL<101>_XI52/XI11/MM8_g
+ N_BLN<4>_XI52/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI11/MM5 N_XI52/XI11/NET34_XI52/XI11/MM5_d
+ N_XI52/XI11/NET33_XI52/XI11/MM5_g N_VDD_XI52/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI11/MM4 N_XI52/XI11/NET33_XI52/XI11/MM4_d
+ N_XI52/XI11/NET34_XI52/XI11/MM4_g N_VDD_XI52/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI11/MM10 N_XI52/XI11/NET35_XI52/XI11/MM10_d
+ N_XI52/XI11/NET36_XI52/XI11/MM10_g N_VDD_XI52/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI11/MM11 N_XI52/XI11/NET36_XI52/XI11/MM11_d
+ N_XI52/XI11/NET35_XI52/XI11/MM11_g N_VDD_XI52/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI12/MM2 N_XI52/XI12/NET34_XI52/XI12/MM2_d
+ N_XI52/XI12/NET33_XI52/XI12/MM2_g N_VSS_XI52/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI12/MM3 N_XI52/XI12/NET33_XI52/XI12/MM3_d N_WL<100>_XI52/XI12/MM3_g
+ N_BLN<3>_XI52/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI12/MM0 N_XI52/XI12/NET34_XI52/XI12/MM0_d N_WL<100>_XI52/XI12/MM0_g
+ N_BL<3>_XI52/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI12/MM1 N_XI52/XI12/NET33_XI52/XI12/MM1_d
+ N_XI52/XI12/NET34_XI52/XI12/MM1_g N_VSS_XI52/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI12/MM9 N_XI52/XI12/NET36_XI52/XI12/MM9_d N_WL<101>_XI52/XI12/MM9_g
+ N_BL<3>_XI52/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI12/MM6 N_XI52/XI12/NET35_XI52/XI12/MM6_d
+ N_XI52/XI12/NET36_XI52/XI12/MM6_g N_VSS_XI52/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI12/MM7 N_XI52/XI12/NET36_XI52/XI12/MM7_d
+ N_XI52/XI12/NET35_XI52/XI12/MM7_g N_VSS_XI52/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI12/MM8 N_XI52/XI12/NET35_XI52/XI12/MM8_d N_WL<101>_XI52/XI12/MM8_g
+ N_BLN<3>_XI52/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI12/MM5 N_XI52/XI12/NET34_XI52/XI12/MM5_d
+ N_XI52/XI12/NET33_XI52/XI12/MM5_g N_VDD_XI52/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI12/MM4 N_XI52/XI12/NET33_XI52/XI12/MM4_d
+ N_XI52/XI12/NET34_XI52/XI12/MM4_g N_VDD_XI52/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI12/MM10 N_XI52/XI12/NET35_XI52/XI12/MM10_d
+ N_XI52/XI12/NET36_XI52/XI12/MM10_g N_VDD_XI52/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI12/MM11 N_XI52/XI12/NET36_XI52/XI12/MM11_d
+ N_XI52/XI12/NET35_XI52/XI12/MM11_g N_VDD_XI52/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI13/MM2 N_XI52/XI13/NET34_XI52/XI13/MM2_d
+ N_XI52/XI13/NET33_XI52/XI13/MM2_g N_VSS_XI52/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI13/MM3 N_XI52/XI13/NET33_XI52/XI13/MM3_d N_WL<100>_XI52/XI13/MM3_g
+ N_BLN<2>_XI52/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI13/MM0 N_XI52/XI13/NET34_XI52/XI13/MM0_d N_WL<100>_XI52/XI13/MM0_g
+ N_BL<2>_XI52/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI13/MM1 N_XI52/XI13/NET33_XI52/XI13/MM1_d
+ N_XI52/XI13/NET34_XI52/XI13/MM1_g N_VSS_XI52/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI13/MM9 N_XI52/XI13/NET36_XI52/XI13/MM9_d N_WL<101>_XI52/XI13/MM9_g
+ N_BL<2>_XI52/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI13/MM6 N_XI52/XI13/NET35_XI52/XI13/MM6_d
+ N_XI52/XI13/NET36_XI52/XI13/MM6_g N_VSS_XI52/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI13/MM7 N_XI52/XI13/NET36_XI52/XI13/MM7_d
+ N_XI52/XI13/NET35_XI52/XI13/MM7_g N_VSS_XI52/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI13/MM8 N_XI52/XI13/NET35_XI52/XI13/MM8_d N_WL<101>_XI52/XI13/MM8_g
+ N_BLN<2>_XI52/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI13/MM5 N_XI52/XI13/NET34_XI52/XI13/MM5_d
+ N_XI52/XI13/NET33_XI52/XI13/MM5_g N_VDD_XI52/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI13/MM4 N_XI52/XI13/NET33_XI52/XI13/MM4_d
+ N_XI52/XI13/NET34_XI52/XI13/MM4_g N_VDD_XI52/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI13/MM10 N_XI52/XI13/NET35_XI52/XI13/MM10_d
+ N_XI52/XI13/NET36_XI52/XI13/MM10_g N_VDD_XI52/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI13/MM11 N_XI52/XI13/NET36_XI52/XI13/MM11_d
+ N_XI52/XI13/NET35_XI52/XI13/MM11_g N_VDD_XI52/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI14/MM2 N_XI52/XI14/NET34_XI52/XI14/MM2_d
+ N_XI52/XI14/NET33_XI52/XI14/MM2_g N_VSS_XI52/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI14/MM3 N_XI52/XI14/NET33_XI52/XI14/MM3_d N_WL<100>_XI52/XI14/MM3_g
+ N_BLN<1>_XI52/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI14/MM0 N_XI52/XI14/NET34_XI52/XI14/MM0_d N_WL<100>_XI52/XI14/MM0_g
+ N_BL<1>_XI52/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI14/MM1 N_XI52/XI14/NET33_XI52/XI14/MM1_d
+ N_XI52/XI14/NET34_XI52/XI14/MM1_g N_VSS_XI52/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI14/MM9 N_XI52/XI14/NET36_XI52/XI14/MM9_d N_WL<101>_XI52/XI14/MM9_g
+ N_BL<1>_XI52/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI14/MM6 N_XI52/XI14/NET35_XI52/XI14/MM6_d
+ N_XI52/XI14/NET36_XI52/XI14/MM6_g N_VSS_XI52/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI14/MM7 N_XI52/XI14/NET36_XI52/XI14/MM7_d
+ N_XI52/XI14/NET35_XI52/XI14/MM7_g N_VSS_XI52/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI14/MM8 N_XI52/XI14/NET35_XI52/XI14/MM8_d N_WL<101>_XI52/XI14/MM8_g
+ N_BLN<1>_XI52/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI14/MM5 N_XI52/XI14/NET34_XI52/XI14/MM5_d
+ N_XI52/XI14/NET33_XI52/XI14/MM5_g N_VDD_XI52/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI14/MM4 N_XI52/XI14/NET33_XI52/XI14/MM4_d
+ N_XI52/XI14/NET34_XI52/XI14/MM4_g N_VDD_XI52/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI14/MM10 N_XI52/XI14/NET35_XI52/XI14/MM10_d
+ N_XI52/XI14/NET36_XI52/XI14/MM10_g N_VDD_XI52/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI14/MM11 N_XI52/XI14/NET36_XI52/XI14/MM11_d
+ N_XI52/XI14/NET35_XI52/XI14/MM11_g N_VDD_XI52/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI15/MM2 N_XI52/XI15/NET34_XI52/XI15/MM2_d
+ N_XI52/XI15/NET33_XI52/XI15/MM2_g N_VSS_XI52/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI15/MM3 N_XI52/XI15/NET33_XI52/XI15/MM3_d N_WL<100>_XI52/XI15/MM3_g
+ N_BLN<0>_XI52/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI15/MM0 N_XI52/XI15/NET34_XI52/XI15/MM0_d N_WL<100>_XI52/XI15/MM0_g
+ N_BL<0>_XI52/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI15/MM1 N_XI52/XI15/NET33_XI52/XI15/MM1_d
+ N_XI52/XI15/NET34_XI52/XI15/MM1_g N_VSS_XI52/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI15/MM9 N_XI52/XI15/NET36_XI52/XI15/MM9_d N_WL<101>_XI52/XI15/MM9_g
+ N_BL<0>_XI52/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI15/MM6 N_XI52/XI15/NET35_XI52/XI15/MM6_d
+ N_XI52/XI15/NET36_XI52/XI15/MM6_g N_VSS_XI52/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI15/MM7 N_XI52/XI15/NET36_XI52/XI15/MM7_d
+ N_XI52/XI15/NET35_XI52/XI15/MM7_g N_VSS_XI52/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI52/XI15/MM8 N_XI52/XI15/NET35_XI52/XI15/MM8_d N_WL<101>_XI52/XI15/MM8_g
+ N_BLN<0>_XI52/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI52/XI15/MM5 N_XI52/XI15/NET34_XI52/XI15/MM5_d
+ N_XI52/XI15/NET33_XI52/XI15/MM5_g N_VDD_XI52/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI15/MM4 N_XI52/XI15/NET33_XI52/XI15/MM4_d
+ N_XI52/XI15/NET34_XI52/XI15/MM4_g N_VDD_XI52/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI15/MM10 N_XI52/XI15/NET35_XI52/XI15/MM10_d
+ N_XI52/XI15/NET36_XI52/XI15/MM10_g N_VDD_XI52/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI52/XI15/MM11 N_XI52/XI15/NET36_XI52/XI15/MM11_d
+ N_XI52/XI15/NET35_XI52/XI15/MM11_g N_VDD_XI52/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI0/MM2 N_XI53/XI0/NET34_XI53/XI0/MM2_d N_XI53/XI0/NET33_XI53/XI0/MM2_g
+ N_VSS_XI53/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI0/MM3 N_XI53/XI0/NET33_XI53/XI0/MM3_d N_WL<102>_XI53/XI0/MM3_g
+ N_BLN<15>_XI53/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI0/MM0 N_XI53/XI0/NET34_XI53/XI0/MM0_d N_WL<102>_XI53/XI0/MM0_g
+ N_BL<15>_XI53/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI0/MM1 N_XI53/XI0/NET33_XI53/XI0/MM1_d N_XI53/XI0/NET34_XI53/XI0/MM1_g
+ N_VSS_XI53/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI0/MM9 N_XI53/XI0/NET36_XI53/XI0/MM9_d N_WL<103>_XI53/XI0/MM9_g
+ N_BL<15>_XI53/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI0/MM6 N_XI53/XI0/NET35_XI53/XI0/MM6_d N_XI53/XI0/NET36_XI53/XI0/MM6_g
+ N_VSS_XI53/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI0/MM7 N_XI53/XI0/NET36_XI53/XI0/MM7_d N_XI53/XI0/NET35_XI53/XI0/MM7_g
+ N_VSS_XI53/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI0/MM8 N_XI53/XI0/NET35_XI53/XI0/MM8_d N_WL<103>_XI53/XI0/MM8_g
+ N_BLN<15>_XI53/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI0/MM5 N_XI53/XI0/NET34_XI53/XI0/MM5_d N_XI53/XI0/NET33_XI53/XI0/MM5_g
+ N_VDD_XI53/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI0/MM4 N_XI53/XI0/NET33_XI53/XI0/MM4_d N_XI53/XI0/NET34_XI53/XI0/MM4_g
+ N_VDD_XI53/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI0/MM10 N_XI53/XI0/NET35_XI53/XI0/MM10_d N_XI53/XI0/NET36_XI53/XI0/MM10_g
+ N_VDD_XI53/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI0/MM11 N_XI53/XI0/NET36_XI53/XI0/MM11_d N_XI53/XI0/NET35_XI53/XI0/MM11_g
+ N_VDD_XI53/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI1/MM2 N_XI53/XI1/NET34_XI53/XI1/MM2_d N_XI53/XI1/NET33_XI53/XI1/MM2_g
+ N_VSS_XI53/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI1/MM3 N_XI53/XI1/NET33_XI53/XI1/MM3_d N_WL<102>_XI53/XI1/MM3_g
+ N_BLN<14>_XI53/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI1/MM0 N_XI53/XI1/NET34_XI53/XI1/MM0_d N_WL<102>_XI53/XI1/MM0_g
+ N_BL<14>_XI53/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI1/MM1 N_XI53/XI1/NET33_XI53/XI1/MM1_d N_XI53/XI1/NET34_XI53/XI1/MM1_g
+ N_VSS_XI53/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI1/MM9 N_XI53/XI1/NET36_XI53/XI1/MM9_d N_WL<103>_XI53/XI1/MM9_g
+ N_BL<14>_XI53/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI1/MM6 N_XI53/XI1/NET35_XI53/XI1/MM6_d N_XI53/XI1/NET36_XI53/XI1/MM6_g
+ N_VSS_XI53/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI1/MM7 N_XI53/XI1/NET36_XI53/XI1/MM7_d N_XI53/XI1/NET35_XI53/XI1/MM7_g
+ N_VSS_XI53/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI1/MM8 N_XI53/XI1/NET35_XI53/XI1/MM8_d N_WL<103>_XI53/XI1/MM8_g
+ N_BLN<14>_XI53/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI1/MM5 N_XI53/XI1/NET34_XI53/XI1/MM5_d N_XI53/XI1/NET33_XI53/XI1/MM5_g
+ N_VDD_XI53/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI1/MM4 N_XI53/XI1/NET33_XI53/XI1/MM4_d N_XI53/XI1/NET34_XI53/XI1/MM4_g
+ N_VDD_XI53/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI1/MM10 N_XI53/XI1/NET35_XI53/XI1/MM10_d N_XI53/XI1/NET36_XI53/XI1/MM10_g
+ N_VDD_XI53/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI1/MM11 N_XI53/XI1/NET36_XI53/XI1/MM11_d N_XI53/XI1/NET35_XI53/XI1/MM11_g
+ N_VDD_XI53/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI2/MM2 N_XI53/XI2/NET34_XI53/XI2/MM2_d N_XI53/XI2/NET33_XI53/XI2/MM2_g
+ N_VSS_XI53/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI2/MM3 N_XI53/XI2/NET33_XI53/XI2/MM3_d N_WL<102>_XI53/XI2/MM3_g
+ N_BLN<13>_XI53/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI2/MM0 N_XI53/XI2/NET34_XI53/XI2/MM0_d N_WL<102>_XI53/XI2/MM0_g
+ N_BL<13>_XI53/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI2/MM1 N_XI53/XI2/NET33_XI53/XI2/MM1_d N_XI53/XI2/NET34_XI53/XI2/MM1_g
+ N_VSS_XI53/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI2/MM9 N_XI53/XI2/NET36_XI53/XI2/MM9_d N_WL<103>_XI53/XI2/MM9_g
+ N_BL<13>_XI53/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI2/MM6 N_XI53/XI2/NET35_XI53/XI2/MM6_d N_XI53/XI2/NET36_XI53/XI2/MM6_g
+ N_VSS_XI53/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI2/MM7 N_XI53/XI2/NET36_XI53/XI2/MM7_d N_XI53/XI2/NET35_XI53/XI2/MM7_g
+ N_VSS_XI53/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI2/MM8 N_XI53/XI2/NET35_XI53/XI2/MM8_d N_WL<103>_XI53/XI2/MM8_g
+ N_BLN<13>_XI53/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI2/MM5 N_XI53/XI2/NET34_XI53/XI2/MM5_d N_XI53/XI2/NET33_XI53/XI2/MM5_g
+ N_VDD_XI53/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI2/MM4 N_XI53/XI2/NET33_XI53/XI2/MM4_d N_XI53/XI2/NET34_XI53/XI2/MM4_g
+ N_VDD_XI53/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI2/MM10 N_XI53/XI2/NET35_XI53/XI2/MM10_d N_XI53/XI2/NET36_XI53/XI2/MM10_g
+ N_VDD_XI53/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI2/MM11 N_XI53/XI2/NET36_XI53/XI2/MM11_d N_XI53/XI2/NET35_XI53/XI2/MM11_g
+ N_VDD_XI53/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI3/MM2 N_XI53/XI3/NET34_XI53/XI3/MM2_d N_XI53/XI3/NET33_XI53/XI3/MM2_g
+ N_VSS_XI53/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI3/MM3 N_XI53/XI3/NET33_XI53/XI3/MM3_d N_WL<102>_XI53/XI3/MM3_g
+ N_BLN<12>_XI53/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI3/MM0 N_XI53/XI3/NET34_XI53/XI3/MM0_d N_WL<102>_XI53/XI3/MM0_g
+ N_BL<12>_XI53/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI3/MM1 N_XI53/XI3/NET33_XI53/XI3/MM1_d N_XI53/XI3/NET34_XI53/XI3/MM1_g
+ N_VSS_XI53/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI3/MM9 N_XI53/XI3/NET36_XI53/XI3/MM9_d N_WL<103>_XI53/XI3/MM9_g
+ N_BL<12>_XI53/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI3/MM6 N_XI53/XI3/NET35_XI53/XI3/MM6_d N_XI53/XI3/NET36_XI53/XI3/MM6_g
+ N_VSS_XI53/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI3/MM7 N_XI53/XI3/NET36_XI53/XI3/MM7_d N_XI53/XI3/NET35_XI53/XI3/MM7_g
+ N_VSS_XI53/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI3/MM8 N_XI53/XI3/NET35_XI53/XI3/MM8_d N_WL<103>_XI53/XI3/MM8_g
+ N_BLN<12>_XI53/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI3/MM5 N_XI53/XI3/NET34_XI53/XI3/MM5_d N_XI53/XI3/NET33_XI53/XI3/MM5_g
+ N_VDD_XI53/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI3/MM4 N_XI53/XI3/NET33_XI53/XI3/MM4_d N_XI53/XI3/NET34_XI53/XI3/MM4_g
+ N_VDD_XI53/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI3/MM10 N_XI53/XI3/NET35_XI53/XI3/MM10_d N_XI53/XI3/NET36_XI53/XI3/MM10_g
+ N_VDD_XI53/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI3/MM11 N_XI53/XI3/NET36_XI53/XI3/MM11_d N_XI53/XI3/NET35_XI53/XI3/MM11_g
+ N_VDD_XI53/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI4/MM2 N_XI53/XI4/NET34_XI53/XI4/MM2_d N_XI53/XI4/NET33_XI53/XI4/MM2_g
+ N_VSS_XI53/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI4/MM3 N_XI53/XI4/NET33_XI53/XI4/MM3_d N_WL<102>_XI53/XI4/MM3_g
+ N_BLN<11>_XI53/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI4/MM0 N_XI53/XI4/NET34_XI53/XI4/MM0_d N_WL<102>_XI53/XI4/MM0_g
+ N_BL<11>_XI53/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI4/MM1 N_XI53/XI4/NET33_XI53/XI4/MM1_d N_XI53/XI4/NET34_XI53/XI4/MM1_g
+ N_VSS_XI53/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI4/MM9 N_XI53/XI4/NET36_XI53/XI4/MM9_d N_WL<103>_XI53/XI4/MM9_g
+ N_BL<11>_XI53/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI4/MM6 N_XI53/XI4/NET35_XI53/XI4/MM6_d N_XI53/XI4/NET36_XI53/XI4/MM6_g
+ N_VSS_XI53/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI4/MM7 N_XI53/XI4/NET36_XI53/XI4/MM7_d N_XI53/XI4/NET35_XI53/XI4/MM7_g
+ N_VSS_XI53/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI4/MM8 N_XI53/XI4/NET35_XI53/XI4/MM8_d N_WL<103>_XI53/XI4/MM8_g
+ N_BLN<11>_XI53/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI4/MM5 N_XI53/XI4/NET34_XI53/XI4/MM5_d N_XI53/XI4/NET33_XI53/XI4/MM5_g
+ N_VDD_XI53/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI4/MM4 N_XI53/XI4/NET33_XI53/XI4/MM4_d N_XI53/XI4/NET34_XI53/XI4/MM4_g
+ N_VDD_XI53/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI4/MM10 N_XI53/XI4/NET35_XI53/XI4/MM10_d N_XI53/XI4/NET36_XI53/XI4/MM10_g
+ N_VDD_XI53/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI4/MM11 N_XI53/XI4/NET36_XI53/XI4/MM11_d N_XI53/XI4/NET35_XI53/XI4/MM11_g
+ N_VDD_XI53/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI5/MM2 N_XI53/XI5/NET34_XI53/XI5/MM2_d N_XI53/XI5/NET33_XI53/XI5/MM2_g
+ N_VSS_XI53/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI5/MM3 N_XI53/XI5/NET33_XI53/XI5/MM3_d N_WL<102>_XI53/XI5/MM3_g
+ N_BLN<10>_XI53/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI5/MM0 N_XI53/XI5/NET34_XI53/XI5/MM0_d N_WL<102>_XI53/XI5/MM0_g
+ N_BL<10>_XI53/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI5/MM1 N_XI53/XI5/NET33_XI53/XI5/MM1_d N_XI53/XI5/NET34_XI53/XI5/MM1_g
+ N_VSS_XI53/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI5/MM9 N_XI53/XI5/NET36_XI53/XI5/MM9_d N_WL<103>_XI53/XI5/MM9_g
+ N_BL<10>_XI53/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI5/MM6 N_XI53/XI5/NET35_XI53/XI5/MM6_d N_XI53/XI5/NET36_XI53/XI5/MM6_g
+ N_VSS_XI53/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI5/MM7 N_XI53/XI5/NET36_XI53/XI5/MM7_d N_XI53/XI5/NET35_XI53/XI5/MM7_g
+ N_VSS_XI53/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI5/MM8 N_XI53/XI5/NET35_XI53/XI5/MM8_d N_WL<103>_XI53/XI5/MM8_g
+ N_BLN<10>_XI53/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI5/MM5 N_XI53/XI5/NET34_XI53/XI5/MM5_d N_XI53/XI5/NET33_XI53/XI5/MM5_g
+ N_VDD_XI53/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI5/MM4 N_XI53/XI5/NET33_XI53/XI5/MM4_d N_XI53/XI5/NET34_XI53/XI5/MM4_g
+ N_VDD_XI53/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI5/MM10 N_XI53/XI5/NET35_XI53/XI5/MM10_d N_XI53/XI5/NET36_XI53/XI5/MM10_g
+ N_VDD_XI53/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI5/MM11 N_XI53/XI5/NET36_XI53/XI5/MM11_d N_XI53/XI5/NET35_XI53/XI5/MM11_g
+ N_VDD_XI53/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI6/MM2 N_XI53/XI6/NET34_XI53/XI6/MM2_d N_XI53/XI6/NET33_XI53/XI6/MM2_g
+ N_VSS_XI53/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM3 N_XI53/XI6/NET33_XI53/XI6/MM3_d N_WL<102>_XI53/XI6/MM3_g
+ N_BLN<9>_XI53/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM0 N_XI53/XI6/NET34_XI53/XI6/MM0_d N_WL<102>_XI53/XI6/MM0_g
+ N_BL<9>_XI53/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM1 N_XI53/XI6/NET33_XI53/XI6/MM1_d N_XI53/XI6/NET34_XI53/XI6/MM1_g
+ N_VSS_XI53/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM9 N_XI53/XI6/NET36_XI53/XI6/MM9_d N_WL<103>_XI53/XI6/MM9_g
+ N_BL<9>_XI53/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM6 N_XI53/XI6/NET35_XI53/XI6/MM6_d N_XI53/XI6/NET36_XI53/XI6/MM6_g
+ N_VSS_XI53/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM7 N_XI53/XI6/NET36_XI53/XI6/MM7_d N_XI53/XI6/NET35_XI53/XI6/MM7_g
+ N_VSS_XI53/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM8 N_XI53/XI6/NET35_XI53/XI6/MM8_d N_WL<103>_XI53/XI6/MM8_g
+ N_BLN<9>_XI53/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI6/MM5 N_XI53/XI6/NET34_XI53/XI6/MM5_d N_XI53/XI6/NET33_XI53/XI6/MM5_g
+ N_VDD_XI53/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI6/MM4 N_XI53/XI6/NET33_XI53/XI6/MM4_d N_XI53/XI6/NET34_XI53/XI6/MM4_g
+ N_VDD_XI53/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI6/MM10 N_XI53/XI6/NET35_XI53/XI6/MM10_d N_XI53/XI6/NET36_XI53/XI6/MM10_g
+ N_VDD_XI53/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI6/MM11 N_XI53/XI6/NET36_XI53/XI6/MM11_d N_XI53/XI6/NET35_XI53/XI6/MM11_g
+ N_VDD_XI53/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI7/MM2 N_XI53/XI7/NET34_XI53/XI7/MM2_d N_XI53/XI7/NET33_XI53/XI7/MM2_g
+ N_VSS_XI53/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM3 N_XI53/XI7/NET33_XI53/XI7/MM3_d N_WL<102>_XI53/XI7/MM3_g
+ N_BLN<8>_XI53/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM0 N_XI53/XI7/NET34_XI53/XI7/MM0_d N_WL<102>_XI53/XI7/MM0_g
+ N_BL<8>_XI53/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM1 N_XI53/XI7/NET33_XI53/XI7/MM1_d N_XI53/XI7/NET34_XI53/XI7/MM1_g
+ N_VSS_XI53/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM9 N_XI53/XI7/NET36_XI53/XI7/MM9_d N_WL<103>_XI53/XI7/MM9_g
+ N_BL<8>_XI53/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM6 N_XI53/XI7/NET35_XI53/XI7/MM6_d N_XI53/XI7/NET36_XI53/XI7/MM6_g
+ N_VSS_XI53/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM7 N_XI53/XI7/NET36_XI53/XI7/MM7_d N_XI53/XI7/NET35_XI53/XI7/MM7_g
+ N_VSS_XI53/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM8 N_XI53/XI7/NET35_XI53/XI7/MM8_d N_WL<103>_XI53/XI7/MM8_g
+ N_BLN<8>_XI53/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI7/MM5 N_XI53/XI7/NET34_XI53/XI7/MM5_d N_XI53/XI7/NET33_XI53/XI7/MM5_g
+ N_VDD_XI53/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI7/MM4 N_XI53/XI7/NET33_XI53/XI7/MM4_d N_XI53/XI7/NET34_XI53/XI7/MM4_g
+ N_VDD_XI53/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI7/MM10 N_XI53/XI7/NET35_XI53/XI7/MM10_d N_XI53/XI7/NET36_XI53/XI7/MM10_g
+ N_VDD_XI53/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI7/MM11 N_XI53/XI7/NET36_XI53/XI7/MM11_d N_XI53/XI7/NET35_XI53/XI7/MM11_g
+ N_VDD_XI53/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI8/MM2 N_XI53/XI8/NET34_XI53/XI8/MM2_d N_XI53/XI8/NET33_XI53/XI8/MM2_g
+ N_VSS_XI53/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM3 N_XI53/XI8/NET33_XI53/XI8/MM3_d N_WL<102>_XI53/XI8/MM3_g
+ N_BLN<7>_XI53/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM0 N_XI53/XI8/NET34_XI53/XI8/MM0_d N_WL<102>_XI53/XI8/MM0_g
+ N_BL<7>_XI53/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM1 N_XI53/XI8/NET33_XI53/XI8/MM1_d N_XI53/XI8/NET34_XI53/XI8/MM1_g
+ N_VSS_XI53/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM9 N_XI53/XI8/NET36_XI53/XI8/MM9_d N_WL<103>_XI53/XI8/MM9_g
+ N_BL<7>_XI53/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM6 N_XI53/XI8/NET35_XI53/XI8/MM6_d N_XI53/XI8/NET36_XI53/XI8/MM6_g
+ N_VSS_XI53/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM7 N_XI53/XI8/NET36_XI53/XI8/MM7_d N_XI53/XI8/NET35_XI53/XI8/MM7_g
+ N_VSS_XI53/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM8 N_XI53/XI8/NET35_XI53/XI8/MM8_d N_WL<103>_XI53/XI8/MM8_g
+ N_BLN<7>_XI53/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI8/MM5 N_XI53/XI8/NET34_XI53/XI8/MM5_d N_XI53/XI8/NET33_XI53/XI8/MM5_g
+ N_VDD_XI53/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI8/MM4 N_XI53/XI8/NET33_XI53/XI8/MM4_d N_XI53/XI8/NET34_XI53/XI8/MM4_g
+ N_VDD_XI53/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI8/MM10 N_XI53/XI8/NET35_XI53/XI8/MM10_d N_XI53/XI8/NET36_XI53/XI8/MM10_g
+ N_VDD_XI53/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI8/MM11 N_XI53/XI8/NET36_XI53/XI8/MM11_d N_XI53/XI8/NET35_XI53/XI8/MM11_g
+ N_VDD_XI53/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI9/MM2 N_XI53/XI9/NET34_XI53/XI9/MM2_d N_XI53/XI9/NET33_XI53/XI9/MM2_g
+ N_VSS_XI53/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM3 N_XI53/XI9/NET33_XI53/XI9/MM3_d N_WL<102>_XI53/XI9/MM3_g
+ N_BLN<6>_XI53/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM0 N_XI53/XI9/NET34_XI53/XI9/MM0_d N_WL<102>_XI53/XI9/MM0_g
+ N_BL<6>_XI53/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM1 N_XI53/XI9/NET33_XI53/XI9/MM1_d N_XI53/XI9/NET34_XI53/XI9/MM1_g
+ N_VSS_XI53/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM9 N_XI53/XI9/NET36_XI53/XI9/MM9_d N_WL<103>_XI53/XI9/MM9_g
+ N_BL<6>_XI53/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM6 N_XI53/XI9/NET35_XI53/XI9/MM6_d N_XI53/XI9/NET36_XI53/XI9/MM6_g
+ N_VSS_XI53/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM7 N_XI53/XI9/NET36_XI53/XI9/MM7_d N_XI53/XI9/NET35_XI53/XI9/MM7_g
+ N_VSS_XI53/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM8 N_XI53/XI9/NET35_XI53/XI9/MM8_d N_WL<103>_XI53/XI9/MM8_g
+ N_BLN<6>_XI53/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI9/MM5 N_XI53/XI9/NET34_XI53/XI9/MM5_d N_XI53/XI9/NET33_XI53/XI9/MM5_g
+ N_VDD_XI53/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI9/MM4 N_XI53/XI9/NET33_XI53/XI9/MM4_d N_XI53/XI9/NET34_XI53/XI9/MM4_g
+ N_VDD_XI53/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI9/MM10 N_XI53/XI9/NET35_XI53/XI9/MM10_d N_XI53/XI9/NET36_XI53/XI9/MM10_g
+ N_VDD_XI53/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI9/MM11 N_XI53/XI9/NET36_XI53/XI9/MM11_d N_XI53/XI9/NET35_XI53/XI9/MM11_g
+ N_VDD_XI53/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI10/MM2 N_XI53/XI10/NET34_XI53/XI10/MM2_d
+ N_XI53/XI10/NET33_XI53/XI10/MM2_g N_VSS_XI53/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI10/MM3 N_XI53/XI10/NET33_XI53/XI10/MM3_d N_WL<102>_XI53/XI10/MM3_g
+ N_BLN<5>_XI53/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI10/MM0 N_XI53/XI10/NET34_XI53/XI10/MM0_d N_WL<102>_XI53/XI10/MM0_g
+ N_BL<5>_XI53/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI10/MM1 N_XI53/XI10/NET33_XI53/XI10/MM1_d
+ N_XI53/XI10/NET34_XI53/XI10/MM1_g N_VSS_XI53/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI10/MM9 N_XI53/XI10/NET36_XI53/XI10/MM9_d N_WL<103>_XI53/XI10/MM9_g
+ N_BL<5>_XI53/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI10/MM6 N_XI53/XI10/NET35_XI53/XI10/MM6_d
+ N_XI53/XI10/NET36_XI53/XI10/MM6_g N_VSS_XI53/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI10/MM7 N_XI53/XI10/NET36_XI53/XI10/MM7_d
+ N_XI53/XI10/NET35_XI53/XI10/MM7_g N_VSS_XI53/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI10/MM8 N_XI53/XI10/NET35_XI53/XI10/MM8_d N_WL<103>_XI53/XI10/MM8_g
+ N_BLN<5>_XI53/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI10/MM5 N_XI53/XI10/NET34_XI53/XI10/MM5_d
+ N_XI53/XI10/NET33_XI53/XI10/MM5_g N_VDD_XI53/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI10/MM4 N_XI53/XI10/NET33_XI53/XI10/MM4_d
+ N_XI53/XI10/NET34_XI53/XI10/MM4_g N_VDD_XI53/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI10/MM10 N_XI53/XI10/NET35_XI53/XI10/MM10_d
+ N_XI53/XI10/NET36_XI53/XI10/MM10_g N_VDD_XI53/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI10/MM11 N_XI53/XI10/NET36_XI53/XI10/MM11_d
+ N_XI53/XI10/NET35_XI53/XI10/MM11_g N_VDD_XI53/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI11/MM2 N_XI53/XI11/NET34_XI53/XI11/MM2_d
+ N_XI53/XI11/NET33_XI53/XI11/MM2_g N_VSS_XI53/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI11/MM3 N_XI53/XI11/NET33_XI53/XI11/MM3_d N_WL<102>_XI53/XI11/MM3_g
+ N_BLN<4>_XI53/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI11/MM0 N_XI53/XI11/NET34_XI53/XI11/MM0_d N_WL<102>_XI53/XI11/MM0_g
+ N_BL<4>_XI53/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI11/MM1 N_XI53/XI11/NET33_XI53/XI11/MM1_d
+ N_XI53/XI11/NET34_XI53/XI11/MM1_g N_VSS_XI53/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI11/MM9 N_XI53/XI11/NET36_XI53/XI11/MM9_d N_WL<103>_XI53/XI11/MM9_g
+ N_BL<4>_XI53/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI11/MM6 N_XI53/XI11/NET35_XI53/XI11/MM6_d
+ N_XI53/XI11/NET36_XI53/XI11/MM6_g N_VSS_XI53/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI11/MM7 N_XI53/XI11/NET36_XI53/XI11/MM7_d
+ N_XI53/XI11/NET35_XI53/XI11/MM7_g N_VSS_XI53/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI11/MM8 N_XI53/XI11/NET35_XI53/XI11/MM8_d N_WL<103>_XI53/XI11/MM8_g
+ N_BLN<4>_XI53/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI11/MM5 N_XI53/XI11/NET34_XI53/XI11/MM5_d
+ N_XI53/XI11/NET33_XI53/XI11/MM5_g N_VDD_XI53/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI11/MM4 N_XI53/XI11/NET33_XI53/XI11/MM4_d
+ N_XI53/XI11/NET34_XI53/XI11/MM4_g N_VDD_XI53/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI11/MM10 N_XI53/XI11/NET35_XI53/XI11/MM10_d
+ N_XI53/XI11/NET36_XI53/XI11/MM10_g N_VDD_XI53/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI11/MM11 N_XI53/XI11/NET36_XI53/XI11/MM11_d
+ N_XI53/XI11/NET35_XI53/XI11/MM11_g N_VDD_XI53/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI12/MM2 N_XI53/XI12/NET34_XI53/XI12/MM2_d
+ N_XI53/XI12/NET33_XI53/XI12/MM2_g N_VSS_XI53/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI12/MM3 N_XI53/XI12/NET33_XI53/XI12/MM3_d N_WL<102>_XI53/XI12/MM3_g
+ N_BLN<3>_XI53/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI12/MM0 N_XI53/XI12/NET34_XI53/XI12/MM0_d N_WL<102>_XI53/XI12/MM0_g
+ N_BL<3>_XI53/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI12/MM1 N_XI53/XI12/NET33_XI53/XI12/MM1_d
+ N_XI53/XI12/NET34_XI53/XI12/MM1_g N_VSS_XI53/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI12/MM9 N_XI53/XI12/NET36_XI53/XI12/MM9_d N_WL<103>_XI53/XI12/MM9_g
+ N_BL<3>_XI53/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI12/MM6 N_XI53/XI12/NET35_XI53/XI12/MM6_d
+ N_XI53/XI12/NET36_XI53/XI12/MM6_g N_VSS_XI53/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI12/MM7 N_XI53/XI12/NET36_XI53/XI12/MM7_d
+ N_XI53/XI12/NET35_XI53/XI12/MM7_g N_VSS_XI53/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI12/MM8 N_XI53/XI12/NET35_XI53/XI12/MM8_d N_WL<103>_XI53/XI12/MM8_g
+ N_BLN<3>_XI53/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI12/MM5 N_XI53/XI12/NET34_XI53/XI12/MM5_d
+ N_XI53/XI12/NET33_XI53/XI12/MM5_g N_VDD_XI53/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI12/MM4 N_XI53/XI12/NET33_XI53/XI12/MM4_d
+ N_XI53/XI12/NET34_XI53/XI12/MM4_g N_VDD_XI53/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI12/MM10 N_XI53/XI12/NET35_XI53/XI12/MM10_d
+ N_XI53/XI12/NET36_XI53/XI12/MM10_g N_VDD_XI53/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI12/MM11 N_XI53/XI12/NET36_XI53/XI12/MM11_d
+ N_XI53/XI12/NET35_XI53/XI12/MM11_g N_VDD_XI53/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI13/MM2 N_XI53/XI13/NET34_XI53/XI13/MM2_d
+ N_XI53/XI13/NET33_XI53/XI13/MM2_g N_VSS_XI53/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI13/MM3 N_XI53/XI13/NET33_XI53/XI13/MM3_d N_WL<102>_XI53/XI13/MM3_g
+ N_BLN<2>_XI53/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI13/MM0 N_XI53/XI13/NET34_XI53/XI13/MM0_d N_WL<102>_XI53/XI13/MM0_g
+ N_BL<2>_XI53/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI13/MM1 N_XI53/XI13/NET33_XI53/XI13/MM1_d
+ N_XI53/XI13/NET34_XI53/XI13/MM1_g N_VSS_XI53/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI13/MM9 N_XI53/XI13/NET36_XI53/XI13/MM9_d N_WL<103>_XI53/XI13/MM9_g
+ N_BL<2>_XI53/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI13/MM6 N_XI53/XI13/NET35_XI53/XI13/MM6_d
+ N_XI53/XI13/NET36_XI53/XI13/MM6_g N_VSS_XI53/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI13/MM7 N_XI53/XI13/NET36_XI53/XI13/MM7_d
+ N_XI53/XI13/NET35_XI53/XI13/MM7_g N_VSS_XI53/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI13/MM8 N_XI53/XI13/NET35_XI53/XI13/MM8_d N_WL<103>_XI53/XI13/MM8_g
+ N_BLN<2>_XI53/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI13/MM5 N_XI53/XI13/NET34_XI53/XI13/MM5_d
+ N_XI53/XI13/NET33_XI53/XI13/MM5_g N_VDD_XI53/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI13/MM4 N_XI53/XI13/NET33_XI53/XI13/MM4_d
+ N_XI53/XI13/NET34_XI53/XI13/MM4_g N_VDD_XI53/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI13/MM10 N_XI53/XI13/NET35_XI53/XI13/MM10_d
+ N_XI53/XI13/NET36_XI53/XI13/MM10_g N_VDD_XI53/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI13/MM11 N_XI53/XI13/NET36_XI53/XI13/MM11_d
+ N_XI53/XI13/NET35_XI53/XI13/MM11_g N_VDD_XI53/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI14/MM2 N_XI53/XI14/NET34_XI53/XI14/MM2_d
+ N_XI53/XI14/NET33_XI53/XI14/MM2_g N_VSS_XI53/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI14/MM3 N_XI53/XI14/NET33_XI53/XI14/MM3_d N_WL<102>_XI53/XI14/MM3_g
+ N_BLN<1>_XI53/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI14/MM0 N_XI53/XI14/NET34_XI53/XI14/MM0_d N_WL<102>_XI53/XI14/MM0_g
+ N_BL<1>_XI53/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI14/MM1 N_XI53/XI14/NET33_XI53/XI14/MM1_d
+ N_XI53/XI14/NET34_XI53/XI14/MM1_g N_VSS_XI53/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI14/MM9 N_XI53/XI14/NET36_XI53/XI14/MM9_d N_WL<103>_XI53/XI14/MM9_g
+ N_BL<1>_XI53/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI14/MM6 N_XI53/XI14/NET35_XI53/XI14/MM6_d
+ N_XI53/XI14/NET36_XI53/XI14/MM6_g N_VSS_XI53/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI14/MM7 N_XI53/XI14/NET36_XI53/XI14/MM7_d
+ N_XI53/XI14/NET35_XI53/XI14/MM7_g N_VSS_XI53/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI14/MM8 N_XI53/XI14/NET35_XI53/XI14/MM8_d N_WL<103>_XI53/XI14/MM8_g
+ N_BLN<1>_XI53/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI14/MM5 N_XI53/XI14/NET34_XI53/XI14/MM5_d
+ N_XI53/XI14/NET33_XI53/XI14/MM5_g N_VDD_XI53/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI14/MM4 N_XI53/XI14/NET33_XI53/XI14/MM4_d
+ N_XI53/XI14/NET34_XI53/XI14/MM4_g N_VDD_XI53/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI14/MM10 N_XI53/XI14/NET35_XI53/XI14/MM10_d
+ N_XI53/XI14/NET36_XI53/XI14/MM10_g N_VDD_XI53/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI14/MM11 N_XI53/XI14/NET36_XI53/XI14/MM11_d
+ N_XI53/XI14/NET35_XI53/XI14/MM11_g N_VDD_XI53/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI15/MM2 N_XI53/XI15/NET34_XI53/XI15/MM2_d
+ N_XI53/XI15/NET33_XI53/XI15/MM2_g N_VSS_XI53/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI15/MM3 N_XI53/XI15/NET33_XI53/XI15/MM3_d N_WL<102>_XI53/XI15/MM3_g
+ N_BLN<0>_XI53/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI15/MM0 N_XI53/XI15/NET34_XI53/XI15/MM0_d N_WL<102>_XI53/XI15/MM0_g
+ N_BL<0>_XI53/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI15/MM1 N_XI53/XI15/NET33_XI53/XI15/MM1_d
+ N_XI53/XI15/NET34_XI53/XI15/MM1_g N_VSS_XI53/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI15/MM9 N_XI53/XI15/NET36_XI53/XI15/MM9_d N_WL<103>_XI53/XI15/MM9_g
+ N_BL<0>_XI53/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI15/MM6 N_XI53/XI15/NET35_XI53/XI15/MM6_d
+ N_XI53/XI15/NET36_XI53/XI15/MM6_g N_VSS_XI53/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI15/MM7 N_XI53/XI15/NET36_XI53/XI15/MM7_d
+ N_XI53/XI15/NET35_XI53/XI15/MM7_g N_VSS_XI53/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI53/XI15/MM8 N_XI53/XI15/NET35_XI53/XI15/MM8_d N_WL<103>_XI53/XI15/MM8_g
+ N_BLN<0>_XI53/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI53/XI15/MM5 N_XI53/XI15/NET34_XI53/XI15/MM5_d
+ N_XI53/XI15/NET33_XI53/XI15/MM5_g N_VDD_XI53/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI15/MM4 N_XI53/XI15/NET33_XI53/XI15/MM4_d
+ N_XI53/XI15/NET34_XI53/XI15/MM4_g N_VDD_XI53/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI15/MM10 N_XI53/XI15/NET35_XI53/XI15/MM10_d
+ N_XI53/XI15/NET36_XI53/XI15/MM10_g N_VDD_XI53/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI53/XI15/MM11 N_XI53/XI15/NET36_XI53/XI15/MM11_d
+ N_XI53/XI15/NET35_XI53/XI15/MM11_g N_VDD_XI53/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI0/MM2 N_XI54/XI0/NET34_XI54/XI0/MM2_d N_XI54/XI0/NET33_XI54/XI0/MM2_g
+ N_VSS_XI54/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI0/MM3 N_XI54/XI0/NET33_XI54/XI0/MM3_d N_WL<104>_XI54/XI0/MM3_g
+ N_BLN<15>_XI54/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI0/MM0 N_XI54/XI0/NET34_XI54/XI0/MM0_d N_WL<104>_XI54/XI0/MM0_g
+ N_BL<15>_XI54/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI0/MM1 N_XI54/XI0/NET33_XI54/XI0/MM1_d N_XI54/XI0/NET34_XI54/XI0/MM1_g
+ N_VSS_XI54/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI0/MM9 N_XI54/XI0/NET36_XI54/XI0/MM9_d N_WL<105>_XI54/XI0/MM9_g
+ N_BL<15>_XI54/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI0/MM6 N_XI54/XI0/NET35_XI54/XI0/MM6_d N_XI54/XI0/NET36_XI54/XI0/MM6_g
+ N_VSS_XI54/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI0/MM7 N_XI54/XI0/NET36_XI54/XI0/MM7_d N_XI54/XI0/NET35_XI54/XI0/MM7_g
+ N_VSS_XI54/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI0/MM8 N_XI54/XI0/NET35_XI54/XI0/MM8_d N_WL<105>_XI54/XI0/MM8_g
+ N_BLN<15>_XI54/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI0/MM5 N_XI54/XI0/NET34_XI54/XI0/MM5_d N_XI54/XI0/NET33_XI54/XI0/MM5_g
+ N_VDD_XI54/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI0/MM4 N_XI54/XI0/NET33_XI54/XI0/MM4_d N_XI54/XI0/NET34_XI54/XI0/MM4_g
+ N_VDD_XI54/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI0/MM10 N_XI54/XI0/NET35_XI54/XI0/MM10_d N_XI54/XI0/NET36_XI54/XI0/MM10_g
+ N_VDD_XI54/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI0/MM11 N_XI54/XI0/NET36_XI54/XI0/MM11_d N_XI54/XI0/NET35_XI54/XI0/MM11_g
+ N_VDD_XI54/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI1/MM2 N_XI54/XI1/NET34_XI54/XI1/MM2_d N_XI54/XI1/NET33_XI54/XI1/MM2_g
+ N_VSS_XI54/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI1/MM3 N_XI54/XI1/NET33_XI54/XI1/MM3_d N_WL<104>_XI54/XI1/MM3_g
+ N_BLN<14>_XI54/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI1/MM0 N_XI54/XI1/NET34_XI54/XI1/MM0_d N_WL<104>_XI54/XI1/MM0_g
+ N_BL<14>_XI54/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI1/MM1 N_XI54/XI1/NET33_XI54/XI1/MM1_d N_XI54/XI1/NET34_XI54/XI1/MM1_g
+ N_VSS_XI54/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI1/MM9 N_XI54/XI1/NET36_XI54/XI1/MM9_d N_WL<105>_XI54/XI1/MM9_g
+ N_BL<14>_XI54/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI1/MM6 N_XI54/XI1/NET35_XI54/XI1/MM6_d N_XI54/XI1/NET36_XI54/XI1/MM6_g
+ N_VSS_XI54/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI1/MM7 N_XI54/XI1/NET36_XI54/XI1/MM7_d N_XI54/XI1/NET35_XI54/XI1/MM7_g
+ N_VSS_XI54/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI1/MM8 N_XI54/XI1/NET35_XI54/XI1/MM8_d N_WL<105>_XI54/XI1/MM8_g
+ N_BLN<14>_XI54/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI1/MM5 N_XI54/XI1/NET34_XI54/XI1/MM5_d N_XI54/XI1/NET33_XI54/XI1/MM5_g
+ N_VDD_XI54/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI1/MM4 N_XI54/XI1/NET33_XI54/XI1/MM4_d N_XI54/XI1/NET34_XI54/XI1/MM4_g
+ N_VDD_XI54/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI1/MM10 N_XI54/XI1/NET35_XI54/XI1/MM10_d N_XI54/XI1/NET36_XI54/XI1/MM10_g
+ N_VDD_XI54/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI1/MM11 N_XI54/XI1/NET36_XI54/XI1/MM11_d N_XI54/XI1/NET35_XI54/XI1/MM11_g
+ N_VDD_XI54/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI2/MM2 N_XI54/XI2/NET34_XI54/XI2/MM2_d N_XI54/XI2/NET33_XI54/XI2/MM2_g
+ N_VSS_XI54/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI2/MM3 N_XI54/XI2/NET33_XI54/XI2/MM3_d N_WL<104>_XI54/XI2/MM3_g
+ N_BLN<13>_XI54/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI2/MM0 N_XI54/XI2/NET34_XI54/XI2/MM0_d N_WL<104>_XI54/XI2/MM0_g
+ N_BL<13>_XI54/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI2/MM1 N_XI54/XI2/NET33_XI54/XI2/MM1_d N_XI54/XI2/NET34_XI54/XI2/MM1_g
+ N_VSS_XI54/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI2/MM9 N_XI54/XI2/NET36_XI54/XI2/MM9_d N_WL<105>_XI54/XI2/MM9_g
+ N_BL<13>_XI54/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI2/MM6 N_XI54/XI2/NET35_XI54/XI2/MM6_d N_XI54/XI2/NET36_XI54/XI2/MM6_g
+ N_VSS_XI54/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI2/MM7 N_XI54/XI2/NET36_XI54/XI2/MM7_d N_XI54/XI2/NET35_XI54/XI2/MM7_g
+ N_VSS_XI54/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI2/MM8 N_XI54/XI2/NET35_XI54/XI2/MM8_d N_WL<105>_XI54/XI2/MM8_g
+ N_BLN<13>_XI54/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI2/MM5 N_XI54/XI2/NET34_XI54/XI2/MM5_d N_XI54/XI2/NET33_XI54/XI2/MM5_g
+ N_VDD_XI54/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI2/MM4 N_XI54/XI2/NET33_XI54/XI2/MM4_d N_XI54/XI2/NET34_XI54/XI2/MM4_g
+ N_VDD_XI54/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI2/MM10 N_XI54/XI2/NET35_XI54/XI2/MM10_d N_XI54/XI2/NET36_XI54/XI2/MM10_g
+ N_VDD_XI54/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI2/MM11 N_XI54/XI2/NET36_XI54/XI2/MM11_d N_XI54/XI2/NET35_XI54/XI2/MM11_g
+ N_VDD_XI54/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI3/MM2 N_XI54/XI3/NET34_XI54/XI3/MM2_d N_XI54/XI3/NET33_XI54/XI3/MM2_g
+ N_VSS_XI54/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI3/MM3 N_XI54/XI3/NET33_XI54/XI3/MM3_d N_WL<104>_XI54/XI3/MM3_g
+ N_BLN<12>_XI54/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI3/MM0 N_XI54/XI3/NET34_XI54/XI3/MM0_d N_WL<104>_XI54/XI3/MM0_g
+ N_BL<12>_XI54/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI3/MM1 N_XI54/XI3/NET33_XI54/XI3/MM1_d N_XI54/XI3/NET34_XI54/XI3/MM1_g
+ N_VSS_XI54/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI3/MM9 N_XI54/XI3/NET36_XI54/XI3/MM9_d N_WL<105>_XI54/XI3/MM9_g
+ N_BL<12>_XI54/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI3/MM6 N_XI54/XI3/NET35_XI54/XI3/MM6_d N_XI54/XI3/NET36_XI54/XI3/MM6_g
+ N_VSS_XI54/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI3/MM7 N_XI54/XI3/NET36_XI54/XI3/MM7_d N_XI54/XI3/NET35_XI54/XI3/MM7_g
+ N_VSS_XI54/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI3/MM8 N_XI54/XI3/NET35_XI54/XI3/MM8_d N_WL<105>_XI54/XI3/MM8_g
+ N_BLN<12>_XI54/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI3/MM5 N_XI54/XI3/NET34_XI54/XI3/MM5_d N_XI54/XI3/NET33_XI54/XI3/MM5_g
+ N_VDD_XI54/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI3/MM4 N_XI54/XI3/NET33_XI54/XI3/MM4_d N_XI54/XI3/NET34_XI54/XI3/MM4_g
+ N_VDD_XI54/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI3/MM10 N_XI54/XI3/NET35_XI54/XI3/MM10_d N_XI54/XI3/NET36_XI54/XI3/MM10_g
+ N_VDD_XI54/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI3/MM11 N_XI54/XI3/NET36_XI54/XI3/MM11_d N_XI54/XI3/NET35_XI54/XI3/MM11_g
+ N_VDD_XI54/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI4/MM2 N_XI54/XI4/NET34_XI54/XI4/MM2_d N_XI54/XI4/NET33_XI54/XI4/MM2_g
+ N_VSS_XI54/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI4/MM3 N_XI54/XI4/NET33_XI54/XI4/MM3_d N_WL<104>_XI54/XI4/MM3_g
+ N_BLN<11>_XI54/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI4/MM0 N_XI54/XI4/NET34_XI54/XI4/MM0_d N_WL<104>_XI54/XI4/MM0_g
+ N_BL<11>_XI54/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI4/MM1 N_XI54/XI4/NET33_XI54/XI4/MM1_d N_XI54/XI4/NET34_XI54/XI4/MM1_g
+ N_VSS_XI54/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI4/MM9 N_XI54/XI4/NET36_XI54/XI4/MM9_d N_WL<105>_XI54/XI4/MM9_g
+ N_BL<11>_XI54/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI4/MM6 N_XI54/XI4/NET35_XI54/XI4/MM6_d N_XI54/XI4/NET36_XI54/XI4/MM6_g
+ N_VSS_XI54/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI4/MM7 N_XI54/XI4/NET36_XI54/XI4/MM7_d N_XI54/XI4/NET35_XI54/XI4/MM7_g
+ N_VSS_XI54/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI4/MM8 N_XI54/XI4/NET35_XI54/XI4/MM8_d N_WL<105>_XI54/XI4/MM8_g
+ N_BLN<11>_XI54/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI4/MM5 N_XI54/XI4/NET34_XI54/XI4/MM5_d N_XI54/XI4/NET33_XI54/XI4/MM5_g
+ N_VDD_XI54/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI4/MM4 N_XI54/XI4/NET33_XI54/XI4/MM4_d N_XI54/XI4/NET34_XI54/XI4/MM4_g
+ N_VDD_XI54/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI4/MM10 N_XI54/XI4/NET35_XI54/XI4/MM10_d N_XI54/XI4/NET36_XI54/XI4/MM10_g
+ N_VDD_XI54/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI4/MM11 N_XI54/XI4/NET36_XI54/XI4/MM11_d N_XI54/XI4/NET35_XI54/XI4/MM11_g
+ N_VDD_XI54/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI5/MM2 N_XI54/XI5/NET34_XI54/XI5/MM2_d N_XI54/XI5/NET33_XI54/XI5/MM2_g
+ N_VSS_XI54/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI5/MM3 N_XI54/XI5/NET33_XI54/XI5/MM3_d N_WL<104>_XI54/XI5/MM3_g
+ N_BLN<10>_XI54/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI5/MM0 N_XI54/XI5/NET34_XI54/XI5/MM0_d N_WL<104>_XI54/XI5/MM0_g
+ N_BL<10>_XI54/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI5/MM1 N_XI54/XI5/NET33_XI54/XI5/MM1_d N_XI54/XI5/NET34_XI54/XI5/MM1_g
+ N_VSS_XI54/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI5/MM9 N_XI54/XI5/NET36_XI54/XI5/MM9_d N_WL<105>_XI54/XI5/MM9_g
+ N_BL<10>_XI54/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI5/MM6 N_XI54/XI5/NET35_XI54/XI5/MM6_d N_XI54/XI5/NET36_XI54/XI5/MM6_g
+ N_VSS_XI54/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI5/MM7 N_XI54/XI5/NET36_XI54/XI5/MM7_d N_XI54/XI5/NET35_XI54/XI5/MM7_g
+ N_VSS_XI54/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI5/MM8 N_XI54/XI5/NET35_XI54/XI5/MM8_d N_WL<105>_XI54/XI5/MM8_g
+ N_BLN<10>_XI54/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI5/MM5 N_XI54/XI5/NET34_XI54/XI5/MM5_d N_XI54/XI5/NET33_XI54/XI5/MM5_g
+ N_VDD_XI54/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI5/MM4 N_XI54/XI5/NET33_XI54/XI5/MM4_d N_XI54/XI5/NET34_XI54/XI5/MM4_g
+ N_VDD_XI54/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI5/MM10 N_XI54/XI5/NET35_XI54/XI5/MM10_d N_XI54/XI5/NET36_XI54/XI5/MM10_g
+ N_VDD_XI54/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI5/MM11 N_XI54/XI5/NET36_XI54/XI5/MM11_d N_XI54/XI5/NET35_XI54/XI5/MM11_g
+ N_VDD_XI54/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI6/MM2 N_XI54/XI6/NET34_XI54/XI6/MM2_d N_XI54/XI6/NET33_XI54/XI6/MM2_g
+ N_VSS_XI54/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM3 N_XI54/XI6/NET33_XI54/XI6/MM3_d N_WL<104>_XI54/XI6/MM3_g
+ N_BLN<9>_XI54/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM0 N_XI54/XI6/NET34_XI54/XI6/MM0_d N_WL<104>_XI54/XI6/MM0_g
+ N_BL<9>_XI54/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM1 N_XI54/XI6/NET33_XI54/XI6/MM1_d N_XI54/XI6/NET34_XI54/XI6/MM1_g
+ N_VSS_XI54/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM9 N_XI54/XI6/NET36_XI54/XI6/MM9_d N_WL<105>_XI54/XI6/MM9_g
+ N_BL<9>_XI54/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM6 N_XI54/XI6/NET35_XI54/XI6/MM6_d N_XI54/XI6/NET36_XI54/XI6/MM6_g
+ N_VSS_XI54/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM7 N_XI54/XI6/NET36_XI54/XI6/MM7_d N_XI54/XI6/NET35_XI54/XI6/MM7_g
+ N_VSS_XI54/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM8 N_XI54/XI6/NET35_XI54/XI6/MM8_d N_WL<105>_XI54/XI6/MM8_g
+ N_BLN<9>_XI54/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI6/MM5 N_XI54/XI6/NET34_XI54/XI6/MM5_d N_XI54/XI6/NET33_XI54/XI6/MM5_g
+ N_VDD_XI54/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI6/MM4 N_XI54/XI6/NET33_XI54/XI6/MM4_d N_XI54/XI6/NET34_XI54/XI6/MM4_g
+ N_VDD_XI54/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI6/MM10 N_XI54/XI6/NET35_XI54/XI6/MM10_d N_XI54/XI6/NET36_XI54/XI6/MM10_g
+ N_VDD_XI54/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI6/MM11 N_XI54/XI6/NET36_XI54/XI6/MM11_d N_XI54/XI6/NET35_XI54/XI6/MM11_g
+ N_VDD_XI54/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI7/MM2 N_XI54/XI7/NET34_XI54/XI7/MM2_d N_XI54/XI7/NET33_XI54/XI7/MM2_g
+ N_VSS_XI54/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM3 N_XI54/XI7/NET33_XI54/XI7/MM3_d N_WL<104>_XI54/XI7/MM3_g
+ N_BLN<8>_XI54/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM0 N_XI54/XI7/NET34_XI54/XI7/MM0_d N_WL<104>_XI54/XI7/MM0_g
+ N_BL<8>_XI54/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM1 N_XI54/XI7/NET33_XI54/XI7/MM1_d N_XI54/XI7/NET34_XI54/XI7/MM1_g
+ N_VSS_XI54/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM9 N_XI54/XI7/NET36_XI54/XI7/MM9_d N_WL<105>_XI54/XI7/MM9_g
+ N_BL<8>_XI54/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM6 N_XI54/XI7/NET35_XI54/XI7/MM6_d N_XI54/XI7/NET36_XI54/XI7/MM6_g
+ N_VSS_XI54/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM7 N_XI54/XI7/NET36_XI54/XI7/MM7_d N_XI54/XI7/NET35_XI54/XI7/MM7_g
+ N_VSS_XI54/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM8 N_XI54/XI7/NET35_XI54/XI7/MM8_d N_WL<105>_XI54/XI7/MM8_g
+ N_BLN<8>_XI54/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI7/MM5 N_XI54/XI7/NET34_XI54/XI7/MM5_d N_XI54/XI7/NET33_XI54/XI7/MM5_g
+ N_VDD_XI54/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI7/MM4 N_XI54/XI7/NET33_XI54/XI7/MM4_d N_XI54/XI7/NET34_XI54/XI7/MM4_g
+ N_VDD_XI54/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI7/MM10 N_XI54/XI7/NET35_XI54/XI7/MM10_d N_XI54/XI7/NET36_XI54/XI7/MM10_g
+ N_VDD_XI54/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI7/MM11 N_XI54/XI7/NET36_XI54/XI7/MM11_d N_XI54/XI7/NET35_XI54/XI7/MM11_g
+ N_VDD_XI54/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI8/MM2 N_XI54/XI8/NET34_XI54/XI8/MM2_d N_XI54/XI8/NET33_XI54/XI8/MM2_g
+ N_VSS_XI54/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM3 N_XI54/XI8/NET33_XI54/XI8/MM3_d N_WL<104>_XI54/XI8/MM3_g
+ N_BLN<7>_XI54/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM0 N_XI54/XI8/NET34_XI54/XI8/MM0_d N_WL<104>_XI54/XI8/MM0_g
+ N_BL<7>_XI54/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM1 N_XI54/XI8/NET33_XI54/XI8/MM1_d N_XI54/XI8/NET34_XI54/XI8/MM1_g
+ N_VSS_XI54/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM9 N_XI54/XI8/NET36_XI54/XI8/MM9_d N_WL<105>_XI54/XI8/MM9_g
+ N_BL<7>_XI54/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM6 N_XI54/XI8/NET35_XI54/XI8/MM6_d N_XI54/XI8/NET36_XI54/XI8/MM6_g
+ N_VSS_XI54/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM7 N_XI54/XI8/NET36_XI54/XI8/MM7_d N_XI54/XI8/NET35_XI54/XI8/MM7_g
+ N_VSS_XI54/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM8 N_XI54/XI8/NET35_XI54/XI8/MM8_d N_WL<105>_XI54/XI8/MM8_g
+ N_BLN<7>_XI54/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI8/MM5 N_XI54/XI8/NET34_XI54/XI8/MM5_d N_XI54/XI8/NET33_XI54/XI8/MM5_g
+ N_VDD_XI54/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI8/MM4 N_XI54/XI8/NET33_XI54/XI8/MM4_d N_XI54/XI8/NET34_XI54/XI8/MM4_g
+ N_VDD_XI54/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI8/MM10 N_XI54/XI8/NET35_XI54/XI8/MM10_d N_XI54/XI8/NET36_XI54/XI8/MM10_g
+ N_VDD_XI54/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI8/MM11 N_XI54/XI8/NET36_XI54/XI8/MM11_d N_XI54/XI8/NET35_XI54/XI8/MM11_g
+ N_VDD_XI54/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI9/MM2 N_XI54/XI9/NET34_XI54/XI9/MM2_d N_XI54/XI9/NET33_XI54/XI9/MM2_g
+ N_VSS_XI54/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM3 N_XI54/XI9/NET33_XI54/XI9/MM3_d N_WL<104>_XI54/XI9/MM3_g
+ N_BLN<6>_XI54/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM0 N_XI54/XI9/NET34_XI54/XI9/MM0_d N_WL<104>_XI54/XI9/MM0_g
+ N_BL<6>_XI54/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM1 N_XI54/XI9/NET33_XI54/XI9/MM1_d N_XI54/XI9/NET34_XI54/XI9/MM1_g
+ N_VSS_XI54/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM9 N_XI54/XI9/NET36_XI54/XI9/MM9_d N_WL<105>_XI54/XI9/MM9_g
+ N_BL<6>_XI54/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM6 N_XI54/XI9/NET35_XI54/XI9/MM6_d N_XI54/XI9/NET36_XI54/XI9/MM6_g
+ N_VSS_XI54/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM7 N_XI54/XI9/NET36_XI54/XI9/MM7_d N_XI54/XI9/NET35_XI54/XI9/MM7_g
+ N_VSS_XI54/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM8 N_XI54/XI9/NET35_XI54/XI9/MM8_d N_WL<105>_XI54/XI9/MM8_g
+ N_BLN<6>_XI54/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI9/MM5 N_XI54/XI9/NET34_XI54/XI9/MM5_d N_XI54/XI9/NET33_XI54/XI9/MM5_g
+ N_VDD_XI54/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI9/MM4 N_XI54/XI9/NET33_XI54/XI9/MM4_d N_XI54/XI9/NET34_XI54/XI9/MM4_g
+ N_VDD_XI54/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI9/MM10 N_XI54/XI9/NET35_XI54/XI9/MM10_d N_XI54/XI9/NET36_XI54/XI9/MM10_g
+ N_VDD_XI54/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI9/MM11 N_XI54/XI9/NET36_XI54/XI9/MM11_d N_XI54/XI9/NET35_XI54/XI9/MM11_g
+ N_VDD_XI54/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI10/MM2 N_XI54/XI10/NET34_XI54/XI10/MM2_d
+ N_XI54/XI10/NET33_XI54/XI10/MM2_g N_VSS_XI54/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI10/MM3 N_XI54/XI10/NET33_XI54/XI10/MM3_d N_WL<104>_XI54/XI10/MM3_g
+ N_BLN<5>_XI54/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI10/MM0 N_XI54/XI10/NET34_XI54/XI10/MM0_d N_WL<104>_XI54/XI10/MM0_g
+ N_BL<5>_XI54/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI10/MM1 N_XI54/XI10/NET33_XI54/XI10/MM1_d
+ N_XI54/XI10/NET34_XI54/XI10/MM1_g N_VSS_XI54/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI10/MM9 N_XI54/XI10/NET36_XI54/XI10/MM9_d N_WL<105>_XI54/XI10/MM9_g
+ N_BL<5>_XI54/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI10/MM6 N_XI54/XI10/NET35_XI54/XI10/MM6_d
+ N_XI54/XI10/NET36_XI54/XI10/MM6_g N_VSS_XI54/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI10/MM7 N_XI54/XI10/NET36_XI54/XI10/MM7_d
+ N_XI54/XI10/NET35_XI54/XI10/MM7_g N_VSS_XI54/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI10/MM8 N_XI54/XI10/NET35_XI54/XI10/MM8_d N_WL<105>_XI54/XI10/MM8_g
+ N_BLN<5>_XI54/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI10/MM5 N_XI54/XI10/NET34_XI54/XI10/MM5_d
+ N_XI54/XI10/NET33_XI54/XI10/MM5_g N_VDD_XI54/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI10/MM4 N_XI54/XI10/NET33_XI54/XI10/MM4_d
+ N_XI54/XI10/NET34_XI54/XI10/MM4_g N_VDD_XI54/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI10/MM10 N_XI54/XI10/NET35_XI54/XI10/MM10_d
+ N_XI54/XI10/NET36_XI54/XI10/MM10_g N_VDD_XI54/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI10/MM11 N_XI54/XI10/NET36_XI54/XI10/MM11_d
+ N_XI54/XI10/NET35_XI54/XI10/MM11_g N_VDD_XI54/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI11/MM2 N_XI54/XI11/NET34_XI54/XI11/MM2_d
+ N_XI54/XI11/NET33_XI54/XI11/MM2_g N_VSS_XI54/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI11/MM3 N_XI54/XI11/NET33_XI54/XI11/MM3_d N_WL<104>_XI54/XI11/MM3_g
+ N_BLN<4>_XI54/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI11/MM0 N_XI54/XI11/NET34_XI54/XI11/MM0_d N_WL<104>_XI54/XI11/MM0_g
+ N_BL<4>_XI54/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI11/MM1 N_XI54/XI11/NET33_XI54/XI11/MM1_d
+ N_XI54/XI11/NET34_XI54/XI11/MM1_g N_VSS_XI54/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI11/MM9 N_XI54/XI11/NET36_XI54/XI11/MM9_d N_WL<105>_XI54/XI11/MM9_g
+ N_BL<4>_XI54/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI11/MM6 N_XI54/XI11/NET35_XI54/XI11/MM6_d
+ N_XI54/XI11/NET36_XI54/XI11/MM6_g N_VSS_XI54/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI11/MM7 N_XI54/XI11/NET36_XI54/XI11/MM7_d
+ N_XI54/XI11/NET35_XI54/XI11/MM7_g N_VSS_XI54/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI11/MM8 N_XI54/XI11/NET35_XI54/XI11/MM8_d N_WL<105>_XI54/XI11/MM8_g
+ N_BLN<4>_XI54/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI11/MM5 N_XI54/XI11/NET34_XI54/XI11/MM5_d
+ N_XI54/XI11/NET33_XI54/XI11/MM5_g N_VDD_XI54/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI11/MM4 N_XI54/XI11/NET33_XI54/XI11/MM4_d
+ N_XI54/XI11/NET34_XI54/XI11/MM4_g N_VDD_XI54/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI11/MM10 N_XI54/XI11/NET35_XI54/XI11/MM10_d
+ N_XI54/XI11/NET36_XI54/XI11/MM10_g N_VDD_XI54/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI11/MM11 N_XI54/XI11/NET36_XI54/XI11/MM11_d
+ N_XI54/XI11/NET35_XI54/XI11/MM11_g N_VDD_XI54/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI12/MM2 N_XI54/XI12/NET34_XI54/XI12/MM2_d
+ N_XI54/XI12/NET33_XI54/XI12/MM2_g N_VSS_XI54/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI12/MM3 N_XI54/XI12/NET33_XI54/XI12/MM3_d N_WL<104>_XI54/XI12/MM3_g
+ N_BLN<3>_XI54/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI12/MM0 N_XI54/XI12/NET34_XI54/XI12/MM0_d N_WL<104>_XI54/XI12/MM0_g
+ N_BL<3>_XI54/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI12/MM1 N_XI54/XI12/NET33_XI54/XI12/MM1_d
+ N_XI54/XI12/NET34_XI54/XI12/MM1_g N_VSS_XI54/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI12/MM9 N_XI54/XI12/NET36_XI54/XI12/MM9_d N_WL<105>_XI54/XI12/MM9_g
+ N_BL<3>_XI54/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI12/MM6 N_XI54/XI12/NET35_XI54/XI12/MM6_d
+ N_XI54/XI12/NET36_XI54/XI12/MM6_g N_VSS_XI54/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI12/MM7 N_XI54/XI12/NET36_XI54/XI12/MM7_d
+ N_XI54/XI12/NET35_XI54/XI12/MM7_g N_VSS_XI54/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI12/MM8 N_XI54/XI12/NET35_XI54/XI12/MM8_d N_WL<105>_XI54/XI12/MM8_g
+ N_BLN<3>_XI54/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI12/MM5 N_XI54/XI12/NET34_XI54/XI12/MM5_d
+ N_XI54/XI12/NET33_XI54/XI12/MM5_g N_VDD_XI54/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI12/MM4 N_XI54/XI12/NET33_XI54/XI12/MM4_d
+ N_XI54/XI12/NET34_XI54/XI12/MM4_g N_VDD_XI54/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI12/MM10 N_XI54/XI12/NET35_XI54/XI12/MM10_d
+ N_XI54/XI12/NET36_XI54/XI12/MM10_g N_VDD_XI54/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI12/MM11 N_XI54/XI12/NET36_XI54/XI12/MM11_d
+ N_XI54/XI12/NET35_XI54/XI12/MM11_g N_VDD_XI54/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI13/MM2 N_XI54/XI13/NET34_XI54/XI13/MM2_d
+ N_XI54/XI13/NET33_XI54/XI13/MM2_g N_VSS_XI54/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI13/MM3 N_XI54/XI13/NET33_XI54/XI13/MM3_d N_WL<104>_XI54/XI13/MM3_g
+ N_BLN<2>_XI54/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI13/MM0 N_XI54/XI13/NET34_XI54/XI13/MM0_d N_WL<104>_XI54/XI13/MM0_g
+ N_BL<2>_XI54/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI13/MM1 N_XI54/XI13/NET33_XI54/XI13/MM1_d
+ N_XI54/XI13/NET34_XI54/XI13/MM1_g N_VSS_XI54/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI13/MM9 N_XI54/XI13/NET36_XI54/XI13/MM9_d N_WL<105>_XI54/XI13/MM9_g
+ N_BL<2>_XI54/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI13/MM6 N_XI54/XI13/NET35_XI54/XI13/MM6_d
+ N_XI54/XI13/NET36_XI54/XI13/MM6_g N_VSS_XI54/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI13/MM7 N_XI54/XI13/NET36_XI54/XI13/MM7_d
+ N_XI54/XI13/NET35_XI54/XI13/MM7_g N_VSS_XI54/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI13/MM8 N_XI54/XI13/NET35_XI54/XI13/MM8_d N_WL<105>_XI54/XI13/MM8_g
+ N_BLN<2>_XI54/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI13/MM5 N_XI54/XI13/NET34_XI54/XI13/MM5_d
+ N_XI54/XI13/NET33_XI54/XI13/MM5_g N_VDD_XI54/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI13/MM4 N_XI54/XI13/NET33_XI54/XI13/MM4_d
+ N_XI54/XI13/NET34_XI54/XI13/MM4_g N_VDD_XI54/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI13/MM10 N_XI54/XI13/NET35_XI54/XI13/MM10_d
+ N_XI54/XI13/NET36_XI54/XI13/MM10_g N_VDD_XI54/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI13/MM11 N_XI54/XI13/NET36_XI54/XI13/MM11_d
+ N_XI54/XI13/NET35_XI54/XI13/MM11_g N_VDD_XI54/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI14/MM2 N_XI54/XI14/NET34_XI54/XI14/MM2_d
+ N_XI54/XI14/NET33_XI54/XI14/MM2_g N_VSS_XI54/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI14/MM3 N_XI54/XI14/NET33_XI54/XI14/MM3_d N_WL<104>_XI54/XI14/MM3_g
+ N_BLN<1>_XI54/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI14/MM0 N_XI54/XI14/NET34_XI54/XI14/MM0_d N_WL<104>_XI54/XI14/MM0_g
+ N_BL<1>_XI54/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI14/MM1 N_XI54/XI14/NET33_XI54/XI14/MM1_d
+ N_XI54/XI14/NET34_XI54/XI14/MM1_g N_VSS_XI54/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI14/MM9 N_XI54/XI14/NET36_XI54/XI14/MM9_d N_WL<105>_XI54/XI14/MM9_g
+ N_BL<1>_XI54/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI14/MM6 N_XI54/XI14/NET35_XI54/XI14/MM6_d
+ N_XI54/XI14/NET36_XI54/XI14/MM6_g N_VSS_XI54/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI14/MM7 N_XI54/XI14/NET36_XI54/XI14/MM7_d
+ N_XI54/XI14/NET35_XI54/XI14/MM7_g N_VSS_XI54/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI14/MM8 N_XI54/XI14/NET35_XI54/XI14/MM8_d N_WL<105>_XI54/XI14/MM8_g
+ N_BLN<1>_XI54/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI14/MM5 N_XI54/XI14/NET34_XI54/XI14/MM5_d
+ N_XI54/XI14/NET33_XI54/XI14/MM5_g N_VDD_XI54/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI14/MM4 N_XI54/XI14/NET33_XI54/XI14/MM4_d
+ N_XI54/XI14/NET34_XI54/XI14/MM4_g N_VDD_XI54/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI14/MM10 N_XI54/XI14/NET35_XI54/XI14/MM10_d
+ N_XI54/XI14/NET36_XI54/XI14/MM10_g N_VDD_XI54/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI14/MM11 N_XI54/XI14/NET36_XI54/XI14/MM11_d
+ N_XI54/XI14/NET35_XI54/XI14/MM11_g N_VDD_XI54/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI15/MM2 N_XI54/XI15/NET34_XI54/XI15/MM2_d
+ N_XI54/XI15/NET33_XI54/XI15/MM2_g N_VSS_XI54/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI15/MM3 N_XI54/XI15/NET33_XI54/XI15/MM3_d N_WL<104>_XI54/XI15/MM3_g
+ N_BLN<0>_XI54/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI15/MM0 N_XI54/XI15/NET34_XI54/XI15/MM0_d N_WL<104>_XI54/XI15/MM0_g
+ N_BL<0>_XI54/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI15/MM1 N_XI54/XI15/NET33_XI54/XI15/MM1_d
+ N_XI54/XI15/NET34_XI54/XI15/MM1_g N_VSS_XI54/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI15/MM9 N_XI54/XI15/NET36_XI54/XI15/MM9_d N_WL<105>_XI54/XI15/MM9_g
+ N_BL<0>_XI54/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI15/MM6 N_XI54/XI15/NET35_XI54/XI15/MM6_d
+ N_XI54/XI15/NET36_XI54/XI15/MM6_g N_VSS_XI54/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI15/MM7 N_XI54/XI15/NET36_XI54/XI15/MM7_d
+ N_XI54/XI15/NET35_XI54/XI15/MM7_g N_VSS_XI54/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI54/XI15/MM8 N_XI54/XI15/NET35_XI54/XI15/MM8_d N_WL<105>_XI54/XI15/MM8_g
+ N_BLN<0>_XI54/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI54/XI15/MM5 N_XI54/XI15/NET34_XI54/XI15/MM5_d
+ N_XI54/XI15/NET33_XI54/XI15/MM5_g N_VDD_XI54/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI15/MM4 N_XI54/XI15/NET33_XI54/XI15/MM4_d
+ N_XI54/XI15/NET34_XI54/XI15/MM4_g N_VDD_XI54/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI15/MM10 N_XI54/XI15/NET35_XI54/XI15/MM10_d
+ N_XI54/XI15/NET36_XI54/XI15/MM10_g N_VDD_XI54/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI54/XI15/MM11 N_XI54/XI15/NET36_XI54/XI15/MM11_d
+ N_XI54/XI15/NET35_XI54/XI15/MM11_g N_VDD_XI54/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI0/MM2 N_XI55/XI0/NET34_XI55/XI0/MM2_d N_XI55/XI0/NET33_XI55/XI0/MM2_g
+ N_VSS_XI55/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI0/MM3 N_XI55/XI0/NET33_XI55/XI0/MM3_d N_WL<106>_XI55/XI0/MM3_g
+ N_BLN<15>_XI55/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI0/MM0 N_XI55/XI0/NET34_XI55/XI0/MM0_d N_WL<106>_XI55/XI0/MM0_g
+ N_BL<15>_XI55/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI0/MM1 N_XI55/XI0/NET33_XI55/XI0/MM1_d N_XI55/XI0/NET34_XI55/XI0/MM1_g
+ N_VSS_XI55/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI0/MM9 N_XI55/XI0/NET36_XI55/XI0/MM9_d N_WL<107>_XI55/XI0/MM9_g
+ N_BL<15>_XI55/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI0/MM6 N_XI55/XI0/NET35_XI55/XI0/MM6_d N_XI55/XI0/NET36_XI55/XI0/MM6_g
+ N_VSS_XI55/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI0/MM7 N_XI55/XI0/NET36_XI55/XI0/MM7_d N_XI55/XI0/NET35_XI55/XI0/MM7_g
+ N_VSS_XI55/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI0/MM8 N_XI55/XI0/NET35_XI55/XI0/MM8_d N_WL<107>_XI55/XI0/MM8_g
+ N_BLN<15>_XI55/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI0/MM5 N_XI55/XI0/NET34_XI55/XI0/MM5_d N_XI55/XI0/NET33_XI55/XI0/MM5_g
+ N_VDD_XI55/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI0/MM4 N_XI55/XI0/NET33_XI55/XI0/MM4_d N_XI55/XI0/NET34_XI55/XI0/MM4_g
+ N_VDD_XI55/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI0/MM10 N_XI55/XI0/NET35_XI55/XI0/MM10_d N_XI55/XI0/NET36_XI55/XI0/MM10_g
+ N_VDD_XI55/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI0/MM11 N_XI55/XI0/NET36_XI55/XI0/MM11_d N_XI55/XI0/NET35_XI55/XI0/MM11_g
+ N_VDD_XI55/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI1/MM2 N_XI55/XI1/NET34_XI55/XI1/MM2_d N_XI55/XI1/NET33_XI55/XI1/MM2_g
+ N_VSS_XI55/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI1/MM3 N_XI55/XI1/NET33_XI55/XI1/MM3_d N_WL<106>_XI55/XI1/MM3_g
+ N_BLN<14>_XI55/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI1/MM0 N_XI55/XI1/NET34_XI55/XI1/MM0_d N_WL<106>_XI55/XI1/MM0_g
+ N_BL<14>_XI55/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI1/MM1 N_XI55/XI1/NET33_XI55/XI1/MM1_d N_XI55/XI1/NET34_XI55/XI1/MM1_g
+ N_VSS_XI55/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI1/MM9 N_XI55/XI1/NET36_XI55/XI1/MM9_d N_WL<107>_XI55/XI1/MM9_g
+ N_BL<14>_XI55/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI1/MM6 N_XI55/XI1/NET35_XI55/XI1/MM6_d N_XI55/XI1/NET36_XI55/XI1/MM6_g
+ N_VSS_XI55/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI1/MM7 N_XI55/XI1/NET36_XI55/XI1/MM7_d N_XI55/XI1/NET35_XI55/XI1/MM7_g
+ N_VSS_XI55/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI1/MM8 N_XI55/XI1/NET35_XI55/XI1/MM8_d N_WL<107>_XI55/XI1/MM8_g
+ N_BLN<14>_XI55/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI1/MM5 N_XI55/XI1/NET34_XI55/XI1/MM5_d N_XI55/XI1/NET33_XI55/XI1/MM5_g
+ N_VDD_XI55/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI1/MM4 N_XI55/XI1/NET33_XI55/XI1/MM4_d N_XI55/XI1/NET34_XI55/XI1/MM4_g
+ N_VDD_XI55/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI1/MM10 N_XI55/XI1/NET35_XI55/XI1/MM10_d N_XI55/XI1/NET36_XI55/XI1/MM10_g
+ N_VDD_XI55/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI1/MM11 N_XI55/XI1/NET36_XI55/XI1/MM11_d N_XI55/XI1/NET35_XI55/XI1/MM11_g
+ N_VDD_XI55/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI2/MM2 N_XI55/XI2/NET34_XI55/XI2/MM2_d N_XI55/XI2/NET33_XI55/XI2/MM2_g
+ N_VSS_XI55/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI2/MM3 N_XI55/XI2/NET33_XI55/XI2/MM3_d N_WL<106>_XI55/XI2/MM3_g
+ N_BLN<13>_XI55/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI2/MM0 N_XI55/XI2/NET34_XI55/XI2/MM0_d N_WL<106>_XI55/XI2/MM0_g
+ N_BL<13>_XI55/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI2/MM1 N_XI55/XI2/NET33_XI55/XI2/MM1_d N_XI55/XI2/NET34_XI55/XI2/MM1_g
+ N_VSS_XI55/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI2/MM9 N_XI55/XI2/NET36_XI55/XI2/MM9_d N_WL<107>_XI55/XI2/MM9_g
+ N_BL<13>_XI55/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI2/MM6 N_XI55/XI2/NET35_XI55/XI2/MM6_d N_XI55/XI2/NET36_XI55/XI2/MM6_g
+ N_VSS_XI55/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI2/MM7 N_XI55/XI2/NET36_XI55/XI2/MM7_d N_XI55/XI2/NET35_XI55/XI2/MM7_g
+ N_VSS_XI55/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI2/MM8 N_XI55/XI2/NET35_XI55/XI2/MM8_d N_WL<107>_XI55/XI2/MM8_g
+ N_BLN<13>_XI55/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI2/MM5 N_XI55/XI2/NET34_XI55/XI2/MM5_d N_XI55/XI2/NET33_XI55/XI2/MM5_g
+ N_VDD_XI55/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI2/MM4 N_XI55/XI2/NET33_XI55/XI2/MM4_d N_XI55/XI2/NET34_XI55/XI2/MM4_g
+ N_VDD_XI55/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI2/MM10 N_XI55/XI2/NET35_XI55/XI2/MM10_d N_XI55/XI2/NET36_XI55/XI2/MM10_g
+ N_VDD_XI55/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI2/MM11 N_XI55/XI2/NET36_XI55/XI2/MM11_d N_XI55/XI2/NET35_XI55/XI2/MM11_g
+ N_VDD_XI55/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI3/MM2 N_XI55/XI3/NET34_XI55/XI3/MM2_d N_XI55/XI3/NET33_XI55/XI3/MM2_g
+ N_VSS_XI55/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI3/MM3 N_XI55/XI3/NET33_XI55/XI3/MM3_d N_WL<106>_XI55/XI3/MM3_g
+ N_BLN<12>_XI55/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI3/MM0 N_XI55/XI3/NET34_XI55/XI3/MM0_d N_WL<106>_XI55/XI3/MM0_g
+ N_BL<12>_XI55/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI3/MM1 N_XI55/XI3/NET33_XI55/XI3/MM1_d N_XI55/XI3/NET34_XI55/XI3/MM1_g
+ N_VSS_XI55/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI3/MM9 N_XI55/XI3/NET36_XI55/XI3/MM9_d N_WL<107>_XI55/XI3/MM9_g
+ N_BL<12>_XI55/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI3/MM6 N_XI55/XI3/NET35_XI55/XI3/MM6_d N_XI55/XI3/NET36_XI55/XI3/MM6_g
+ N_VSS_XI55/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI3/MM7 N_XI55/XI3/NET36_XI55/XI3/MM7_d N_XI55/XI3/NET35_XI55/XI3/MM7_g
+ N_VSS_XI55/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI3/MM8 N_XI55/XI3/NET35_XI55/XI3/MM8_d N_WL<107>_XI55/XI3/MM8_g
+ N_BLN<12>_XI55/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI3/MM5 N_XI55/XI3/NET34_XI55/XI3/MM5_d N_XI55/XI3/NET33_XI55/XI3/MM5_g
+ N_VDD_XI55/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI3/MM4 N_XI55/XI3/NET33_XI55/XI3/MM4_d N_XI55/XI3/NET34_XI55/XI3/MM4_g
+ N_VDD_XI55/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI3/MM10 N_XI55/XI3/NET35_XI55/XI3/MM10_d N_XI55/XI3/NET36_XI55/XI3/MM10_g
+ N_VDD_XI55/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI3/MM11 N_XI55/XI3/NET36_XI55/XI3/MM11_d N_XI55/XI3/NET35_XI55/XI3/MM11_g
+ N_VDD_XI55/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI4/MM2 N_XI55/XI4/NET34_XI55/XI4/MM2_d N_XI55/XI4/NET33_XI55/XI4/MM2_g
+ N_VSS_XI55/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI4/MM3 N_XI55/XI4/NET33_XI55/XI4/MM3_d N_WL<106>_XI55/XI4/MM3_g
+ N_BLN<11>_XI55/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI4/MM0 N_XI55/XI4/NET34_XI55/XI4/MM0_d N_WL<106>_XI55/XI4/MM0_g
+ N_BL<11>_XI55/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI4/MM1 N_XI55/XI4/NET33_XI55/XI4/MM1_d N_XI55/XI4/NET34_XI55/XI4/MM1_g
+ N_VSS_XI55/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI4/MM9 N_XI55/XI4/NET36_XI55/XI4/MM9_d N_WL<107>_XI55/XI4/MM9_g
+ N_BL<11>_XI55/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI4/MM6 N_XI55/XI4/NET35_XI55/XI4/MM6_d N_XI55/XI4/NET36_XI55/XI4/MM6_g
+ N_VSS_XI55/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI4/MM7 N_XI55/XI4/NET36_XI55/XI4/MM7_d N_XI55/XI4/NET35_XI55/XI4/MM7_g
+ N_VSS_XI55/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI4/MM8 N_XI55/XI4/NET35_XI55/XI4/MM8_d N_WL<107>_XI55/XI4/MM8_g
+ N_BLN<11>_XI55/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI4/MM5 N_XI55/XI4/NET34_XI55/XI4/MM5_d N_XI55/XI4/NET33_XI55/XI4/MM5_g
+ N_VDD_XI55/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI4/MM4 N_XI55/XI4/NET33_XI55/XI4/MM4_d N_XI55/XI4/NET34_XI55/XI4/MM4_g
+ N_VDD_XI55/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI4/MM10 N_XI55/XI4/NET35_XI55/XI4/MM10_d N_XI55/XI4/NET36_XI55/XI4/MM10_g
+ N_VDD_XI55/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI4/MM11 N_XI55/XI4/NET36_XI55/XI4/MM11_d N_XI55/XI4/NET35_XI55/XI4/MM11_g
+ N_VDD_XI55/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI5/MM2 N_XI55/XI5/NET34_XI55/XI5/MM2_d N_XI55/XI5/NET33_XI55/XI5/MM2_g
+ N_VSS_XI55/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI5/MM3 N_XI55/XI5/NET33_XI55/XI5/MM3_d N_WL<106>_XI55/XI5/MM3_g
+ N_BLN<10>_XI55/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI5/MM0 N_XI55/XI5/NET34_XI55/XI5/MM0_d N_WL<106>_XI55/XI5/MM0_g
+ N_BL<10>_XI55/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI5/MM1 N_XI55/XI5/NET33_XI55/XI5/MM1_d N_XI55/XI5/NET34_XI55/XI5/MM1_g
+ N_VSS_XI55/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI5/MM9 N_XI55/XI5/NET36_XI55/XI5/MM9_d N_WL<107>_XI55/XI5/MM9_g
+ N_BL<10>_XI55/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI5/MM6 N_XI55/XI5/NET35_XI55/XI5/MM6_d N_XI55/XI5/NET36_XI55/XI5/MM6_g
+ N_VSS_XI55/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI5/MM7 N_XI55/XI5/NET36_XI55/XI5/MM7_d N_XI55/XI5/NET35_XI55/XI5/MM7_g
+ N_VSS_XI55/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI5/MM8 N_XI55/XI5/NET35_XI55/XI5/MM8_d N_WL<107>_XI55/XI5/MM8_g
+ N_BLN<10>_XI55/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI5/MM5 N_XI55/XI5/NET34_XI55/XI5/MM5_d N_XI55/XI5/NET33_XI55/XI5/MM5_g
+ N_VDD_XI55/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI5/MM4 N_XI55/XI5/NET33_XI55/XI5/MM4_d N_XI55/XI5/NET34_XI55/XI5/MM4_g
+ N_VDD_XI55/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI5/MM10 N_XI55/XI5/NET35_XI55/XI5/MM10_d N_XI55/XI5/NET36_XI55/XI5/MM10_g
+ N_VDD_XI55/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI5/MM11 N_XI55/XI5/NET36_XI55/XI5/MM11_d N_XI55/XI5/NET35_XI55/XI5/MM11_g
+ N_VDD_XI55/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI6/MM2 N_XI55/XI6/NET34_XI55/XI6/MM2_d N_XI55/XI6/NET33_XI55/XI6/MM2_g
+ N_VSS_XI55/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM3 N_XI55/XI6/NET33_XI55/XI6/MM3_d N_WL<106>_XI55/XI6/MM3_g
+ N_BLN<9>_XI55/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM0 N_XI55/XI6/NET34_XI55/XI6/MM0_d N_WL<106>_XI55/XI6/MM0_g
+ N_BL<9>_XI55/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM1 N_XI55/XI6/NET33_XI55/XI6/MM1_d N_XI55/XI6/NET34_XI55/XI6/MM1_g
+ N_VSS_XI55/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM9 N_XI55/XI6/NET36_XI55/XI6/MM9_d N_WL<107>_XI55/XI6/MM9_g
+ N_BL<9>_XI55/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM6 N_XI55/XI6/NET35_XI55/XI6/MM6_d N_XI55/XI6/NET36_XI55/XI6/MM6_g
+ N_VSS_XI55/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM7 N_XI55/XI6/NET36_XI55/XI6/MM7_d N_XI55/XI6/NET35_XI55/XI6/MM7_g
+ N_VSS_XI55/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM8 N_XI55/XI6/NET35_XI55/XI6/MM8_d N_WL<107>_XI55/XI6/MM8_g
+ N_BLN<9>_XI55/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI6/MM5 N_XI55/XI6/NET34_XI55/XI6/MM5_d N_XI55/XI6/NET33_XI55/XI6/MM5_g
+ N_VDD_XI55/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI6/MM4 N_XI55/XI6/NET33_XI55/XI6/MM4_d N_XI55/XI6/NET34_XI55/XI6/MM4_g
+ N_VDD_XI55/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI6/MM10 N_XI55/XI6/NET35_XI55/XI6/MM10_d N_XI55/XI6/NET36_XI55/XI6/MM10_g
+ N_VDD_XI55/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI6/MM11 N_XI55/XI6/NET36_XI55/XI6/MM11_d N_XI55/XI6/NET35_XI55/XI6/MM11_g
+ N_VDD_XI55/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI7/MM2 N_XI55/XI7/NET34_XI55/XI7/MM2_d N_XI55/XI7/NET33_XI55/XI7/MM2_g
+ N_VSS_XI55/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM3 N_XI55/XI7/NET33_XI55/XI7/MM3_d N_WL<106>_XI55/XI7/MM3_g
+ N_BLN<8>_XI55/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM0 N_XI55/XI7/NET34_XI55/XI7/MM0_d N_WL<106>_XI55/XI7/MM0_g
+ N_BL<8>_XI55/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM1 N_XI55/XI7/NET33_XI55/XI7/MM1_d N_XI55/XI7/NET34_XI55/XI7/MM1_g
+ N_VSS_XI55/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM9 N_XI55/XI7/NET36_XI55/XI7/MM9_d N_WL<107>_XI55/XI7/MM9_g
+ N_BL<8>_XI55/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM6 N_XI55/XI7/NET35_XI55/XI7/MM6_d N_XI55/XI7/NET36_XI55/XI7/MM6_g
+ N_VSS_XI55/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM7 N_XI55/XI7/NET36_XI55/XI7/MM7_d N_XI55/XI7/NET35_XI55/XI7/MM7_g
+ N_VSS_XI55/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM8 N_XI55/XI7/NET35_XI55/XI7/MM8_d N_WL<107>_XI55/XI7/MM8_g
+ N_BLN<8>_XI55/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI7/MM5 N_XI55/XI7/NET34_XI55/XI7/MM5_d N_XI55/XI7/NET33_XI55/XI7/MM5_g
+ N_VDD_XI55/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI7/MM4 N_XI55/XI7/NET33_XI55/XI7/MM4_d N_XI55/XI7/NET34_XI55/XI7/MM4_g
+ N_VDD_XI55/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI7/MM10 N_XI55/XI7/NET35_XI55/XI7/MM10_d N_XI55/XI7/NET36_XI55/XI7/MM10_g
+ N_VDD_XI55/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI7/MM11 N_XI55/XI7/NET36_XI55/XI7/MM11_d N_XI55/XI7/NET35_XI55/XI7/MM11_g
+ N_VDD_XI55/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI8/MM2 N_XI55/XI8/NET34_XI55/XI8/MM2_d N_XI55/XI8/NET33_XI55/XI8/MM2_g
+ N_VSS_XI55/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM3 N_XI55/XI8/NET33_XI55/XI8/MM3_d N_WL<106>_XI55/XI8/MM3_g
+ N_BLN<7>_XI55/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM0 N_XI55/XI8/NET34_XI55/XI8/MM0_d N_WL<106>_XI55/XI8/MM0_g
+ N_BL<7>_XI55/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM1 N_XI55/XI8/NET33_XI55/XI8/MM1_d N_XI55/XI8/NET34_XI55/XI8/MM1_g
+ N_VSS_XI55/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM9 N_XI55/XI8/NET36_XI55/XI8/MM9_d N_WL<107>_XI55/XI8/MM9_g
+ N_BL<7>_XI55/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM6 N_XI55/XI8/NET35_XI55/XI8/MM6_d N_XI55/XI8/NET36_XI55/XI8/MM6_g
+ N_VSS_XI55/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM7 N_XI55/XI8/NET36_XI55/XI8/MM7_d N_XI55/XI8/NET35_XI55/XI8/MM7_g
+ N_VSS_XI55/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM8 N_XI55/XI8/NET35_XI55/XI8/MM8_d N_WL<107>_XI55/XI8/MM8_g
+ N_BLN<7>_XI55/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI8/MM5 N_XI55/XI8/NET34_XI55/XI8/MM5_d N_XI55/XI8/NET33_XI55/XI8/MM5_g
+ N_VDD_XI55/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI8/MM4 N_XI55/XI8/NET33_XI55/XI8/MM4_d N_XI55/XI8/NET34_XI55/XI8/MM4_g
+ N_VDD_XI55/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI8/MM10 N_XI55/XI8/NET35_XI55/XI8/MM10_d N_XI55/XI8/NET36_XI55/XI8/MM10_g
+ N_VDD_XI55/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI8/MM11 N_XI55/XI8/NET36_XI55/XI8/MM11_d N_XI55/XI8/NET35_XI55/XI8/MM11_g
+ N_VDD_XI55/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI9/MM2 N_XI55/XI9/NET34_XI55/XI9/MM2_d N_XI55/XI9/NET33_XI55/XI9/MM2_g
+ N_VSS_XI55/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM3 N_XI55/XI9/NET33_XI55/XI9/MM3_d N_WL<106>_XI55/XI9/MM3_g
+ N_BLN<6>_XI55/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM0 N_XI55/XI9/NET34_XI55/XI9/MM0_d N_WL<106>_XI55/XI9/MM0_g
+ N_BL<6>_XI55/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM1 N_XI55/XI9/NET33_XI55/XI9/MM1_d N_XI55/XI9/NET34_XI55/XI9/MM1_g
+ N_VSS_XI55/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM9 N_XI55/XI9/NET36_XI55/XI9/MM9_d N_WL<107>_XI55/XI9/MM9_g
+ N_BL<6>_XI55/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM6 N_XI55/XI9/NET35_XI55/XI9/MM6_d N_XI55/XI9/NET36_XI55/XI9/MM6_g
+ N_VSS_XI55/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM7 N_XI55/XI9/NET36_XI55/XI9/MM7_d N_XI55/XI9/NET35_XI55/XI9/MM7_g
+ N_VSS_XI55/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM8 N_XI55/XI9/NET35_XI55/XI9/MM8_d N_WL<107>_XI55/XI9/MM8_g
+ N_BLN<6>_XI55/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI9/MM5 N_XI55/XI9/NET34_XI55/XI9/MM5_d N_XI55/XI9/NET33_XI55/XI9/MM5_g
+ N_VDD_XI55/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI9/MM4 N_XI55/XI9/NET33_XI55/XI9/MM4_d N_XI55/XI9/NET34_XI55/XI9/MM4_g
+ N_VDD_XI55/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI9/MM10 N_XI55/XI9/NET35_XI55/XI9/MM10_d N_XI55/XI9/NET36_XI55/XI9/MM10_g
+ N_VDD_XI55/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI9/MM11 N_XI55/XI9/NET36_XI55/XI9/MM11_d N_XI55/XI9/NET35_XI55/XI9/MM11_g
+ N_VDD_XI55/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI10/MM2 N_XI55/XI10/NET34_XI55/XI10/MM2_d
+ N_XI55/XI10/NET33_XI55/XI10/MM2_g N_VSS_XI55/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI10/MM3 N_XI55/XI10/NET33_XI55/XI10/MM3_d N_WL<106>_XI55/XI10/MM3_g
+ N_BLN<5>_XI55/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI10/MM0 N_XI55/XI10/NET34_XI55/XI10/MM0_d N_WL<106>_XI55/XI10/MM0_g
+ N_BL<5>_XI55/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI10/MM1 N_XI55/XI10/NET33_XI55/XI10/MM1_d
+ N_XI55/XI10/NET34_XI55/XI10/MM1_g N_VSS_XI55/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI10/MM9 N_XI55/XI10/NET36_XI55/XI10/MM9_d N_WL<107>_XI55/XI10/MM9_g
+ N_BL<5>_XI55/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI10/MM6 N_XI55/XI10/NET35_XI55/XI10/MM6_d
+ N_XI55/XI10/NET36_XI55/XI10/MM6_g N_VSS_XI55/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI10/MM7 N_XI55/XI10/NET36_XI55/XI10/MM7_d
+ N_XI55/XI10/NET35_XI55/XI10/MM7_g N_VSS_XI55/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI10/MM8 N_XI55/XI10/NET35_XI55/XI10/MM8_d N_WL<107>_XI55/XI10/MM8_g
+ N_BLN<5>_XI55/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI10/MM5 N_XI55/XI10/NET34_XI55/XI10/MM5_d
+ N_XI55/XI10/NET33_XI55/XI10/MM5_g N_VDD_XI55/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI10/MM4 N_XI55/XI10/NET33_XI55/XI10/MM4_d
+ N_XI55/XI10/NET34_XI55/XI10/MM4_g N_VDD_XI55/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI10/MM10 N_XI55/XI10/NET35_XI55/XI10/MM10_d
+ N_XI55/XI10/NET36_XI55/XI10/MM10_g N_VDD_XI55/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI10/MM11 N_XI55/XI10/NET36_XI55/XI10/MM11_d
+ N_XI55/XI10/NET35_XI55/XI10/MM11_g N_VDD_XI55/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI11/MM2 N_XI55/XI11/NET34_XI55/XI11/MM2_d
+ N_XI55/XI11/NET33_XI55/XI11/MM2_g N_VSS_XI55/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI11/MM3 N_XI55/XI11/NET33_XI55/XI11/MM3_d N_WL<106>_XI55/XI11/MM3_g
+ N_BLN<4>_XI55/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI11/MM0 N_XI55/XI11/NET34_XI55/XI11/MM0_d N_WL<106>_XI55/XI11/MM0_g
+ N_BL<4>_XI55/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI11/MM1 N_XI55/XI11/NET33_XI55/XI11/MM1_d
+ N_XI55/XI11/NET34_XI55/XI11/MM1_g N_VSS_XI55/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI11/MM9 N_XI55/XI11/NET36_XI55/XI11/MM9_d N_WL<107>_XI55/XI11/MM9_g
+ N_BL<4>_XI55/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI11/MM6 N_XI55/XI11/NET35_XI55/XI11/MM6_d
+ N_XI55/XI11/NET36_XI55/XI11/MM6_g N_VSS_XI55/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI11/MM7 N_XI55/XI11/NET36_XI55/XI11/MM7_d
+ N_XI55/XI11/NET35_XI55/XI11/MM7_g N_VSS_XI55/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI11/MM8 N_XI55/XI11/NET35_XI55/XI11/MM8_d N_WL<107>_XI55/XI11/MM8_g
+ N_BLN<4>_XI55/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI11/MM5 N_XI55/XI11/NET34_XI55/XI11/MM5_d
+ N_XI55/XI11/NET33_XI55/XI11/MM5_g N_VDD_XI55/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI11/MM4 N_XI55/XI11/NET33_XI55/XI11/MM4_d
+ N_XI55/XI11/NET34_XI55/XI11/MM4_g N_VDD_XI55/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI11/MM10 N_XI55/XI11/NET35_XI55/XI11/MM10_d
+ N_XI55/XI11/NET36_XI55/XI11/MM10_g N_VDD_XI55/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI11/MM11 N_XI55/XI11/NET36_XI55/XI11/MM11_d
+ N_XI55/XI11/NET35_XI55/XI11/MM11_g N_VDD_XI55/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI12/MM2 N_XI55/XI12/NET34_XI55/XI12/MM2_d
+ N_XI55/XI12/NET33_XI55/XI12/MM2_g N_VSS_XI55/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI12/MM3 N_XI55/XI12/NET33_XI55/XI12/MM3_d N_WL<106>_XI55/XI12/MM3_g
+ N_BLN<3>_XI55/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI12/MM0 N_XI55/XI12/NET34_XI55/XI12/MM0_d N_WL<106>_XI55/XI12/MM0_g
+ N_BL<3>_XI55/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI12/MM1 N_XI55/XI12/NET33_XI55/XI12/MM1_d
+ N_XI55/XI12/NET34_XI55/XI12/MM1_g N_VSS_XI55/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI12/MM9 N_XI55/XI12/NET36_XI55/XI12/MM9_d N_WL<107>_XI55/XI12/MM9_g
+ N_BL<3>_XI55/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI12/MM6 N_XI55/XI12/NET35_XI55/XI12/MM6_d
+ N_XI55/XI12/NET36_XI55/XI12/MM6_g N_VSS_XI55/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI12/MM7 N_XI55/XI12/NET36_XI55/XI12/MM7_d
+ N_XI55/XI12/NET35_XI55/XI12/MM7_g N_VSS_XI55/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI12/MM8 N_XI55/XI12/NET35_XI55/XI12/MM8_d N_WL<107>_XI55/XI12/MM8_g
+ N_BLN<3>_XI55/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI12/MM5 N_XI55/XI12/NET34_XI55/XI12/MM5_d
+ N_XI55/XI12/NET33_XI55/XI12/MM5_g N_VDD_XI55/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI12/MM4 N_XI55/XI12/NET33_XI55/XI12/MM4_d
+ N_XI55/XI12/NET34_XI55/XI12/MM4_g N_VDD_XI55/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI12/MM10 N_XI55/XI12/NET35_XI55/XI12/MM10_d
+ N_XI55/XI12/NET36_XI55/XI12/MM10_g N_VDD_XI55/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI12/MM11 N_XI55/XI12/NET36_XI55/XI12/MM11_d
+ N_XI55/XI12/NET35_XI55/XI12/MM11_g N_VDD_XI55/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI13/MM2 N_XI55/XI13/NET34_XI55/XI13/MM2_d
+ N_XI55/XI13/NET33_XI55/XI13/MM2_g N_VSS_XI55/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI13/MM3 N_XI55/XI13/NET33_XI55/XI13/MM3_d N_WL<106>_XI55/XI13/MM3_g
+ N_BLN<2>_XI55/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI13/MM0 N_XI55/XI13/NET34_XI55/XI13/MM0_d N_WL<106>_XI55/XI13/MM0_g
+ N_BL<2>_XI55/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI13/MM1 N_XI55/XI13/NET33_XI55/XI13/MM1_d
+ N_XI55/XI13/NET34_XI55/XI13/MM1_g N_VSS_XI55/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI13/MM9 N_XI55/XI13/NET36_XI55/XI13/MM9_d N_WL<107>_XI55/XI13/MM9_g
+ N_BL<2>_XI55/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI13/MM6 N_XI55/XI13/NET35_XI55/XI13/MM6_d
+ N_XI55/XI13/NET36_XI55/XI13/MM6_g N_VSS_XI55/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI13/MM7 N_XI55/XI13/NET36_XI55/XI13/MM7_d
+ N_XI55/XI13/NET35_XI55/XI13/MM7_g N_VSS_XI55/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI13/MM8 N_XI55/XI13/NET35_XI55/XI13/MM8_d N_WL<107>_XI55/XI13/MM8_g
+ N_BLN<2>_XI55/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI13/MM5 N_XI55/XI13/NET34_XI55/XI13/MM5_d
+ N_XI55/XI13/NET33_XI55/XI13/MM5_g N_VDD_XI55/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI13/MM4 N_XI55/XI13/NET33_XI55/XI13/MM4_d
+ N_XI55/XI13/NET34_XI55/XI13/MM4_g N_VDD_XI55/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI13/MM10 N_XI55/XI13/NET35_XI55/XI13/MM10_d
+ N_XI55/XI13/NET36_XI55/XI13/MM10_g N_VDD_XI55/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI13/MM11 N_XI55/XI13/NET36_XI55/XI13/MM11_d
+ N_XI55/XI13/NET35_XI55/XI13/MM11_g N_VDD_XI55/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI14/MM2 N_XI55/XI14/NET34_XI55/XI14/MM2_d
+ N_XI55/XI14/NET33_XI55/XI14/MM2_g N_VSS_XI55/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI14/MM3 N_XI55/XI14/NET33_XI55/XI14/MM3_d N_WL<106>_XI55/XI14/MM3_g
+ N_BLN<1>_XI55/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI14/MM0 N_XI55/XI14/NET34_XI55/XI14/MM0_d N_WL<106>_XI55/XI14/MM0_g
+ N_BL<1>_XI55/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI14/MM1 N_XI55/XI14/NET33_XI55/XI14/MM1_d
+ N_XI55/XI14/NET34_XI55/XI14/MM1_g N_VSS_XI55/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI14/MM9 N_XI55/XI14/NET36_XI55/XI14/MM9_d N_WL<107>_XI55/XI14/MM9_g
+ N_BL<1>_XI55/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI14/MM6 N_XI55/XI14/NET35_XI55/XI14/MM6_d
+ N_XI55/XI14/NET36_XI55/XI14/MM6_g N_VSS_XI55/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI14/MM7 N_XI55/XI14/NET36_XI55/XI14/MM7_d
+ N_XI55/XI14/NET35_XI55/XI14/MM7_g N_VSS_XI55/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI14/MM8 N_XI55/XI14/NET35_XI55/XI14/MM8_d N_WL<107>_XI55/XI14/MM8_g
+ N_BLN<1>_XI55/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI14/MM5 N_XI55/XI14/NET34_XI55/XI14/MM5_d
+ N_XI55/XI14/NET33_XI55/XI14/MM5_g N_VDD_XI55/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI14/MM4 N_XI55/XI14/NET33_XI55/XI14/MM4_d
+ N_XI55/XI14/NET34_XI55/XI14/MM4_g N_VDD_XI55/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI14/MM10 N_XI55/XI14/NET35_XI55/XI14/MM10_d
+ N_XI55/XI14/NET36_XI55/XI14/MM10_g N_VDD_XI55/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI14/MM11 N_XI55/XI14/NET36_XI55/XI14/MM11_d
+ N_XI55/XI14/NET35_XI55/XI14/MM11_g N_VDD_XI55/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI15/MM2 N_XI55/XI15/NET34_XI55/XI15/MM2_d
+ N_XI55/XI15/NET33_XI55/XI15/MM2_g N_VSS_XI55/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI15/MM3 N_XI55/XI15/NET33_XI55/XI15/MM3_d N_WL<106>_XI55/XI15/MM3_g
+ N_BLN<0>_XI55/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI15/MM0 N_XI55/XI15/NET34_XI55/XI15/MM0_d N_WL<106>_XI55/XI15/MM0_g
+ N_BL<0>_XI55/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI15/MM1 N_XI55/XI15/NET33_XI55/XI15/MM1_d
+ N_XI55/XI15/NET34_XI55/XI15/MM1_g N_VSS_XI55/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI15/MM9 N_XI55/XI15/NET36_XI55/XI15/MM9_d N_WL<107>_XI55/XI15/MM9_g
+ N_BL<0>_XI55/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI15/MM6 N_XI55/XI15/NET35_XI55/XI15/MM6_d
+ N_XI55/XI15/NET36_XI55/XI15/MM6_g N_VSS_XI55/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI15/MM7 N_XI55/XI15/NET36_XI55/XI15/MM7_d
+ N_XI55/XI15/NET35_XI55/XI15/MM7_g N_VSS_XI55/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI55/XI15/MM8 N_XI55/XI15/NET35_XI55/XI15/MM8_d N_WL<107>_XI55/XI15/MM8_g
+ N_BLN<0>_XI55/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI55/XI15/MM5 N_XI55/XI15/NET34_XI55/XI15/MM5_d
+ N_XI55/XI15/NET33_XI55/XI15/MM5_g N_VDD_XI55/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI15/MM4 N_XI55/XI15/NET33_XI55/XI15/MM4_d
+ N_XI55/XI15/NET34_XI55/XI15/MM4_g N_VDD_XI55/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI15/MM10 N_XI55/XI15/NET35_XI55/XI15/MM10_d
+ N_XI55/XI15/NET36_XI55/XI15/MM10_g N_VDD_XI55/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI55/XI15/MM11 N_XI55/XI15/NET36_XI55/XI15/MM11_d
+ N_XI55/XI15/NET35_XI55/XI15/MM11_g N_VDD_XI55/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI0/MM2 N_XI56/XI0/NET34_XI56/XI0/MM2_d N_XI56/XI0/NET33_XI56/XI0/MM2_g
+ N_VSS_XI56/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI0/MM3 N_XI56/XI0/NET33_XI56/XI0/MM3_d N_WL<108>_XI56/XI0/MM3_g
+ N_BLN<15>_XI56/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI0/MM0 N_XI56/XI0/NET34_XI56/XI0/MM0_d N_WL<108>_XI56/XI0/MM0_g
+ N_BL<15>_XI56/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI0/MM1 N_XI56/XI0/NET33_XI56/XI0/MM1_d N_XI56/XI0/NET34_XI56/XI0/MM1_g
+ N_VSS_XI56/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI0/MM9 N_XI56/XI0/NET36_XI56/XI0/MM9_d N_WL<109>_XI56/XI0/MM9_g
+ N_BL<15>_XI56/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI0/MM6 N_XI56/XI0/NET35_XI56/XI0/MM6_d N_XI56/XI0/NET36_XI56/XI0/MM6_g
+ N_VSS_XI56/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI0/MM7 N_XI56/XI0/NET36_XI56/XI0/MM7_d N_XI56/XI0/NET35_XI56/XI0/MM7_g
+ N_VSS_XI56/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI0/MM8 N_XI56/XI0/NET35_XI56/XI0/MM8_d N_WL<109>_XI56/XI0/MM8_g
+ N_BLN<15>_XI56/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI0/MM5 N_XI56/XI0/NET34_XI56/XI0/MM5_d N_XI56/XI0/NET33_XI56/XI0/MM5_g
+ N_VDD_XI56/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI0/MM4 N_XI56/XI0/NET33_XI56/XI0/MM4_d N_XI56/XI0/NET34_XI56/XI0/MM4_g
+ N_VDD_XI56/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI0/MM10 N_XI56/XI0/NET35_XI56/XI0/MM10_d N_XI56/XI0/NET36_XI56/XI0/MM10_g
+ N_VDD_XI56/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI0/MM11 N_XI56/XI0/NET36_XI56/XI0/MM11_d N_XI56/XI0/NET35_XI56/XI0/MM11_g
+ N_VDD_XI56/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI1/MM2 N_XI56/XI1/NET34_XI56/XI1/MM2_d N_XI56/XI1/NET33_XI56/XI1/MM2_g
+ N_VSS_XI56/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI1/MM3 N_XI56/XI1/NET33_XI56/XI1/MM3_d N_WL<108>_XI56/XI1/MM3_g
+ N_BLN<14>_XI56/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI1/MM0 N_XI56/XI1/NET34_XI56/XI1/MM0_d N_WL<108>_XI56/XI1/MM0_g
+ N_BL<14>_XI56/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI1/MM1 N_XI56/XI1/NET33_XI56/XI1/MM1_d N_XI56/XI1/NET34_XI56/XI1/MM1_g
+ N_VSS_XI56/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI1/MM9 N_XI56/XI1/NET36_XI56/XI1/MM9_d N_WL<109>_XI56/XI1/MM9_g
+ N_BL<14>_XI56/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI1/MM6 N_XI56/XI1/NET35_XI56/XI1/MM6_d N_XI56/XI1/NET36_XI56/XI1/MM6_g
+ N_VSS_XI56/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI1/MM7 N_XI56/XI1/NET36_XI56/XI1/MM7_d N_XI56/XI1/NET35_XI56/XI1/MM7_g
+ N_VSS_XI56/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI1/MM8 N_XI56/XI1/NET35_XI56/XI1/MM8_d N_WL<109>_XI56/XI1/MM8_g
+ N_BLN<14>_XI56/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI1/MM5 N_XI56/XI1/NET34_XI56/XI1/MM5_d N_XI56/XI1/NET33_XI56/XI1/MM5_g
+ N_VDD_XI56/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI1/MM4 N_XI56/XI1/NET33_XI56/XI1/MM4_d N_XI56/XI1/NET34_XI56/XI1/MM4_g
+ N_VDD_XI56/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI1/MM10 N_XI56/XI1/NET35_XI56/XI1/MM10_d N_XI56/XI1/NET36_XI56/XI1/MM10_g
+ N_VDD_XI56/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI1/MM11 N_XI56/XI1/NET36_XI56/XI1/MM11_d N_XI56/XI1/NET35_XI56/XI1/MM11_g
+ N_VDD_XI56/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI2/MM2 N_XI56/XI2/NET34_XI56/XI2/MM2_d N_XI56/XI2/NET33_XI56/XI2/MM2_g
+ N_VSS_XI56/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI2/MM3 N_XI56/XI2/NET33_XI56/XI2/MM3_d N_WL<108>_XI56/XI2/MM3_g
+ N_BLN<13>_XI56/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI2/MM0 N_XI56/XI2/NET34_XI56/XI2/MM0_d N_WL<108>_XI56/XI2/MM0_g
+ N_BL<13>_XI56/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI2/MM1 N_XI56/XI2/NET33_XI56/XI2/MM1_d N_XI56/XI2/NET34_XI56/XI2/MM1_g
+ N_VSS_XI56/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI2/MM9 N_XI56/XI2/NET36_XI56/XI2/MM9_d N_WL<109>_XI56/XI2/MM9_g
+ N_BL<13>_XI56/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI2/MM6 N_XI56/XI2/NET35_XI56/XI2/MM6_d N_XI56/XI2/NET36_XI56/XI2/MM6_g
+ N_VSS_XI56/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI2/MM7 N_XI56/XI2/NET36_XI56/XI2/MM7_d N_XI56/XI2/NET35_XI56/XI2/MM7_g
+ N_VSS_XI56/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI2/MM8 N_XI56/XI2/NET35_XI56/XI2/MM8_d N_WL<109>_XI56/XI2/MM8_g
+ N_BLN<13>_XI56/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI2/MM5 N_XI56/XI2/NET34_XI56/XI2/MM5_d N_XI56/XI2/NET33_XI56/XI2/MM5_g
+ N_VDD_XI56/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI2/MM4 N_XI56/XI2/NET33_XI56/XI2/MM4_d N_XI56/XI2/NET34_XI56/XI2/MM4_g
+ N_VDD_XI56/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI2/MM10 N_XI56/XI2/NET35_XI56/XI2/MM10_d N_XI56/XI2/NET36_XI56/XI2/MM10_g
+ N_VDD_XI56/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI2/MM11 N_XI56/XI2/NET36_XI56/XI2/MM11_d N_XI56/XI2/NET35_XI56/XI2/MM11_g
+ N_VDD_XI56/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI3/MM2 N_XI56/XI3/NET34_XI56/XI3/MM2_d N_XI56/XI3/NET33_XI56/XI3/MM2_g
+ N_VSS_XI56/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI3/MM3 N_XI56/XI3/NET33_XI56/XI3/MM3_d N_WL<108>_XI56/XI3/MM3_g
+ N_BLN<12>_XI56/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI3/MM0 N_XI56/XI3/NET34_XI56/XI3/MM0_d N_WL<108>_XI56/XI3/MM0_g
+ N_BL<12>_XI56/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI3/MM1 N_XI56/XI3/NET33_XI56/XI3/MM1_d N_XI56/XI3/NET34_XI56/XI3/MM1_g
+ N_VSS_XI56/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI3/MM9 N_XI56/XI3/NET36_XI56/XI3/MM9_d N_WL<109>_XI56/XI3/MM9_g
+ N_BL<12>_XI56/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI3/MM6 N_XI56/XI3/NET35_XI56/XI3/MM6_d N_XI56/XI3/NET36_XI56/XI3/MM6_g
+ N_VSS_XI56/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI3/MM7 N_XI56/XI3/NET36_XI56/XI3/MM7_d N_XI56/XI3/NET35_XI56/XI3/MM7_g
+ N_VSS_XI56/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI3/MM8 N_XI56/XI3/NET35_XI56/XI3/MM8_d N_WL<109>_XI56/XI3/MM8_g
+ N_BLN<12>_XI56/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI3/MM5 N_XI56/XI3/NET34_XI56/XI3/MM5_d N_XI56/XI3/NET33_XI56/XI3/MM5_g
+ N_VDD_XI56/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI3/MM4 N_XI56/XI3/NET33_XI56/XI3/MM4_d N_XI56/XI3/NET34_XI56/XI3/MM4_g
+ N_VDD_XI56/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI3/MM10 N_XI56/XI3/NET35_XI56/XI3/MM10_d N_XI56/XI3/NET36_XI56/XI3/MM10_g
+ N_VDD_XI56/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI3/MM11 N_XI56/XI3/NET36_XI56/XI3/MM11_d N_XI56/XI3/NET35_XI56/XI3/MM11_g
+ N_VDD_XI56/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI4/MM2 N_XI56/XI4/NET34_XI56/XI4/MM2_d N_XI56/XI4/NET33_XI56/XI4/MM2_g
+ N_VSS_XI56/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI4/MM3 N_XI56/XI4/NET33_XI56/XI4/MM3_d N_WL<108>_XI56/XI4/MM3_g
+ N_BLN<11>_XI56/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI4/MM0 N_XI56/XI4/NET34_XI56/XI4/MM0_d N_WL<108>_XI56/XI4/MM0_g
+ N_BL<11>_XI56/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI4/MM1 N_XI56/XI4/NET33_XI56/XI4/MM1_d N_XI56/XI4/NET34_XI56/XI4/MM1_g
+ N_VSS_XI56/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI4/MM9 N_XI56/XI4/NET36_XI56/XI4/MM9_d N_WL<109>_XI56/XI4/MM9_g
+ N_BL<11>_XI56/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI4/MM6 N_XI56/XI4/NET35_XI56/XI4/MM6_d N_XI56/XI4/NET36_XI56/XI4/MM6_g
+ N_VSS_XI56/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI4/MM7 N_XI56/XI4/NET36_XI56/XI4/MM7_d N_XI56/XI4/NET35_XI56/XI4/MM7_g
+ N_VSS_XI56/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI4/MM8 N_XI56/XI4/NET35_XI56/XI4/MM8_d N_WL<109>_XI56/XI4/MM8_g
+ N_BLN<11>_XI56/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI4/MM5 N_XI56/XI4/NET34_XI56/XI4/MM5_d N_XI56/XI4/NET33_XI56/XI4/MM5_g
+ N_VDD_XI56/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI4/MM4 N_XI56/XI4/NET33_XI56/XI4/MM4_d N_XI56/XI4/NET34_XI56/XI4/MM4_g
+ N_VDD_XI56/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI4/MM10 N_XI56/XI4/NET35_XI56/XI4/MM10_d N_XI56/XI4/NET36_XI56/XI4/MM10_g
+ N_VDD_XI56/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI4/MM11 N_XI56/XI4/NET36_XI56/XI4/MM11_d N_XI56/XI4/NET35_XI56/XI4/MM11_g
+ N_VDD_XI56/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI5/MM2 N_XI56/XI5/NET34_XI56/XI5/MM2_d N_XI56/XI5/NET33_XI56/XI5/MM2_g
+ N_VSS_XI56/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI5/MM3 N_XI56/XI5/NET33_XI56/XI5/MM3_d N_WL<108>_XI56/XI5/MM3_g
+ N_BLN<10>_XI56/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI5/MM0 N_XI56/XI5/NET34_XI56/XI5/MM0_d N_WL<108>_XI56/XI5/MM0_g
+ N_BL<10>_XI56/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI5/MM1 N_XI56/XI5/NET33_XI56/XI5/MM1_d N_XI56/XI5/NET34_XI56/XI5/MM1_g
+ N_VSS_XI56/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI5/MM9 N_XI56/XI5/NET36_XI56/XI5/MM9_d N_WL<109>_XI56/XI5/MM9_g
+ N_BL<10>_XI56/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI5/MM6 N_XI56/XI5/NET35_XI56/XI5/MM6_d N_XI56/XI5/NET36_XI56/XI5/MM6_g
+ N_VSS_XI56/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI5/MM7 N_XI56/XI5/NET36_XI56/XI5/MM7_d N_XI56/XI5/NET35_XI56/XI5/MM7_g
+ N_VSS_XI56/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI5/MM8 N_XI56/XI5/NET35_XI56/XI5/MM8_d N_WL<109>_XI56/XI5/MM8_g
+ N_BLN<10>_XI56/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI5/MM5 N_XI56/XI5/NET34_XI56/XI5/MM5_d N_XI56/XI5/NET33_XI56/XI5/MM5_g
+ N_VDD_XI56/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI5/MM4 N_XI56/XI5/NET33_XI56/XI5/MM4_d N_XI56/XI5/NET34_XI56/XI5/MM4_g
+ N_VDD_XI56/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI5/MM10 N_XI56/XI5/NET35_XI56/XI5/MM10_d N_XI56/XI5/NET36_XI56/XI5/MM10_g
+ N_VDD_XI56/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI5/MM11 N_XI56/XI5/NET36_XI56/XI5/MM11_d N_XI56/XI5/NET35_XI56/XI5/MM11_g
+ N_VDD_XI56/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI6/MM2 N_XI56/XI6/NET34_XI56/XI6/MM2_d N_XI56/XI6/NET33_XI56/XI6/MM2_g
+ N_VSS_XI56/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM3 N_XI56/XI6/NET33_XI56/XI6/MM3_d N_WL<108>_XI56/XI6/MM3_g
+ N_BLN<9>_XI56/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM0 N_XI56/XI6/NET34_XI56/XI6/MM0_d N_WL<108>_XI56/XI6/MM0_g
+ N_BL<9>_XI56/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM1 N_XI56/XI6/NET33_XI56/XI6/MM1_d N_XI56/XI6/NET34_XI56/XI6/MM1_g
+ N_VSS_XI56/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM9 N_XI56/XI6/NET36_XI56/XI6/MM9_d N_WL<109>_XI56/XI6/MM9_g
+ N_BL<9>_XI56/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM6 N_XI56/XI6/NET35_XI56/XI6/MM6_d N_XI56/XI6/NET36_XI56/XI6/MM6_g
+ N_VSS_XI56/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM7 N_XI56/XI6/NET36_XI56/XI6/MM7_d N_XI56/XI6/NET35_XI56/XI6/MM7_g
+ N_VSS_XI56/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM8 N_XI56/XI6/NET35_XI56/XI6/MM8_d N_WL<109>_XI56/XI6/MM8_g
+ N_BLN<9>_XI56/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI6/MM5 N_XI56/XI6/NET34_XI56/XI6/MM5_d N_XI56/XI6/NET33_XI56/XI6/MM5_g
+ N_VDD_XI56/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI6/MM4 N_XI56/XI6/NET33_XI56/XI6/MM4_d N_XI56/XI6/NET34_XI56/XI6/MM4_g
+ N_VDD_XI56/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI6/MM10 N_XI56/XI6/NET35_XI56/XI6/MM10_d N_XI56/XI6/NET36_XI56/XI6/MM10_g
+ N_VDD_XI56/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI6/MM11 N_XI56/XI6/NET36_XI56/XI6/MM11_d N_XI56/XI6/NET35_XI56/XI6/MM11_g
+ N_VDD_XI56/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI7/MM2 N_XI56/XI7/NET34_XI56/XI7/MM2_d N_XI56/XI7/NET33_XI56/XI7/MM2_g
+ N_VSS_XI56/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM3 N_XI56/XI7/NET33_XI56/XI7/MM3_d N_WL<108>_XI56/XI7/MM3_g
+ N_BLN<8>_XI56/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM0 N_XI56/XI7/NET34_XI56/XI7/MM0_d N_WL<108>_XI56/XI7/MM0_g
+ N_BL<8>_XI56/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM1 N_XI56/XI7/NET33_XI56/XI7/MM1_d N_XI56/XI7/NET34_XI56/XI7/MM1_g
+ N_VSS_XI56/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM9 N_XI56/XI7/NET36_XI56/XI7/MM9_d N_WL<109>_XI56/XI7/MM9_g
+ N_BL<8>_XI56/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM6 N_XI56/XI7/NET35_XI56/XI7/MM6_d N_XI56/XI7/NET36_XI56/XI7/MM6_g
+ N_VSS_XI56/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM7 N_XI56/XI7/NET36_XI56/XI7/MM7_d N_XI56/XI7/NET35_XI56/XI7/MM7_g
+ N_VSS_XI56/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM8 N_XI56/XI7/NET35_XI56/XI7/MM8_d N_WL<109>_XI56/XI7/MM8_g
+ N_BLN<8>_XI56/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI7/MM5 N_XI56/XI7/NET34_XI56/XI7/MM5_d N_XI56/XI7/NET33_XI56/XI7/MM5_g
+ N_VDD_XI56/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI7/MM4 N_XI56/XI7/NET33_XI56/XI7/MM4_d N_XI56/XI7/NET34_XI56/XI7/MM4_g
+ N_VDD_XI56/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI7/MM10 N_XI56/XI7/NET35_XI56/XI7/MM10_d N_XI56/XI7/NET36_XI56/XI7/MM10_g
+ N_VDD_XI56/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI7/MM11 N_XI56/XI7/NET36_XI56/XI7/MM11_d N_XI56/XI7/NET35_XI56/XI7/MM11_g
+ N_VDD_XI56/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI8/MM2 N_XI56/XI8/NET34_XI56/XI8/MM2_d N_XI56/XI8/NET33_XI56/XI8/MM2_g
+ N_VSS_XI56/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM3 N_XI56/XI8/NET33_XI56/XI8/MM3_d N_WL<108>_XI56/XI8/MM3_g
+ N_BLN<7>_XI56/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM0 N_XI56/XI8/NET34_XI56/XI8/MM0_d N_WL<108>_XI56/XI8/MM0_g
+ N_BL<7>_XI56/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM1 N_XI56/XI8/NET33_XI56/XI8/MM1_d N_XI56/XI8/NET34_XI56/XI8/MM1_g
+ N_VSS_XI56/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM9 N_XI56/XI8/NET36_XI56/XI8/MM9_d N_WL<109>_XI56/XI8/MM9_g
+ N_BL<7>_XI56/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM6 N_XI56/XI8/NET35_XI56/XI8/MM6_d N_XI56/XI8/NET36_XI56/XI8/MM6_g
+ N_VSS_XI56/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM7 N_XI56/XI8/NET36_XI56/XI8/MM7_d N_XI56/XI8/NET35_XI56/XI8/MM7_g
+ N_VSS_XI56/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM8 N_XI56/XI8/NET35_XI56/XI8/MM8_d N_WL<109>_XI56/XI8/MM8_g
+ N_BLN<7>_XI56/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI8/MM5 N_XI56/XI8/NET34_XI56/XI8/MM5_d N_XI56/XI8/NET33_XI56/XI8/MM5_g
+ N_VDD_XI56/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI8/MM4 N_XI56/XI8/NET33_XI56/XI8/MM4_d N_XI56/XI8/NET34_XI56/XI8/MM4_g
+ N_VDD_XI56/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI8/MM10 N_XI56/XI8/NET35_XI56/XI8/MM10_d N_XI56/XI8/NET36_XI56/XI8/MM10_g
+ N_VDD_XI56/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI8/MM11 N_XI56/XI8/NET36_XI56/XI8/MM11_d N_XI56/XI8/NET35_XI56/XI8/MM11_g
+ N_VDD_XI56/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI9/MM2 N_XI56/XI9/NET34_XI56/XI9/MM2_d N_XI56/XI9/NET33_XI56/XI9/MM2_g
+ N_VSS_XI56/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM3 N_XI56/XI9/NET33_XI56/XI9/MM3_d N_WL<108>_XI56/XI9/MM3_g
+ N_BLN<6>_XI56/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM0 N_XI56/XI9/NET34_XI56/XI9/MM0_d N_WL<108>_XI56/XI9/MM0_g
+ N_BL<6>_XI56/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM1 N_XI56/XI9/NET33_XI56/XI9/MM1_d N_XI56/XI9/NET34_XI56/XI9/MM1_g
+ N_VSS_XI56/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM9 N_XI56/XI9/NET36_XI56/XI9/MM9_d N_WL<109>_XI56/XI9/MM9_g
+ N_BL<6>_XI56/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM6 N_XI56/XI9/NET35_XI56/XI9/MM6_d N_XI56/XI9/NET36_XI56/XI9/MM6_g
+ N_VSS_XI56/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM7 N_XI56/XI9/NET36_XI56/XI9/MM7_d N_XI56/XI9/NET35_XI56/XI9/MM7_g
+ N_VSS_XI56/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM8 N_XI56/XI9/NET35_XI56/XI9/MM8_d N_WL<109>_XI56/XI9/MM8_g
+ N_BLN<6>_XI56/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI9/MM5 N_XI56/XI9/NET34_XI56/XI9/MM5_d N_XI56/XI9/NET33_XI56/XI9/MM5_g
+ N_VDD_XI56/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI9/MM4 N_XI56/XI9/NET33_XI56/XI9/MM4_d N_XI56/XI9/NET34_XI56/XI9/MM4_g
+ N_VDD_XI56/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI9/MM10 N_XI56/XI9/NET35_XI56/XI9/MM10_d N_XI56/XI9/NET36_XI56/XI9/MM10_g
+ N_VDD_XI56/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI9/MM11 N_XI56/XI9/NET36_XI56/XI9/MM11_d N_XI56/XI9/NET35_XI56/XI9/MM11_g
+ N_VDD_XI56/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI10/MM2 N_XI56/XI10/NET34_XI56/XI10/MM2_d
+ N_XI56/XI10/NET33_XI56/XI10/MM2_g N_VSS_XI56/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI10/MM3 N_XI56/XI10/NET33_XI56/XI10/MM3_d N_WL<108>_XI56/XI10/MM3_g
+ N_BLN<5>_XI56/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI10/MM0 N_XI56/XI10/NET34_XI56/XI10/MM0_d N_WL<108>_XI56/XI10/MM0_g
+ N_BL<5>_XI56/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI10/MM1 N_XI56/XI10/NET33_XI56/XI10/MM1_d
+ N_XI56/XI10/NET34_XI56/XI10/MM1_g N_VSS_XI56/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI10/MM9 N_XI56/XI10/NET36_XI56/XI10/MM9_d N_WL<109>_XI56/XI10/MM9_g
+ N_BL<5>_XI56/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI10/MM6 N_XI56/XI10/NET35_XI56/XI10/MM6_d
+ N_XI56/XI10/NET36_XI56/XI10/MM6_g N_VSS_XI56/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI10/MM7 N_XI56/XI10/NET36_XI56/XI10/MM7_d
+ N_XI56/XI10/NET35_XI56/XI10/MM7_g N_VSS_XI56/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI10/MM8 N_XI56/XI10/NET35_XI56/XI10/MM8_d N_WL<109>_XI56/XI10/MM8_g
+ N_BLN<5>_XI56/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI10/MM5 N_XI56/XI10/NET34_XI56/XI10/MM5_d
+ N_XI56/XI10/NET33_XI56/XI10/MM5_g N_VDD_XI56/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI10/MM4 N_XI56/XI10/NET33_XI56/XI10/MM4_d
+ N_XI56/XI10/NET34_XI56/XI10/MM4_g N_VDD_XI56/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI10/MM10 N_XI56/XI10/NET35_XI56/XI10/MM10_d
+ N_XI56/XI10/NET36_XI56/XI10/MM10_g N_VDD_XI56/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI10/MM11 N_XI56/XI10/NET36_XI56/XI10/MM11_d
+ N_XI56/XI10/NET35_XI56/XI10/MM11_g N_VDD_XI56/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI11/MM2 N_XI56/XI11/NET34_XI56/XI11/MM2_d
+ N_XI56/XI11/NET33_XI56/XI11/MM2_g N_VSS_XI56/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI11/MM3 N_XI56/XI11/NET33_XI56/XI11/MM3_d N_WL<108>_XI56/XI11/MM3_g
+ N_BLN<4>_XI56/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI11/MM0 N_XI56/XI11/NET34_XI56/XI11/MM0_d N_WL<108>_XI56/XI11/MM0_g
+ N_BL<4>_XI56/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI11/MM1 N_XI56/XI11/NET33_XI56/XI11/MM1_d
+ N_XI56/XI11/NET34_XI56/XI11/MM1_g N_VSS_XI56/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI11/MM9 N_XI56/XI11/NET36_XI56/XI11/MM9_d N_WL<109>_XI56/XI11/MM9_g
+ N_BL<4>_XI56/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI11/MM6 N_XI56/XI11/NET35_XI56/XI11/MM6_d
+ N_XI56/XI11/NET36_XI56/XI11/MM6_g N_VSS_XI56/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI11/MM7 N_XI56/XI11/NET36_XI56/XI11/MM7_d
+ N_XI56/XI11/NET35_XI56/XI11/MM7_g N_VSS_XI56/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI11/MM8 N_XI56/XI11/NET35_XI56/XI11/MM8_d N_WL<109>_XI56/XI11/MM8_g
+ N_BLN<4>_XI56/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI11/MM5 N_XI56/XI11/NET34_XI56/XI11/MM5_d
+ N_XI56/XI11/NET33_XI56/XI11/MM5_g N_VDD_XI56/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI11/MM4 N_XI56/XI11/NET33_XI56/XI11/MM4_d
+ N_XI56/XI11/NET34_XI56/XI11/MM4_g N_VDD_XI56/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI11/MM10 N_XI56/XI11/NET35_XI56/XI11/MM10_d
+ N_XI56/XI11/NET36_XI56/XI11/MM10_g N_VDD_XI56/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI11/MM11 N_XI56/XI11/NET36_XI56/XI11/MM11_d
+ N_XI56/XI11/NET35_XI56/XI11/MM11_g N_VDD_XI56/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI12/MM2 N_XI56/XI12/NET34_XI56/XI12/MM2_d
+ N_XI56/XI12/NET33_XI56/XI12/MM2_g N_VSS_XI56/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI12/MM3 N_XI56/XI12/NET33_XI56/XI12/MM3_d N_WL<108>_XI56/XI12/MM3_g
+ N_BLN<3>_XI56/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI12/MM0 N_XI56/XI12/NET34_XI56/XI12/MM0_d N_WL<108>_XI56/XI12/MM0_g
+ N_BL<3>_XI56/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI12/MM1 N_XI56/XI12/NET33_XI56/XI12/MM1_d
+ N_XI56/XI12/NET34_XI56/XI12/MM1_g N_VSS_XI56/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI12/MM9 N_XI56/XI12/NET36_XI56/XI12/MM9_d N_WL<109>_XI56/XI12/MM9_g
+ N_BL<3>_XI56/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI12/MM6 N_XI56/XI12/NET35_XI56/XI12/MM6_d
+ N_XI56/XI12/NET36_XI56/XI12/MM6_g N_VSS_XI56/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI12/MM7 N_XI56/XI12/NET36_XI56/XI12/MM7_d
+ N_XI56/XI12/NET35_XI56/XI12/MM7_g N_VSS_XI56/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI12/MM8 N_XI56/XI12/NET35_XI56/XI12/MM8_d N_WL<109>_XI56/XI12/MM8_g
+ N_BLN<3>_XI56/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI12/MM5 N_XI56/XI12/NET34_XI56/XI12/MM5_d
+ N_XI56/XI12/NET33_XI56/XI12/MM5_g N_VDD_XI56/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI12/MM4 N_XI56/XI12/NET33_XI56/XI12/MM4_d
+ N_XI56/XI12/NET34_XI56/XI12/MM4_g N_VDD_XI56/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI12/MM10 N_XI56/XI12/NET35_XI56/XI12/MM10_d
+ N_XI56/XI12/NET36_XI56/XI12/MM10_g N_VDD_XI56/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI12/MM11 N_XI56/XI12/NET36_XI56/XI12/MM11_d
+ N_XI56/XI12/NET35_XI56/XI12/MM11_g N_VDD_XI56/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI13/MM2 N_XI56/XI13/NET34_XI56/XI13/MM2_d
+ N_XI56/XI13/NET33_XI56/XI13/MM2_g N_VSS_XI56/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI13/MM3 N_XI56/XI13/NET33_XI56/XI13/MM3_d N_WL<108>_XI56/XI13/MM3_g
+ N_BLN<2>_XI56/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI13/MM0 N_XI56/XI13/NET34_XI56/XI13/MM0_d N_WL<108>_XI56/XI13/MM0_g
+ N_BL<2>_XI56/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI13/MM1 N_XI56/XI13/NET33_XI56/XI13/MM1_d
+ N_XI56/XI13/NET34_XI56/XI13/MM1_g N_VSS_XI56/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI13/MM9 N_XI56/XI13/NET36_XI56/XI13/MM9_d N_WL<109>_XI56/XI13/MM9_g
+ N_BL<2>_XI56/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI13/MM6 N_XI56/XI13/NET35_XI56/XI13/MM6_d
+ N_XI56/XI13/NET36_XI56/XI13/MM6_g N_VSS_XI56/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI13/MM7 N_XI56/XI13/NET36_XI56/XI13/MM7_d
+ N_XI56/XI13/NET35_XI56/XI13/MM7_g N_VSS_XI56/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI13/MM8 N_XI56/XI13/NET35_XI56/XI13/MM8_d N_WL<109>_XI56/XI13/MM8_g
+ N_BLN<2>_XI56/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI13/MM5 N_XI56/XI13/NET34_XI56/XI13/MM5_d
+ N_XI56/XI13/NET33_XI56/XI13/MM5_g N_VDD_XI56/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI13/MM4 N_XI56/XI13/NET33_XI56/XI13/MM4_d
+ N_XI56/XI13/NET34_XI56/XI13/MM4_g N_VDD_XI56/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI13/MM10 N_XI56/XI13/NET35_XI56/XI13/MM10_d
+ N_XI56/XI13/NET36_XI56/XI13/MM10_g N_VDD_XI56/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI13/MM11 N_XI56/XI13/NET36_XI56/XI13/MM11_d
+ N_XI56/XI13/NET35_XI56/XI13/MM11_g N_VDD_XI56/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI14/MM2 N_XI56/XI14/NET34_XI56/XI14/MM2_d
+ N_XI56/XI14/NET33_XI56/XI14/MM2_g N_VSS_XI56/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI14/MM3 N_XI56/XI14/NET33_XI56/XI14/MM3_d N_WL<108>_XI56/XI14/MM3_g
+ N_BLN<1>_XI56/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI14/MM0 N_XI56/XI14/NET34_XI56/XI14/MM0_d N_WL<108>_XI56/XI14/MM0_g
+ N_BL<1>_XI56/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI14/MM1 N_XI56/XI14/NET33_XI56/XI14/MM1_d
+ N_XI56/XI14/NET34_XI56/XI14/MM1_g N_VSS_XI56/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI14/MM9 N_XI56/XI14/NET36_XI56/XI14/MM9_d N_WL<109>_XI56/XI14/MM9_g
+ N_BL<1>_XI56/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI14/MM6 N_XI56/XI14/NET35_XI56/XI14/MM6_d
+ N_XI56/XI14/NET36_XI56/XI14/MM6_g N_VSS_XI56/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI14/MM7 N_XI56/XI14/NET36_XI56/XI14/MM7_d
+ N_XI56/XI14/NET35_XI56/XI14/MM7_g N_VSS_XI56/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI14/MM8 N_XI56/XI14/NET35_XI56/XI14/MM8_d N_WL<109>_XI56/XI14/MM8_g
+ N_BLN<1>_XI56/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI14/MM5 N_XI56/XI14/NET34_XI56/XI14/MM5_d
+ N_XI56/XI14/NET33_XI56/XI14/MM5_g N_VDD_XI56/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI14/MM4 N_XI56/XI14/NET33_XI56/XI14/MM4_d
+ N_XI56/XI14/NET34_XI56/XI14/MM4_g N_VDD_XI56/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI14/MM10 N_XI56/XI14/NET35_XI56/XI14/MM10_d
+ N_XI56/XI14/NET36_XI56/XI14/MM10_g N_VDD_XI56/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI14/MM11 N_XI56/XI14/NET36_XI56/XI14/MM11_d
+ N_XI56/XI14/NET35_XI56/XI14/MM11_g N_VDD_XI56/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI15/MM2 N_XI56/XI15/NET34_XI56/XI15/MM2_d
+ N_XI56/XI15/NET33_XI56/XI15/MM2_g N_VSS_XI56/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI15/MM3 N_XI56/XI15/NET33_XI56/XI15/MM3_d N_WL<108>_XI56/XI15/MM3_g
+ N_BLN<0>_XI56/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI15/MM0 N_XI56/XI15/NET34_XI56/XI15/MM0_d N_WL<108>_XI56/XI15/MM0_g
+ N_BL<0>_XI56/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI15/MM1 N_XI56/XI15/NET33_XI56/XI15/MM1_d
+ N_XI56/XI15/NET34_XI56/XI15/MM1_g N_VSS_XI56/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI15/MM9 N_XI56/XI15/NET36_XI56/XI15/MM9_d N_WL<109>_XI56/XI15/MM9_g
+ N_BL<0>_XI56/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI15/MM6 N_XI56/XI15/NET35_XI56/XI15/MM6_d
+ N_XI56/XI15/NET36_XI56/XI15/MM6_g N_VSS_XI56/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI15/MM7 N_XI56/XI15/NET36_XI56/XI15/MM7_d
+ N_XI56/XI15/NET35_XI56/XI15/MM7_g N_VSS_XI56/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI56/XI15/MM8 N_XI56/XI15/NET35_XI56/XI15/MM8_d N_WL<109>_XI56/XI15/MM8_g
+ N_BLN<0>_XI56/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI56/XI15/MM5 N_XI56/XI15/NET34_XI56/XI15/MM5_d
+ N_XI56/XI15/NET33_XI56/XI15/MM5_g N_VDD_XI56/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI15/MM4 N_XI56/XI15/NET33_XI56/XI15/MM4_d
+ N_XI56/XI15/NET34_XI56/XI15/MM4_g N_VDD_XI56/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI15/MM10 N_XI56/XI15/NET35_XI56/XI15/MM10_d
+ N_XI56/XI15/NET36_XI56/XI15/MM10_g N_VDD_XI56/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI56/XI15/MM11 N_XI56/XI15/NET36_XI56/XI15/MM11_d
+ N_XI56/XI15/NET35_XI56/XI15/MM11_g N_VDD_XI56/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI0/MM2 N_XI57/XI0/NET34_XI57/XI0/MM2_d N_XI57/XI0/NET33_XI57/XI0/MM2_g
+ N_VSS_XI57/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI0/MM3 N_XI57/XI0/NET33_XI57/XI0/MM3_d N_WL<110>_XI57/XI0/MM3_g
+ N_BLN<15>_XI57/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI0/MM0 N_XI57/XI0/NET34_XI57/XI0/MM0_d N_WL<110>_XI57/XI0/MM0_g
+ N_BL<15>_XI57/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI0/MM1 N_XI57/XI0/NET33_XI57/XI0/MM1_d N_XI57/XI0/NET34_XI57/XI0/MM1_g
+ N_VSS_XI57/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI0/MM9 N_XI57/XI0/NET36_XI57/XI0/MM9_d N_WL<111>_XI57/XI0/MM9_g
+ N_BL<15>_XI57/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI0/MM6 N_XI57/XI0/NET35_XI57/XI0/MM6_d N_XI57/XI0/NET36_XI57/XI0/MM6_g
+ N_VSS_XI57/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI0/MM7 N_XI57/XI0/NET36_XI57/XI0/MM7_d N_XI57/XI0/NET35_XI57/XI0/MM7_g
+ N_VSS_XI57/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI0/MM8 N_XI57/XI0/NET35_XI57/XI0/MM8_d N_WL<111>_XI57/XI0/MM8_g
+ N_BLN<15>_XI57/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI0/MM5 N_XI57/XI0/NET34_XI57/XI0/MM5_d N_XI57/XI0/NET33_XI57/XI0/MM5_g
+ N_VDD_XI57/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI0/MM4 N_XI57/XI0/NET33_XI57/XI0/MM4_d N_XI57/XI0/NET34_XI57/XI0/MM4_g
+ N_VDD_XI57/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI0/MM10 N_XI57/XI0/NET35_XI57/XI0/MM10_d N_XI57/XI0/NET36_XI57/XI0/MM10_g
+ N_VDD_XI57/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI0/MM11 N_XI57/XI0/NET36_XI57/XI0/MM11_d N_XI57/XI0/NET35_XI57/XI0/MM11_g
+ N_VDD_XI57/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI1/MM2 N_XI57/XI1/NET34_XI57/XI1/MM2_d N_XI57/XI1/NET33_XI57/XI1/MM2_g
+ N_VSS_XI57/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI1/MM3 N_XI57/XI1/NET33_XI57/XI1/MM3_d N_WL<110>_XI57/XI1/MM3_g
+ N_BLN<14>_XI57/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI1/MM0 N_XI57/XI1/NET34_XI57/XI1/MM0_d N_WL<110>_XI57/XI1/MM0_g
+ N_BL<14>_XI57/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI1/MM1 N_XI57/XI1/NET33_XI57/XI1/MM1_d N_XI57/XI1/NET34_XI57/XI1/MM1_g
+ N_VSS_XI57/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI1/MM9 N_XI57/XI1/NET36_XI57/XI1/MM9_d N_WL<111>_XI57/XI1/MM9_g
+ N_BL<14>_XI57/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI1/MM6 N_XI57/XI1/NET35_XI57/XI1/MM6_d N_XI57/XI1/NET36_XI57/XI1/MM6_g
+ N_VSS_XI57/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI1/MM7 N_XI57/XI1/NET36_XI57/XI1/MM7_d N_XI57/XI1/NET35_XI57/XI1/MM7_g
+ N_VSS_XI57/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI1/MM8 N_XI57/XI1/NET35_XI57/XI1/MM8_d N_WL<111>_XI57/XI1/MM8_g
+ N_BLN<14>_XI57/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI1/MM5 N_XI57/XI1/NET34_XI57/XI1/MM5_d N_XI57/XI1/NET33_XI57/XI1/MM5_g
+ N_VDD_XI57/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI1/MM4 N_XI57/XI1/NET33_XI57/XI1/MM4_d N_XI57/XI1/NET34_XI57/XI1/MM4_g
+ N_VDD_XI57/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI1/MM10 N_XI57/XI1/NET35_XI57/XI1/MM10_d N_XI57/XI1/NET36_XI57/XI1/MM10_g
+ N_VDD_XI57/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI1/MM11 N_XI57/XI1/NET36_XI57/XI1/MM11_d N_XI57/XI1/NET35_XI57/XI1/MM11_g
+ N_VDD_XI57/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI2/MM2 N_XI57/XI2/NET34_XI57/XI2/MM2_d N_XI57/XI2/NET33_XI57/XI2/MM2_g
+ N_VSS_XI57/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI2/MM3 N_XI57/XI2/NET33_XI57/XI2/MM3_d N_WL<110>_XI57/XI2/MM3_g
+ N_BLN<13>_XI57/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI2/MM0 N_XI57/XI2/NET34_XI57/XI2/MM0_d N_WL<110>_XI57/XI2/MM0_g
+ N_BL<13>_XI57/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI2/MM1 N_XI57/XI2/NET33_XI57/XI2/MM1_d N_XI57/XI2/NET34_XI57/XI2/MM1_g
+ N_VSS_XI57/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI2/MM9 N_XI57/XI2/NET36_XI57/XI2/MM9_d N_WL<111>_XI57/XI2/MM9_g
+ N_BL<13>_XI57/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI2/MM6 N_XI57/XI2/NET35_XI57/XI2/MM6_d N_XI57/XI2/NET36_XI57/XI2/MM6_g
+ N_VSS_XI57/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI2/MM7 N_XI57/XI2/NET36_XI57/XI2/MM7_d N_XI57/XI2/NET35_XI57/XI2/MM7_g
+ N_VSS_XI57/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI2/MM8 N_XI57/XI2/NET35_XI57/XI2/MM8_d N_WL<111>_XI57/XI2/MM8_g
+ N_BLN<13>_XI57/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI2/MM5 N_XI57/XI2/NET34_XI57/XI2/MM5_d N_XI57/XI2/NET33_XI57/XI2/MM5_g
+ N_VDD_XI57/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI2/MM4 N_XI57/XI2/NET33_XI57/XI2/MM4_d N_XI57/XI2/NET34_XI57/XI2/MM4_g
+ N_VDD_XI57/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI2/MM10 N_XI57/XI2/NET35_XI57/XI2/MM10_d N_XI57/XI2/NET36_XI57/XI2/MM10_g
+ N_VDD_XI57/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI2/MM11 N_XI57/XI2/NET36_XI57/XI2/MM11_d N_XI57/XI2/NET35_XI57/XI2/MM11_g
+ N_VDD_XI57/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI3/MM2 N_XI57/XI3/NET34_XI57/XI3/MM2_d N_XI57/XI3/NET33_XI57/XI3/MM2_g
+ N_VSS_XI57/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI3/MM3 N_XI57/XI3/NET33_XI57/XI3/MM3_d N_WL<110>_XI57/XI3/MM3_g
+ N_BLN<12>_XI57/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI3/MM0 N_XI57/XI3/NET34_XI57/XI3/MM0_d N_WL<110>_XI57/XI3/MM0_g
+ N_BL<12>_XI57/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI3/MM1 N_XI57/XI3/NET33_XI57/XI3/MM1_d N_XI57/XI3/NET34_XI57/XI3/MM1_g
+ N_VSS_XI57/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI3/MM9 N_XI57/XI3/NET36_XI57/XI3/MM9_d N_WL<111>_XI57/XI3/MM9_g
+ N_BL<12>_XI57/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI3/MM6 N_XI57/XI3/NET35_XI57/XI3/MM6_d N_XI57/XI3/NET36_XI57/XI3/MM6_g
+ N_VSS_XI57/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI3/MM7 N_XI57/XI3/NET36_XI57/XI3/MM7_d N_XI57/XI3/NET35_XI57/XI3/MM7_g
+ N_VSS_XI57/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI3/MM8 N_XI57/XI3/NET35_XI57/XI3/MM8_d N_WL<111>_XI57/XI3/MM8_g
+ N_BLN<12>_XI57/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI3/MM5 N_XI57/XI3/NET34_XI57/XI3/MM5_d N_XI57/XI3/NET33_XI57/XI3/MM5_g
+ N_VDD_XI57/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI3/MM4 N_XI57/XI3/NET33_XI57/XI3/MM4_d N_XI57/XI3/NET34_XI57/XI3/MM4_g
+ N_VDD_XI57/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI3/MM10 N_XI57/XI3/NET35_XI57/XI3/MM10_d N_XI57/XI3/NET36_XI57/XI3/MM10_g
+ N_VDD_XI57/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI3/MM11 N_XI57/XI3/NET36_XI57/XI3/MM11_d N_XI57/XI3/NET35_XI57/XI3/MM11_g
+ N_VDD_XI57/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI4/MM2 N_XI57/XI4/NET34_XI57/XI4/MM2_d N_XI57/XI4/NET33_XI57/XI4/MM2_g
+ N_VSS_XI57/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI4/MM3 N_XI57/XI4/NET33_XI57/XI4/MM3_d N_WL<110>_XI57/XI4/MM3_g
+ N_BLN<11>_XI57/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI4/MM0 N_XI57/XI4/NET34_XI57/XI4/MM0_d N_WL<110>_XI57/XI4/MM0_g
+ N_BL<11>_XI57/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI4/MM1 N_XI57/XI4/NET33_XI57/XI4/MM1_d N_XI57/XI4/NET34_XI57/XI4/MM1_g
+ N_VSS_XI57/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI4/MM9 N_XI57/XI4/NET36_XI57/XI4/MM9_d N_WL<111>_XI57/XI4/MM9_g
+ N_BL<11>_XI57/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI4/MM6 N_XI57/XI4/NET35_XI57/XI4/MM6_d N_XI57/XI4/NET36_XI57/XI4/MM6_g
+ N_VSS_XI57/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI4/MM7 N_XI57/XI4/NET36_XI57/XI4/MM7_d N_XI57/XI4/NET35_XI57/XI4/MM7_g
+ N_VSS_XI57/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI4/MM8 N_XI57/XI4/NET35_XI57/XI4/MM8_d N_WL<111>_XI57/XI4/MM8_g
+ N_BLN<11>_XI57/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI4/MM5 N_XI57/XI4/NET34_XI57/XI4/MM5_d N_XI57/XI4/NET33_XI57/XI4/MM5_g
+ N_VDD_XI57/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI4/MM4 N_XI57/XI4/NET33_XI57/XI4/MM4_d N_XI57/XI4/NET34_XI57/XI4/MM4_g
+ N_VDD_XI57/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI4/MM10 N_XI57/XI4/NET35_XI57/XI4/MM10_d N_XI57/XI4/NET36_XI57/XI4/MM10_g
+ N_VDD_XI57/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI4/MM11 N_XI57/XI4/NET36_XI57/XI4/MM11_d N_XI57/XI4/NET35_XI57/XI4/MM11_g
+ N_VDD_XI57/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI5/MM2 N_XI57/XI5/NET34_XI57/XI5/MM2_d N_XI57/XI5/NET33_XI57/XI5/MM2_g
+ N_VSS_XI57/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI5/MM3 N_XI57/XI5/NET33_XI57/XI5/MM3_d N_WL<110>_XI57/XI5/MM3_g
+ N_BLN<10>_XI57/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI5/MM0 N_XI57/XI5/NET34_XI57/XI5/MM0_d N_WL<110>_XI57/XI5/MM0_g
+ N_BL<10>_XI57/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI5/MM1 N_XI57/XI5/NET33_XI57/XI5/MM1_d N_XI57/XI5/NET34_XI57/XI5/MM1_g
+ N_VSS_XI57/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI5/MM9 N_XI57/XI5/NET36_XI57/XI5/MM9_d N_WL<111>_XI57/XI5/MM9_g
+ N_BL<10>_XI57/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI5/MM6 N_XI57/XI5/NET35_XI57/XI5/MM6_d N_XI57/XI5/NET36_XI57/XI5/MM6_g
+ N_VSS_XI57/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI5/MM7 N_XI57/XI5/NET36_XI57/XI5/MM7_d N_XI57/XI5/NET35_XI57/XI5/MM7_g
+ N_VSS_XI57/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI5/MM8 N_XI57/XI5/NET35_XI57/XI5/MM8_d N_WL<111>_XI57/XI5/MM8_g
+ N_BLN<10>_XI57/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI5/MM5 N_XI57/XI5/NET34_XI57/XI5/MM5_d N_XI57/XI5/NET33_XI57/XI5/MM5_g
+ N_VDD_XI57/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI5/MM4 N_XI57/XI5/NET33_XI57/XI5/MM4_d N_XI57/XI5/NET34_XI57/XI5/MM4_g
+ N_VDD_XI57/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI5/MM10 N_XI57/XI5/NET35_XI57/XI5/MM10_d N_XI57/XI5/NET36_XI57/XI5/MM10_g
+ N_VDD_XI57/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI5/MM11 N_XI57/XI5/NET36_XI57/XI5/MM11_d N_XI57/XI5/NET35_XI57/XI5/MM11_g
+ N_VDD_XI57/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI6/MM2 N_XI57/XI6/NET34_XI57/XI6/MM2_d N_XI57/XI6/NET33_XI57/XI6/MM2_g
+ N_VSS_XI57/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM3 N_XI57/XI6/NET33_XI57/XI6/MM3_d N_WL<110>_XI57/XI6/MM3_g
+ N_BLN<9>_XI57/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM0 N_XI57/XI6/NET34_XI57/XI6/MM0_d N_WL<110>_XI57/XI6/MM0_g
+ N_BL<9>_XI57/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM1 N_XI57/XI6/NET33_XI57/XI6/MM1_d N_XI57/XI6/NET34_XI57/XI6/MM1_g
+ N_VSS_XI57/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM9 N_XI57/XI6/NET36_XI57/XI6/MM9_d N_WL<111>_XI57/XI6/MM9_g
+ N_BL<9>_XI57/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM6 N_XI57/XI6/NET35_XI57/XI6/MM6_d N_XI57/XI6/NET36_XI57/XI6/MM6_g
+ N_VSS_XI57/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM7 N_XI57/XI6/NET36_XI57/XI6/MM7_d N_XI57/XI6/NET35_XI57/XI6/MM7_g
+ N_VSS_XI57/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM8 N_XI57/XI6/NET35_XI57/XI6/MM8_d N_WL<111>_XI57/XI6/MM8_g
+ N_BLN<9>_XI57/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI6/MM5 N_XI57/XI6/NET34_XI57/XI6/MM5_d N_XI57/XI6/NET33_XI57/XI6/MM5_g
+ N_VDD_XI57/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI6/MM4 N_XI57/XI6/NET33_XI57/XI6/MM4_d N_XI57/XI6/NET34_XI57/XI6/MM4_g
+ N_VDD_XI57/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI6/MM10 N_XI57/XI6/NET35_XI57/XI6/MM10_d N_XI57/XI6/NET36_XI57/XI6/MM10_g
+ N_VDD_XI57/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI6/MM11 N_XI57/XI6/NET36_XI57/XI6/MM11_d N_XI57/XI6/NET35_XI57/XI6/MM11_g
+ N_VDD_XI57/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI7/MM2 N_XI57/XI7/NET34_XI57/XI7/MM2_d N_XI57/XI7/NET33_XI57/XI7/MM2_g
+ N_VSS_XI57/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM3 N_XI57/XI7/NET33_XI57/XI7/MM3_d N_WL<110>_XI57/XI7/MM3_g
+ N_BLN<8>_XI57/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM0 N_XI57/XI7/NET34_XI57/XI7/MM0_d N_WL<110>_XI57/XI7/MM0_g
+ N_BL<8>_XI57/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM1 N_XI57/XI7/NET33_XI57/XI7/MM1_d N_XI57/XI7/NET34_XI57/XI7/MM1_g
+ N_VSS_XI57/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM9 N_XI57/XI7/NET36_XI57/XI7/MM9_d N_WL<111>_XI57/XI7/MM9_g
+ N_BL<8>_XI57/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM6 N_XI57/XI7/NET35_XI57/XI7/MM6_d N_XI57/XI7/NET36_XI57/XI7/MM6_g
+ N_VSS_XI57/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM7 N_XI57/XI7/NET36_XI57/XI7/MM7_d N_XI57/XI7/NET35_XI57/XI7/MM7_g
+ N_VSS_XI57/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM8 N_XI57/XI7/NET35_XI57/XI7/MM8_d N_WL<111>_XI57/XI7/MM8_g
+ N_BLN<8>_XI57/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI7/MM5 N_XI57/XI7/NET34_XI57/XI7/MM5_d N_XI57/XI7/NET33_XI57/XI7/MM5_g
+ N_VDD_XI57/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI7/MM4 N_XI57/XI7/NET33_XI57/XI7/MM4_d N_XI57/XI7/NET34_XI57/XI7/MM4_g
+ N_VDD_XI57/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI7/MM10 N_XI57/XI7/NET35_XI57/XI7/MM10_d N_XI57/XI7/NET36_XI57/XI7/MM10_g
+ N_VDD_XI57/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI7/MM11 N_XI57/XI7/NET36_XI57/XI7/MM11_d N_XI57/XI7/NET35_XI57/XI7/MM11_g
+ N_VDD_XI57/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI8/MM2 N_XI57/XI8/NET34_XI57/XI8/MM2_d N_XI57/XI8/NET33_XI57/XI8/MM2_g
+ N_VSS_XI57/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM3 N_XI57/XI8/NET33_XI57/XI8/MM3_d N_WL<110>_XI57/XI8/MM3_g
+ N_BLN<7>_XI57/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM0 N_XI57/XI8/NET34_XI57/XI8/MM0_d N_WL<110>_XI57/XI8/MM0_g
+ N_BL<7>_XI57/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM1 N_XI57/XI8/NET33_XI57/XI8/MM1_d N_XI57/XI8/NET34_XI57/XI8/MM1_g
+ N_VSS_XI57/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM9 N_XI57/XI8/NET36_XI57/XI8/MM9_d N_WL<111>_XI57/XI8/MM9_g
+ N_BL<7>_XI57/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM6 N_XI57/XI8/NET35_XI57/XI8/MM6_d N_XI57/XI8/NET36_XI57/XI8/MM6_g
+ N_VSS_XI57/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM7 N_XI57/XI8/NET36_XI57/XI8/MM7_d N_XI57/XI8/NET35_XI57/XI8/MM7_g
+ N_VSS_XI57/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM8 N_XI57/XI8/NET35_XI57/XI8/MM8_d N_WL<111>_XI57/XI8/MM8_g
+ N_BLN<7>_XI57/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI8/MM5 N_XI57/XI8/NET34_XI57/XI8/MM5_d N_XI57/XI8/NET33_XI57/XI8/MM5_g
+ N_VDD_XI57/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI8/MM4 N_XI57/XI8/NET33_XI57/XI8/MM4_d N_XI57/XI8/NET34_XI57/XI8/MM4_g
+ N_VDD_XI57/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI8/MM10 N_XI57/XI8/NET35_XI57/XI8/MM10_d N_XI57/XI8/NET36_XI57/XI8/MM10_g
+ N_VDD_XI57/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI8/MM11 N_XI57/XI8/NET36_XI57/XI8/MM11_d N_XI57/XI8/NET35_XI57/XI8/MM11_g
+ N_VDD_XI57/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI9/MM2 N_XI57/XI9/NET34_XI57/XI9/MM2_d N_XI57/XI9/NET33_XI57/XI9/MM2_g
+ N_VSS_XI57/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM3 N_XI57/XI9/NET33_XI57/XI9/MM3_d N_WL<110>_XI57/XI9/MM3_g
+ N_BLN<6>_XI57/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM0 N_XI57/XI9/NET34_XI57/XI9/MM0_d N_WL<110>_XI57/XI9/MM0_g
+ N_BL<6>_XI57/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM1 N_XI57/XI9/NET33_XI57/XI9/MM1_d N_XI57/XI9/NET34_XI57/XI9/MM1_g
+ N_VSS_XI57/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM9 N_XI57/XI9/NET36_XI57/XI9/MM9_d N_WL<111>_XI57/XI9/MM9_g
+ N_BL<6>_XI57/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM6 N_XI57/XI9/NET35_XI57/XI9/MM6_d N_XI57/XI9/NET36_XI57/XI9/MM6_g
+ N_VSS_XI57/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM7 N_XI57/XI9/NET36_XI57/XI9/MM7_d N_XI57/XI9/NET35_XI57/XI9/MM7_g
+ N_VSS_XI57/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM8 N_XI57/XI9/NET35_XI57/XI9/MM8_d N_WL<111>_XI57/XI9/MM8_g
+ N_BLN<6>_XI57/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI9/MM5 N_XI57/XI9/NET34_XI57/XI9/MM5_d N_XI57/XI9/NET33_XI57/XI9/MM5_g
+ N_VDD_XI57/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI9/MM4 N_XI57/XI9/NET33_XI57/XI9/MM4_d N_XI57/XI9/NET34_XI57/XI9/MM4_g
+ N_VDD_XI57/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI9/MM10 N_XI57/XI9/NET35_XI57/XI9/MM10_d N_XI57/XI9/NET36_XI57/XI9/MM10_g
+ N_VDD_XI57/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI9/MM11 N_XI57/XI9/NET36_XI57/XI9/MM11_d N_XI57/XI9/NET35_XI57/XI9/MM11_g
+ N_VDD_XI57/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI10/MM2 N_XI57/XI10/NET34_XI57/XI10/MM2_d
+ N_XI57/XI10/NET33_XI57/XI10/MM2_g N_VSS_XI57/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI10/MM3 N_XI57/XI10/NET33_XI57/XI10/MM3_d N_WL<110>_XI57/XI10/MM3_g
+ N_BLN<5>_XI57/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI10/MM0 N_XI57/XI10/NET34_XI57/XI10/MM0_d N_WL<110>_XI57/XI10/MM0_g
+ N_BL<5>_XI57/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI10/MM1 N_XI57/XI10/NET33_XI57/XI10/MM1_d
+ N_XI57/XI10/NET34_XI57/XI10/MM1_g N_VSS_XI57/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI10/MM9 N_XI57/XI10/NET36_XI57/XI10/MM9_d N_WL<111>_XI57/XI10/MM9_g
+ N_BL<5>_XI57/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI10/MM6 N_XI57/XI10/NET35_XI57/XI10/MM6_d
+ N_XI57/XI10/NET36_XI57/XI10/MM6_g N_VSS_XI57/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI10/MM7 N_XI57/XI10/NET36_XI57/XI10/MM7_d
+ N_XI57/XI10/NET35_XI57/XI10/MM7_g N_VSS_XI57/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI10/MM8 N_XI57/XI10/NET35_XI57/XI10/MM8_d N_WL<111>_XI57/XI10/MM8_g
+ N_BLN<5>_XI57/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI10/MM5 N_XI57/XI10/NET34_XI57/XI10/MM5_d
+ N_XI57/XI10/NET33_XI57/XI10/MM5_g N_VDD_XI57/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI10/MM4 N_XI57/XI10/NET33_XI57/XI10/MM4_d
+ N_XI57/XI10/NET34_XI57/XI10/MM4_g N_VDD_XI57/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI10/MM10 N_XI57/XI10/NET35_XI57/XI10/MM10_d
+ N_XI57/XI10/NET36_XI57/XI10/MM10_g N_VDD_XI57/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI10/MM11 N_XI57/XI10/NET36_XI57/XI10/MM11_d
+ N_XI57/XI10/NET35_XI57/XI10/MM11_g N_VDD_XI57/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI11/MM2 N_XI57/XI11/NET34_XI57/XI11/MM2_d
+ N_XI57/XI11/NET33_XI57/XI11/MM2_g N_VSS_XI57/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI11/MM3 N_XI57/XI11/NET33_XI57/XI11/MM3_d N_WL<110>_XI57/XI11/MM3_g
+ N_BLN<4>_XI57/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI11/MM0 N_XI57/XI11/NET34_XI57/XI11/MM0_d N_WL<110>_XI57/XI11/MM0_g
+ N_BL<4>_XI57/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI11/MM1 N_XI57/XI11/NET33_XI57/XI11/MM1_d
+ N_XI57/XI11/NET34_XI57/XI11/MM1_g N_VSS_XI57/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI11/MM9 N_XI57/XI11/NET36_XI57/XI11/MM9_d N_WL<111>_XI57/XI11/MM9_g
+ N_BL<4>_XI57/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI11/MM6 N_XI57/XI11/NET35_XI57/XI11/MM6_d
+ N_XI57/XI11/NET36_XI57/XI11/MM6_g N_VSS_XI57/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI11/MM7 N_XI57/XI11/NET36_XI57/XI11/MM7_d
+ N_XI57/XI11/NET35_XI57/XI11/MM7_g N_VSS_XI57/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI11/MM8 N_XI57/XI11/NET35_XI57/XI11/MM8_d N_WL<111>_XI57/XI11/MM8_g
+ N_BLN<4>_XI57/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI11/MM5 N_XI57/XI11/NET34_XI57/XI11/MM5_d
+ N_XI57/XI11/NET33_XI57/XI11/MM5_g N_VDD_XI57/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI11/MM4 N_XI57/XI11/NET33_XI57/XI11/MM4_d
+ N_XI57/XI11/NET34_XI57/XI11/MM4_g N_VDD_XI57/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI11/MM10 N_XI57/XI11/NET35_XI57/XI11/MM10_d
+ N_XI57/XI11/NET36_XI57/XI11/MM10_g N_VDD_XI57/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI11/MM11 N_XI57/XI11/NET36_XI57/XI11/MM11_d
+ N_XI57/XI11/NET35_XI57/XI11/MM11_g N_VDD_XI57/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI12/MM2 N_XI57/XI12/NET34_XI57/XI12/MM2_d
+ N_XI57/XI12/NET33_XI57/XI12/MM2_g N_VSS_XI57/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI12/MM3 N_XI57/XI12/NET33_XI57/XI12/MM3_d N_WL<110>_XI57/XI12/MM3_g
+ N_BLN<3>_XI57/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI12/MM0 N_XI57/XI12/NET34_XI57/XI12/MM0_d N_WL<110>_XI57/XI12/MM0_g
+ N_BL<3>_XI57/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI12/MM1 N_XI57/XI12/NET33_XI57/XI12/MM1_d
+ N_XI57/XI12/NET34_XI57/XI12/MM1_g N_VSS_XI57/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI12/MM9 N_XI57/XI12/NET36_XI57/XI12/MM9_d N_WL<111>_XI57/XI12/MM9_g
+ N_BL<3>_XI57/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI12/MM6 N_XI57/XI12/NET35_XI57/XI12/MM6_d
+ N_XI57/XI12/NET36_XI57/XI12/MM6_g N_VSS_XI57/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI12/MM7 N_XI57/XI12/NET36_XI57/XI12/MM7_d
+ N_XI57/XI12/NET35_XI57/XI12/MM7_g N_VSS_XI57/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI12/MM8 N_XI57/XI12/NET35_XI57/XI12/MM8_d N_WL<111>_XI57/XI12/MM8_g
+ N_BLN<3>_XI57/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI12/MM5 N_XI57/XI12/NET34_XI57/XI12/MM5_d
+ N_XI57/XI12/NET33_XI57/XI12/MM5_g N_VDD_XI57/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI12/MM4 N_XI57/XI12/NET33_XI57/XI12/MM4_d
+ N_XI57/XI12/NET34_XI57/XI12/MM4_g N_VDD_XI57/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI12/MM10 N_XI57/XI12/NET35_XI57/XI12/MM10_d
+ N_XI57/XI12/NET36_XI57/XI12/MM10_g N_VDD_XI57/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI12/MM11 N_XI57/XI12/NET36_XI57/XI12/MM11_d
+ N_XI57/XI12/NET35_XI57/XI12/MM11_g N_VDD_XI57/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI13/MM2 N_XI57/XI13/NET34_XI57/XI13/MM2_d
+ N_XI57/XI13/NET33_XI57/XI13/MM2_g N_VSS_XI57/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI13/MM3 N_XI57/XI13/NET33_XI57/XI13/MM3_d N_WL<110>_XI57/XI13/MM3_g
+ N_BLN<2>_XI57/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI13/MM0 N_XI57/XI13/NET34_XI57/XI13/MM0_d N_WL<110>_XI57/XI13/MM0_g
+ N_BL<2>_XI57/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI13/MM1 N_XI57/XI13/NET33_XI57/XI13/MM1_d
+ N_XI57/XI13/NET34_XI57/XI13/MM1_g N_VSS_XI57/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI13/MM9 N_XI57/XI13/NET36_XI57/XI13/MM9_d N_WL<111>_XI57/XI13/MM9_g
+ N_BL<2>_XI57/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI13/MM6 N_XI57/XI13/NET35_XI57/XI13/MM6_d
+ N_XI57/XI13/NET36_XI57/XI13/MM6_g N_VSS_XI57/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI13/MM7 N_XI57/XI13/NET36_XI57/XI13/MM7_d
+ N_XI57/XI13/NET35_XI57/XI13/MM7_g N_VSS_XI57/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI13/MM8 N_XI57/XI13/NET35_XI57/XI13/MM8_d N_WL<111>_XI57/XI13/MM8_g
+ N_BLN<2>_XI57/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI13/MM5 N_XI57/XI13/NET34_XI57/XI13/MM5_d
+ N_XI57/XI13/NET33_XI57/XI13/MM5_g N_VDD_XI57/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI13/MM4 N_XI57/XI13/NET33_XI57/XI13/MM4_d
+ N_XI57/XI13/NET34_XI57/XI13/MM4_g N_VDD_XI57/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI13/MM10 N_XI57/XI13/NET35_XI57/XI13/MM10_d
+ N_XI57/XI13/NET36_XI57/XI13/MM10_g N_VDD_XI57/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI13/MM11 N_XI57/XI13/NET36_XI57/XI13/MM11_d
+ N_XI57/XI13/NET35_XI57/XI13/MM11_g N_VDD_XI57/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI14/MM2 N_XI57/XI14/NET34_XI57/XI14/MM2_d
+ N_XI57/XI14/NET33_XI57/XI14/MM2_g N_VSS_XI57/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI14/MM3 N_XI57/XI14/NET33_XI57/XI14/MM3_d N_WL<110>_XI57/XI14/MM3_g
+ N_BLN<1>_XI57/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI14/MM0 N_XI57/XI14/NET34_XI57/XI14/MM0_d N_WL<110>_XI57/XI14/MM0_g
+ N_BL<1>_XI57/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI14/MM1 N_XI57/XI14/NET33_XI57/XI14/MM1_d
+ N_XI57/XI14/NET34_XI57/XI14/MM1_g N_VSS_XI57/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI14/MM9 N_XI57/XI14/NET36_XI57/XI14/MM9_d N_WL<111>_XI57/XI14/MM9_g
+ N_BL<1>_XI57/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI14/MM6 N_XI57/XI14/NET35_XI57/XI14/MM6_d
+ N_XI57/XI14/NET36_XI57/XI14/MM6_g N_VSS_XI57/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI14/MM7 N_XI57/XI14/NET36_XI57/XI14/MM7_d
+ N_XI57/XI14/NET35_XI57/XI14/MM7_g N_VSS_XI57/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI14/MM8 N_XI57/XI14/NET35_XI57/XI14/MM8_d N_WL<111>_XI57/XI14/MM8_g
+ N_BLN<1>_XI57/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI14/MM5 N_XI57/XI14/NET34_XI57/XI14/MM5_d
+ N_XI57/XI14/NET33_XI57/XI14/MM5_g N_VDD_XI57/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI14/MM4 N_XI57/XI14/NET33_XI57/XI14/MM4_d
+ N_XI57/XI14/NET34_XI57/XI14/MM4_g N_VDD_XI57/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI14/MM10 N_XI57/XI14/NET35_XI57/XI14/MM10_d
+ N_XI57/XI14/NET36_XI57/XI14/MM10_g N_VDD_XI57/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI14/MM11 N_XI57/XI14/NET36_XI57/XI14/MM11_d
+ N_XI57/XI14/NET35_XI57/XI14/MM11_g N_VDD_XI57/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI15/MM2 N_XI57/XI15/NET34_XI57/XI15/MM2_d
+ N_XI57/XI15/NET33_XI57/XI15/MM2_g N_VSS_XI57/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI15/MM3 N_XI57/XI15/NET33_XI57/XI15/MM3_d N_WL<110>_XI57/XI15/MM3_g
+ N_BLN<0>_XI57/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI15/MM0 N_XI57/XI15/NET34_XI57/XI15/MM0_d N_WL<110>_XI57/XI15/MM0_g
+ N_BL<0>_XI57/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI15/MM1 N_XI57/XI15/NET33_XI57/XI15/MM1_d
+ N_XI57/XI15/NET34_XI57/XI15/MM1_g N_VSS_XI57/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI15/MM9 N_XI57/XI15/NET36_XI57/XI15/MM9_d N_WL<111>_XI57/XI15/MM9_g
+ N_BL<0>_XI57/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI15/MM6 N_XI57/XI15/NET35_XI57/XI15/MM6_d
+ N_XI57/XI15/NET36_XI57/XI15/MM6_g N_VSS_XI57/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI15/MM7 N_XI57/XI15/NET36_XI57/XI15/MM7_d
+ N_XI57/XI15/NET35_XI57/XI15/MM7_g N_VSS_XI57/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI57/XI15/MM8 N_XI57/XI15/NET35_XI57/XI15/MM8_d N_WL<111>_XI57/XI15/MM8_g
+ N_BLN<0>_XI57/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI57/XI15/MM5 N_XI57/XI15/NET34_XI57/XI15/MM5_d
+ N_XI57/XI15/NET33_XI57/XI15/MM5_g N_VDD_XI57/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI15/MM4 N_XI57/XI15/NET33_XI57/XI15/MM4_d
+ N_XI57/XI15/NET34_XI57/XI15/MM4_g N_VDD_XI57/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI15/MM10 N_XI57/XI15/NET35_XI57/XI15/MM10_d
+ N_XI57/XI15/NET36_XI57/XI15/MM10_g N_VDD_XI57/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI57/XI15/MM11 N_XI57/XI15/NET36_XI57/XI15/MM11_d
+ N_XI57/XI15/NET35_XI57/XI15/MM11_g N_VDD_XI57/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI0/MM2 N_XI58/XI0/NET34_XI58/XI0/MM2_d N_XI58/XI0/NET33_XI58/XI0/MM2_g
+ N_VSS_XI58/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI0/MM3 N_XI58/XI0/NET33_XI58/XI0/MM3_d N_WL<112>_XI58/XI0/MM3_g
+ N_BLN<15>_XI58/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI0/MM0 N_XI58/XI0/NET34_XI58/XI0/MM0_d N_WL<112>_XI58/XI0/MM0_g
+ N_BL<15>_XI58/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI0/MM1 N_XI58/XI0/NET33_XI58/XI0/MM1_d N_XI58/XI0/NET34_XI58/XI0/MM1_g
+ N_VSS_XI58/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI0/MM9 N_XI58/XI0/NET36_XI58/XI0/MM9_d N_WL<113>_XI58/XI0/MM9_g
+ N_BL<15>_XI58/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI0/MM6 N_XI58/XI0/NET35_XI58/XI0/MM6_d N_XI58/XI0/NET36_XI58/XI0/MM6_g
+ N_VSS_XI58/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI0/MM7 N_XI58/XI0/NET36_XI58/XI0/MM7_d N_XI58/XI0/NET35_XI58/XI0/MM7_g
+ N_VSS_XI58/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI0/MM8 N_XI58/XI0/NET35_XI58/XI0/MM8_d N_WL<113>_XI58/XI0/MM8_g
+ N_BLN<15>_XI58/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI0/MM5 N_XI58/XI0/NET34_XI58/XI0/MM5_d N_XI58/XI0/NET33_XI58/XI0/MM5_g
+ N_VDD_XI58/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI0/MM4 N_XI58/XI0/NET33_XI58/XI0/MM4_d N_XI58/XI0/NET34_XI58/XI0/MM4_g
+ N_VDD_XI58/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI0/MM10 N_XI58/XI0/NET35_XI58/XI0/MM10_d N_XI58/XI0/NET36_XI58/XI0/MM10_g
+ N_VDD_XI58/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI0/MM11 N_XI58/XI0/NET36_XI58/XI0/MM11_d N_XI58/XI0/NET35_XI58/XI0/MM11_g
+ N_VDD_XI58/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI1/MM2 N_XI58/XI1/NET34_XI58/XI1/MM2_d N_XI58/XI1/NET33_XI58/XI1/MM2_g
+ N_VSS_XI58/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI1/MM3 N_XI58/XI1/NET33_XI58/XI1/MM3_d N_WL<112>_XI58/XI1/MM3_g
+ N_BLN<14>_XI58/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI1/MM0 N_XI58/XI1/NET34_XI58/XI1/MM0_d N_WL<112>_XI58/XI1/MM0_g
+ N_BL<14>_XI58/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI1/MM1 N_XI58/XI1/NET33_XI58/XI1/MM1_d N_XI58/XI1/NET34_XI58/XI1/MM1_g
+ N_VSS_XI58/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI1/MM9 N_XI58/XI1/NET36_XI58/XI1/MM9_d N_WL<113>_XI58/XI1/MM9_g
+ N_BL<14>_XI58/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI1/MM6 N_XI58/XI1/NET35_XI58/XI1/MM6_d N_XI58/XI1/NET36_XI58/XI1/MM6_g
+ N_VSS_XI58/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI1/MM7 N_XI58/XI1/NET36_XI58/XI1/MM7_d N_XI58/XI1/NET35_XI58/XI1/MM7_g
+ N_VSS_XI58/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI1/MM8 N_XI58/XI1/NET35_XI58/XI1/MM8_d N_WL<113>_XI58/XI1/MM8_g
+ N_BLN<14>_XI58/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI1/MM5 N_XI58/XI1/NET34_XI58/XI1/MM5_d N_XI58/XI1/NET33_XI58/XI1/MM5_g
+ N_VDD_XI58/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI1/MM4 N_XI58/XI1/NET33_XI58/XI1/MM4_d N_XI58/XI1/NET34_XI58/XI1/MM4_g
+ N_VDD_XI58/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI1/MM10 N_XI58/XI1/NET35_XI58/XI1/MM10_d N_XI58/XI1/NET36_XI58/XI1/MM10_g
+ N_VDD_XI58/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI1/MM11 N_XI58/XI1/NET36_XI58/XI1/MM11_d N_XI58/XI1/NET35_XI58/XI1/MM11_g
+ N_VDD_XI58/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI2/MM2 N_XI58/XI2/NET34_XI58/XI2/MM2_d N_XI58/XI2/NET33_XI58/XI2/MM2_g
+ N_VSS_XI58/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI2/MM3 N_XI58/XI2/NET33_XI58/XI2/MM3_d N_WL<112>_XI58/XI2/MM3_g
+ N_BLN<13>_XI58/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI2/MM0 N_XI58/XI2/NET34_XI58/XI2/MM0_d N_WL<112>_XI58/XI2/MM0_g
+ N_BL<13>_XI58/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI2/MM1 N_XI58/XI2/NET33_XI58/XI2/MM1_d N_XI58/XI2/NET34_XI58/XI2/MM1_g
+ N_VSS_XI58/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI2/MM9 N_XI58/XI2/NET36_XI58/XI2/MM9_d N_WL<113>_XI58/XI2/MM9_g
+ N_BL<13>_XI58/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI2/MM6 N_XI58/XI2/NET35_XI58/XI2/MM6_d N_XI58/XI2/NET36_XI58/XI2/MM6_g
+ N_VSS_XI58/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI2/MM7 N_XI58/XI2/NET36_XI58/XI2/MM7_d N_XI58/XI2/NET35_XI58/XI2/MM7_g
+ N_VSS_XI58/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI2/MM8 N_XI58/XI2/NET35_XI58/XI2/MM8_d N_WL<113>_XI58/XI2/MM8_g
+ N_BLN<13>_XI58/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI2/MM5 N_XI58/XI2/NET34_XI58/XI2/MM5_d N_XI58/XI2/NET33_XI58/XI2/MM5_g
+ N_VDD_XI58/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI2/MM4 N_XI58/XI2/NET33_XI58/XI2/MM4_d N_XI58/XI2/NET34_XI58/XI2/MM4_g
+ N_VDD_XI58/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI2/MM10 N_XI58/XI2/NET35_XI58/XI2/MM10_d N_XI58/XI2/NET36_XI58/XI2/MM10_g
+ N_VDD_XI58/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI2/MM11 N_XI58/XI2/NET36_XI58/XI2/MM11_d N_XI58/XI2/NET35_XI58/XI2/MM11_g
+ N_VDD_XI58/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI3/MM2 N_XI58/XI3/NET34_XI58/XI3/MM2_d N_XI58/XI3/NET33_XI58/XI3/MM2_g
+ N_VSS_XI58/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI3/MM3 N_XI58/XI3/NET33_XI58/XI3/MM3_d N_WL<112>_XI58/XI3/MM3_g
+ N_BLN<12>_XI58/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI3/MM0 N_XI58/XI3/NET34_XI58/XI3/MM0_d N_WL<112>_XI58/XI3/MM0_g
+ N_BL<12>_XI58/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI3/MM1 N_XI58/XI3/NET33_XI58/XI3/MM1_d N_XI58/XI3/NET34_XI58/XI3/MM1_g
+ N_VSS_XI58/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI3/MM9 N_XI58/XI3/NET36_XI58/XI3/MM9_d N_WL<113>_XI58/XI3/MM9_g
+ N_BL<12>_XI58/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI3/MM6 N_XI58/XI3/NET35_XI58/XI3/MM6_d N_XI58/XI3/NET36_XI58/XI3/MM6_g
+ N_VSS_XI58/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI3/MM7 N_XI58/XI3/NET36_XI58/XI3/MM7_d N_XI58/XI3/NET35_XI58/XI3/MM7_g
+ N_VSS_XI58/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI3/MM8 N_XI58/XI3/NET35_XI58/XI3/MM8_d N_WL<113>_XI58/XI3/MM8_g
+ N_BLN<12>_XI58/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI3/MM5 N_XI58/XI3/NET34_XI58/XI3/MM5_d N_XI58/XI3/NET33_XI58/XI3/MM5_g
+ N_VDD_XI58/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI3/MM4 N_XI58/XI3/NET33_XI58/XI3/MM4_d N_XI58/XI3/NET34_XI58/XI3/MM4_g
+ N_VDD_XI58/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI3/MM10 N_XI58/XI3/NET35_XI58/XI3/MM10_d N_XI58/XI3/NET36_XI58/XI3/MM10_g
+ N_VDD_XI58/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI3/MM11 N_XI58/XI3/NET36_XI58/XI3/MM11_d N_XI58/XI3/NET35_XI58/XI3/MM11_g
+ N_VDD_XI58/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI4/MM2 N_XI58/XI4/NET34_XI58/XI4/MM2_d N_XI58/XI4/NET33_XI58/XI4/MM2_g
+ N_VSS_XI58/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI4/MM3 N_XI58/XI4/NET33_XI58/XI4/MM3_d N_WL<112>_XI58/XI4/MM3_g
+ N_BLN<11>_XI58/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI4/MM0 N_XI58/XI4/NET34_XI58/XI4/MM0_d N_WL<112>_XI58/XI4/MM0_g
+ N_BL<11>_XI58/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI4/MM1 N_XI58/XI4/NET33_XI58/XI4/MM1_d N_XI58/XI4/NET34_XI58/XI4/MM1_g
+ N_VSS_XI58/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI4/MM9 N_XI58/XI4/NET36_XI58/XI4/MM9_d N_WL<113>_XI58/XI4/MM9_g
+ N_BL<11>_XI58/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI4/MM6 N_XI58/XI4/NET35_XI58/XI4/MM6_d N_XI58/XI4/NET36_XI58/XI4/MM6_g
+ N_VSS_XI58/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI4/MM7 N_XI58/XI4/NET36_XI58/XI4/MM7_d N_XI58/XI4/NET35_XI58/XI4/MM7_g
+ N_VSS_XI58/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI4/MM8 N_XI58/XI4/NET35_XI58/XI4/MM8_d N_WL<113>_XI58/XI4/MM8_g
+ N_BLN<11>_XI58/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI4/MM5 N_XI58/XI4/NET34_XI58/XI4/MM5_d N_XI58/XI4/NET33_XI58/XI4/MM5_g
+ N_VDD_XI58/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI4/MM4 N_XI58/XI4/NET33_XI58/XI4/MM4_d N_XI58/XI4/NET34_XI58/XI4/MM4_g
+ N_VDD_XI58/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI4/MM10 N_XI58/XI4/NET35_XI58/XI4/MM10_d N_XI58/XI4/NET36_XI58/XI4/MM10_g
+ N_VDD_XI58/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI4/MM11 N_XI58/XI4/NET36_XI58/XI4/MM11_d N_XI58/XI4/NET35_XI58/XI4/MM11_g
+ N_VDD_XI58/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI5/MM2 N_XI58/XI5/NET34_XI58/XI5/MM2_d N_XI58/XI5/NET33_XI58/XI5/MM2_g
+ N_VSS_XI58/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI5/MM3 N_XI58/XI5/NET33_XI58/XI5/MM3_d N_WL<112>_XI58/XI5/MM3_g
+ N_BLN<10>_XI58/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI5/MM0 N_XI58/XI5/NET34_XI58/XI5/MM0_d N_WL<112>_XI58/XI5/MM0_g
+ N_BL<10>_XI58/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI5/MM1 N_XI58/XI5/NET33_XI58/XI5/MM1_d N_XI58/XI5/NET34_XI58/XI5/MM1_g
+ N_VSS_XI58/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI5/MM9 N_XI58/XI5/NET36_XI58/XI5/MM9_d N_WL<113>_XI58/XI5/MM9_g
+ N_BL<10>_XI58/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI5/MM6 N_XI58/XI5/NET35_XI58/XI5/MM6_d N_XI58/XI5/NET36_XI58/XI5/MM6_g
+ N_VSS_XI58/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI5/MM7 N_XI58/XI5/NET36_XI58/XI5/MM7_d N_XI58/XI5/NET35_XI58/XI5/MM7_g
+ N_VSS_XI58/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI5/MM8 N_XI58/XI5/NET35_XI58/XI5/MM8_d N_WL<113>_XI58/XI5/MM8_g
+ N_BLN<10>_XI58/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI5/MM5 N_XI58/XI5/NET34_XI58/XI5/MM5_d N_XI58/XI5/NET33_XI58/XI5/MM5_g
+ N_VDD_XI58/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI5/MM4 N_XI58/XI5/NET33_XI58/XI5/MM4_d N_XI58/XI5/NET34_XI58/XI5/MM4_g
+ N_VDD_XI58/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI5/MM10 N_XI58/XI5/NET35_XI58/XI5/MM10_d N_XI58/XI5/NET36_XI58/XI5/MM10_g
+ N_VDD_XI58/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI5/MM11 N_XI58/XI5/NET36_XI58/XI5/MM11_d N_XI58/XI5/NET35_XI58/XI5/MM11_g
+ N_VDD_XI58/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI6/MM2 N_XI58/XI6/NET34_XI58/XI6/MM2_d N_XI58/XI6/NET33_XI58/XI6/MM2_g
+ N_VSS_XI58/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM3 N_XI58/XI6/NET33_XI58/XI6/MM3_d N_WL<112>_XI58/XI6/MM3_g
+ N_BLN<9>_XI58/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM0 N_XI58/XI6/NET34_XI58/XI6/MM0_d N_WL<112>_XI58/XI6/MM0_g
+ N_BL<9>_XI58/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM1 N_XI58/XI6/NET33_XI58/XI6/MM1_d N_XI58/XI6/NET34_XI58/XI6/MM1_g
+ N_VSS_XI58/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM9 N_XI58/XI6/NET36_XI58/XI6/MM9_d N_WL<113>_XI58/XI6/MM9_g
+ N_BL<9>_XI58/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM6 N_XI58/XI6/NET35_XI58/XI6/MM6_d N_XI58/XI6/NET36_XI58/XI6/MM6_g
+ N_VSS_XI58/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM7 N_XI58/XI6/NET36_XI58/XI6/MM7_d N_XI58/XI6/NET35_XI58/XI6/MM7_g
+ N_VSS_XI58/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM8 N_XI58/XI6/NET35_XI58/XI6/MM8_d N_WL<113>_XI58/XI6/MM8_g
+ N_BLN<9>_XI58/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI6/MM5 N_XI58/XI6/NET34_XI58/XI6/MM5_d N_XI58/XI6/NET33_XI58/XI6/MM5_g
+ N_VDD_XI58/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI6/MM4 N_XI58/XI6/NET33_XI58/XI6/MM4_d N_XI58/XI6/NET34_XI58/XI6/MM4_g
+ N_VDD_XI58/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI6/MM10 N_XI58/XI6/NET35_XI58/XI6/MM10_d N_XI58/XI6/NET36_XI58/XI6/MM10_g
+ N_VDD_XI58/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI6/MM11 N_XI58/XI6/NET36_XI58/XI6/MM11_d N_XI58/XI6/NET35_XI58/XI6/MM11_g
+ N_VDD_XI58/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI7/MM2 N_XI58/XI7/NET34_XI58/XI7/MM2_d N_XI58/XI7/NET33_XI58/XI7/MM2_g
+ N_VSS_XI58/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM3 N_XI58/XI7/NET33_XI58/XI7/MM3_d N_WL<112>_XI58/XI7/MM3_g
+ N_BLN<8>_XI58/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM0 N_XI58/XI7/NET34_XI58/XI7/MM0_d N_WL<112>_XI58/XI7/MM0_g
+ N_BL<8>_XI58/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM1 N_XI58/XI7/NET33_XI58/XI7/MM1_d N_XI58/XI7/NET34_XI58/XI7/MM1_g
+ N_VSS_XI58/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM9 N_XI58/XI7/NET36_XI58/XI7/MM9_d N_WL<113>_XI58/XI7/MM9_g
+ N_BL<8>_XI58/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM6 N_XI58/XI7/NET35_XI58/XI7/MM6_d N_XI58/XI7/NET36_XI58/XI7/MM6_g
+ N_VSS_XI58/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM7 N_XI58/XI7/NET36_XI58/XI7/MM7_d N_XI58/XI7/NET35_XI58/XI7/MM7_g
+ N_VSS_XI58/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM8 N_XI58/XI7/NET35_XI58/XI7/MM8_d N_WL<113>_XI58/XI7/MM8_g
+ N_BLN<8>_XI58/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI7/MM5 N_XI58/XI7/NET34_XI58/XI7/MM5_d N_XI58/XI7/NET33_XI58/XI7/MM5_g
+ N_VDD_XI58/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI7/MM4 N_XI58/XI7/NET33_XI58/XI7/MM4_d N_XI58/XI7/NET34_XI58/XI7/MM4_g
+ N_VDD_XI58/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI7/MM10 N_XI58/XI7/NET35_XI58/XI7/MM10_d N_XI58/XI7/NET36_XI58/XI7/MM10_g
+ N_VDD_XI58/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI7/MM11 N_XI58/XI7/NET36_XI58/XI7/MM11_d N_XI58/XI7/NET35_XI58/XI7/MM11_g
+ N_VDD_XI58/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI8/MM2 N_XI58/XI8/NET34_XI58/XI8/MM2_d N_XI58/XI8/NET33_XI58/XI8/MM2_g
+ N_VSS_XI58/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM3 N_XI58/XI8/NET33_XI58/XI8/MM3_d N_WL<112>_XI58/XI8/MM3_g
+ N_BLN<7>_XI58/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM0 N_XI58/XI8/NET34_XI58/XI8/MM0_d N_WL<112>_XI58/XI8/MM0_g
+ N_BL<7>_XI58/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM1 N_XI58/XI8/NET33_XI58/XI8/MM1_d N_XI58/XI8/NET34_XI58/XI8/MM1_g
+ N_VSS_XI58/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM9 N_XI58/XI8/NET36_XI58/XI8/MM9_d N_WL<113>_XI58/XI8/MM9_g
+ N_BL<7>_XI58/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM6 N_XI58/XI8/NET35_XI58/XI8/MM6_d N_XI58/XI8/NET36_XI58/XI8/MM6_g
+ N_VSS_XI58/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM7 N_XI58/XI8/NET36_XI58/XI8/MM7_d N_XI58/XI8/NET35_XI58/XI8/MM7_g
+ N_VSS_XI58/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM8 N_XI58/XI8/NET35_XI58/XI8/MM8_d N_WL<113>_XI58/XI8/MM8_g
+ N_BLN<7>_XI58/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI8/MM5 N_XI58/XI8/NET34_XI58/XI8/MM5_d N_XI58/XI8/NET33_XI58/XI8/MM5_g
+ N_VDD_XI58/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI8/MM4 N_XI58/XI8/NET33_XI58/XI8/MM4_d N_XI58/XI8/NET34_XI58/XI8/MM4_g
+ N_VDD_XI58/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI8/MM10 N_XI58/XI8/NET35_XI58/XI8/MM10_d N_XI58/XI8/NET36_XI58/XI8/MM10_g
+ N_VDD_XI58/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI8/MM11 N_XI58/XI8/NET36_XI58/XI8/MM11_d N_XI58/XI8/NET35_XI58/XI8/MM11_g
+ N_VDD_XI58/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI9/MM2 N_XI58/XI9/NET34_XI58/XI9/MM2_d N_XI58/XI9/NET33_XI58/XI9/MM2_g
+ N_VSS_XI58/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM3 N_XI58/XI9/NET33_XI58/XI9/MM3_d N_WL<112>_XI58/XI9/MM3_g
+ N_BLN<6>_XI58/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM0 N_XI58/XI9/NET34_XI58/XI9/MM0_d N_WL<112>_XI58/XI9/MM0_g
+ N_BL<6>_XI58/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM1 N_XI58/XI9/NET33_XI58/XI9/MM1_d N_XI58/XI9/NET34_XI58/XI9/MM1_g
+ N_VSS_XI58/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM9 N_XI58/XI9/NET36_XI58/XI9/MM9_d N_WL<113>_XI58/XI9/MM9_g
+ N_BL<6>_XI58/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM6 N_XI58/XI9/NET35_XI58/XI9/MM6_d N_XI58/XI9/NET36_XI58/XI9/MM6_g
+ N_VSS_XI58/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM7 N_XI58/XI9/NET36_XI58/XI9/MM7_d N_XI58/XI9/NET35_XI58/XI9/MM7_g
+ N_VSS_XI58/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM8 N_XI58/XI9/NET35_XI58/XI9/MM8_d N_WL<113>_XI58/XI9/MM8_g
+ N_BLN<6>_XI58/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI9/MM5 N_XI58/XI9/NET34_XI58/XI9/MM5_d N_XI58/XI9/NET33_XI58/XI9/MM5_g
+ N_VDD_XI58/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI9/MM4 N_XI58/XI9/NET33_XI58/XI9/MM4_d N_XI58/XI9/NET34_XI58/XI9/MM4_g
+ N_VDD_XI58/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI9/MM10 N_XI58/XI9/NET35_XI58/XI9/MM10_d N_XI58/XI9/NET36_XI58/XI9/MM10_g
+ N_VDD_XI58/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI9/MM11 N_XI58/XI9/NET36_XI58/XI9/MM11_d N_XI58/XI9/NET35_XI58/XI9/MM11_g
+ N_VDD_XI58/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI10/MM2 N_XI58/XI10/NET34_XI58/XI10/MM2_d
+ N_XI58/XI10/NET33_XI58/XI10/MM2_g N_VSS_XI58/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI10/MM3 N_XI58/XI10/NET33_XI58/XI10/MM3_d N_WL<112>_XI58/XI10/MM3_g
+ N_BLN<5>_XI58/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI10/MM0 N_XI58/XI10/NET34_XI58/XI10/MM0_d N_WL<112>_XI58/XI10/MM0_g
+ N_BL<5>_XI58/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI10/MM1 N_XI58/XI10/NET33_XI58/XI10/MM1_d
+ N_XI58/XI10/NET34_XI58/XI10/MM1_g N_VSS_XI58/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI10/MM9 N_XI58/XI10/NET36_XI58/XI10/MM9_d N_WL<113>_XI58/XI10/MM9_g
+ N_BL<5>_XI58/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI10/MM6 N_XI58/XI10/NET35_XI58/XI10/MM6_d
+ N_XI58/XI10/NET36_XI58/XI10/MM6_g N_VSS_XI58/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI10/MM7 N_XI58/XI10/NET36_XI58/XI10/MM7_d
+ N_XI58/XI10/NET35_XI58/XI10/MM7_g N_VSS_XI58/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI10/MM8 N_XI58/XI10/NET35_XI58/XI10/MM8_d N_WL<113>_XI58/XI10/MM8_g
+ N_BLN<5>_XI58/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI10/MM5 N_XI58/XI10/NET34_XI58/XI10/MM5_d
+ N_XI58/XI10/NET33_XI58/XI10/MM5_g N_VDD_XI58/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI10/MM4 N_XI58/XI10/NET33_XI58/XI10/MM4_d
+ N_XI58/XI10/NET34_XI58/XI10/MM4_g N_VDD_XI58/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI10/MM10 N_XI58/XI10/NET35_XI58/XI10/MM10_d
+ N_XI58/XI10/NET36_XI58/XI10/MM10_g N_VDD_XI58/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI10/MM11 N_XI58/XI10/NET36_XI58/XI10/MM11_d
+ N_XI58/XI10/NET35_XI58/XI10/MM11_g N_VDD_XI58/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI11/MM2 N_XI58/XI11/NET34_XI58/XI11/MM2_d
+ N_XI58/XI11/NET33_XI58/XI11/MM2_g N_VSS_XI58/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI11/MM3 N_XI58/XI11/NET33_XI58/XI11/MM3_d N_WL<112>_XI58/XI11/MM3_g
+ N_BLN<4>_XI58/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI11/MM0 N_XI58/XI11/NET34_XI58/XI11/MM0_d N_WL<112>_XI58/XI11/MM0_g
+ N_BL<4>_XI58/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI11/MM1 N_XI58/XI11/NET33_XI58/XI11/MM1_d
+ N_XI58/XI11/NET34_XI58/XI11/MM1_g N_VSS_XI58/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI11/MM9 N_XI58/XI11/NET36_XI58/XI11/MM9_d N_WL<113>_XI58/XI11/MM9_g
+ N_BL<4>_XI58/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI11/MM6 N_XI58/XI11/NET35_XI58/XI11/MM6_d
+ N_XI58/XI11/NET36_XI58/XI11/MM6_g N_VSS_XI58/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI11/MM7 N_XI58/XI11/NET36_XI58/XI11/MM7_d
+ N_XI58/XI11/NET35_XI58/XI11/MM7_g N_VSS_XI58/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI11/MM8 N_XI58/XI11/NET35_XI58/XI11/MM8_d N_WL<113>_XI58/XI11/MM8_g
+ N_BLN<4>_XI58/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI11/MM5 N_XI58/XI11/NET34_XI58/XI11/MM5_d
+ N_XI58/XI11/NET33_XI58/XI11/MM5_g N_VDD_XI58/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI11/MM4 N_XI58/XI11/NET33_XI58/XI11/MM4_d
+ N_XI58/XI11/NET34_XI58/XI11/MM4_g N_VDD_XI58/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI11/MM10 N_XI58/XI11/NET35_XI58/XI11/MM10_d
+ N_XI58/XI11/NET36_XI58/XI11/MM10_g N_VDD_XI58/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI11/MM11 N_XI58/XI11/NET36_XI58/XI11/MM11_d
+ N_XI58/XI11/NET35_XI58/XI11/MM11_g N_VDD_XI58/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI12/MM2 N_XI58/XI12/NET34_XI58/XI12/MM2_d
+ N_XI58/XI12/NET33_XI58/XI12/MM2_g N_VSS_XI58/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI12/MM3 N_XI58/XI12/NET33_XI58/XI12/MM3_d N_WL<112>_XI58/XI12/MM3_g
+ N_BLN<3>_XI58/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI12/MM0 N_XI58/XI12/NET34_XI58/XI12/MM0_d N_WL<112>_XI58/XI12/MM0_g
+ N_BL<3>_XI58/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI12/MM1 N_XI58/XI12/NET33_XI58/XI12/MM1_d
+ N_XI58/XI12/NET34_XI58/XI12/MM1_g N_VSS_XI58/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI12/MM9 N_XI58/XI12/NET36_XI58/XI12/MM9_d N_WL<113>_XI58/XI12/MM9_g
+ N_BL<3>_XI58/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI12/MM6 N_XI58/XI12/NET35_XI58/XI12/MM6_d
+ N_XI58/XI12/NET36_XI58/XI12/MM6_g N_VSS_XI58/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI12/MM7 N_XI58/XI12/NET36_XI58/XI12/MM7_d
+ N_XI58/XI12/NET35_XI58/XI12/MM7_g N_VSS_XI58/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI12/MM8 N_XI58/XI12/NET35_XI58/XI12/MM8_d N_WL<113>_XI58/XI12/MM8_g
+ N_BLN<3>_XI58/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI12/MM5 N_XI58/XI12/NET34_XI58/XI12/MM5_d
+ N_XI58/XI12/NET33_XI58/XI12/MM5_g N_VDD_XI58/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI12/MM4 N_XI58/XI12/NET33_XI58/XI12/MM4_d
+ N_XI58/XI12/NET34_XI58/XI12/MM4_g N_VDD_XI58/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI12/MM10 N_XI58/XI12/NET35_XI58/XI12/MM10_d
+ N_XI58/XI12/NET36_XI58/XI12/MM10_g N_VDD_XI58/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI12/MM11 N_XI58/XI12/NET36_XI58/XI12/MM11_d
+ N_XI58/XI12/NET35_XI58/XI12/MM11_g N_VDD_XI58/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI13/MM2 N_XI58/XI13/NET34_XI58/XI13/MM2_d
+ N_XI58/XI13/NET33_XI58/XI13/MM2_g N_VSS_XI58/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI13/MM3 N_XI58/XI13/NET33_XI58/XI13/MM3_d N_WL<112>_XI58/XI13/MM3_g
+ N_BLN<2>_XI58/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI13/MM0 N_XI58/XI13/NET34_XI58/XI13/MM0_d N_WL<112>_XI58/XI13/MM0_g
+ N_BL<2>_XI58/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI13/MM1 N_XI58/XI13/NET33_XI58/XI13/MM1_d
+ N_XI58/XI13/NET34_XI58/XI13/MM1_g N_VSS_XI58/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI13/MM9 N_XI58/XI13/NET36_XI58/XI13/MM9_d N_WL<113>_XI58/XI13/MM9_g
+ N_BL<2>_XI58/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI13/MM6 N_XI58/XI13/NET35_XI58/XI13/MM6_d
+ N_XI58/XI13/NET36_XI58/XI13/MM6_g N_VSS_XI58/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI13/MM7 N_XI58/XI13/NET36_XI58/XI13/MM7_d
+ N_XI58/XI13/NET35_XI58/XI13/MM7_g N_VSS_XI58/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI13/MM8 N_XI58/XI13/NET35_XI58/XI13/MM8_d N_WL<113>_XI58/XI13/MM8_g
+ N_BLN<2>_XI58/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI13/MM5 N_XI58/XI13/NET34_XI58/XI13/MM5_d
+ N_XI58/XI13/NET33_XI58/XI13/MM5_g N_VDD_XI58/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI13/MM4 N_XI58/XI13/NET33_XI58/XI13/MM4_d
+ N_XI58/XI13/NET34_XI58/XI13/MM4_g N_VDD_XI58/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI13/MM10 N_XI58/XI13/NET35_XI58/XI13/MM10_d
+ N_XI58/XI13/NET36_XI58/XI13/MM10_g N_VDD_XI58/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI13/MM11 N_XI58/XI13/NET36_XI58/XI13/MM11_d
+ N_XI58/XI13/NET35_XI58/XI13/MM11_g N_VDD_XI58/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI14/MM2 N_XI58/XI14/NET34_XI58/XI14/MM2_d
+ N_XI58/XI14/NET33_XI58/XI14/MM2_g N_VSS_XI58/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI14/MM3 N_XI58/XI14/NET33_XI58/XI14/MM3_d N_WL<112>_XI58/XI14/MM3_g
+ N_BLN<1>_XI58/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI14/MM0 N_XI58/XI14/NET34_XI58/XI14/MM0_d N_WL<112>_XI58/XI14/MM0_g
+ N_BL<1>_XI58/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI14/MM1 N_XI58/XI14/NET33_XI58/XI14/MM1_d
+ N_XI58/XI14/NET34_XI58/XI14/MM1_g N_VSS_XI58/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI14/MM9 N_XI58/XI14/NET36_XI58/XI14/MM9_d N_WL<113>_XI58/XI14/MM9_g
+ N_BL<1>_XI58/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI14/MM6 N_XI58/XI14/NET35_XI58/XI14/MM6_d
+ N_XI58/XI14/NET36_XI58/XI14/MM6_g N_VSS_XI58/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI14/MM7 N_XI58/XI14/NET36_XI58/XI14/MM7_d
+ N_XI58/XI14/NET35_XI58/XI14/MM7_g N_VSS_XI58/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI14/MM8 N_XI58/XI14/NET35_XI58/XI14/MM8_d N_WL<113>_XI58/XI14/MM8_g
+ N_BLN<1>_XI58/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI14/MM5 N_XI58/XI14/NET34_XI58/XI14/MM5_d
+ N_XI58/XI14/NET33_XI58/XI14/MM5_g N_VDD_XI58/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI14/MM4 N_XI58/XI14/NET33_XI58/XI14/MM4_d
+ N_XI58/XI14/NET34_XI58/XI14/MM4_g N_VDD_XI58/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI14/MM10 N_XI58/XI14/NET35_XI58/XI14/MM10_d
+ N_XI58/XI14/NET36_XI58/XI14/MM10_g N_VDD_XI58/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI14/MM11 N_XI58/XI14/NET36_XI58/XI14/MM11_d
+ N_XI58/XI14/NET35_XI58/XI14/MM11_g N_VDD_XI58/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI15/MM2 N_XI58/XI15/NET34_XI58/XI15/MM2_d
+ N_XI58/XI15/NET33_XI58/XI15/MM2_g N_VSS_XI58/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI15/MM3 N_XI58/XI15/NET33_XI58/XI15/MM3_d N_WL<112>_XI58/XI15/MM3_g
+ N_BLN<0>_XI58/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI15/MM0 N_XI58/XI15/NET34_XI58/XI15/MM0_d N_WL<112>_XI58/XI15/MM0_g
+ N_BL<0>_XI58/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI15/MM1 N_XI58/XI15/NET33_XI58/XI15/MM1_d
+ N_XI58/XI15/NET34_XI58/XI15/MM1_g N_VSS_XI58/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI15/MM9 N_XI58/XI15/NET36_XI58/XI15/MM9_d N_WL<113>_XI58/XI15/MM9_g
+ N_BL<0>_XI58/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI15/MM6 N_XI58/XI15/NET35_XI58/XI15/MM6_d
+ N_XI58/XI15/NET36_XI58/XI15/MM6_g N_VSS_XI58/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI15/MM7 N_XI58/XI15/NET36_XI58/XI15/MM7_d
+ N_XI58/XI15/NET35_XI58/XI15/MM7_g N_VSS_XI58/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI58/XI15/MM8 N_XI58/XI15/NET35_XI58/XI15/MM8_d N_WL<113>_XI58/XI15/MM8_g
+ N_BLN<0>_XI58/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI58/XI15/MM5 N_XI58/XI15/NET34_XI58/XI15/MM5_d
+ N_XI58/XI15/NET33_XI58/XI15/MM5_g N_VDD_XI58/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI15/MM4 N_XI58/XI15/NET33_XI58/XI15/MM4_d
+ N_XI58/XI15/NET34_XI58/XI15/MM4_g N_VDD_XI58/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI15/MM10 N_XI58/XI15/NET35_XI58/XI15/MM10_d
+ N_XI58/XI15/NET36_XI58/XI15/MM10_g N_VDD_XI58/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI58/XI15/MM11 N_XI58/XI15/NET36_XI58/XI15/MM11_d
+ N_XI58/XI15/NET35_XI58/XI15/MM11_g N_VDD_XI58/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI0/MM2 N_XI59/XI0/NET34_XI59/XI0/MM2_d N_XI59/XI0/NET33_XI59/XI0/MM2_g
+ N_VSS_XI59/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI0/MM3 N_XI59/XI0/NET33_XI59/XI0/MM3_d N_WL<114>_XI59/XI0/MM3_g
+ N_BLN<15>_XI59/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI0/MM0 N_XI59/XI0/NET34_XI59/XI0/MM0_d N_WL<114>_XI59/XI0/MM0_g
+ N_BL<15>_XI59/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI0/MM1 N_XI59/XI0/NET33_XI59/XI0/MM1_d N_XI59/XI0/NET34_XI59/XI0/MM1_g
+ N_VSS_XI59/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI0/MM9 N_XI59/XI0/NET36_XI59/XI0/MM9_d N_WL<115>_XI59/XI0/MM9_g
+ N_BL<15>_XI59/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI0/MM6 N_XI59/XI0/NET35_XI59/XI0/MM6_d N_XI59/XI0/NET36_XI59/XI0/MM6_g
+ N_VSS_XI59/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI0/MM7 N_XI59/XI0/NET36_XI59/XI0/MM7_d N_XI59/XI0/NET35_XI59/XI0/MM7_g
+ N_VSS_XI59/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI0/MM8 N_XI59/XI0/NET35_XI59/XI0/MM8_d N_WL<115>_XI59/XI0/MM8_g
+ N_BLN<15>_XI59/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI0/MM5 N_XI59/XI0/NET34_XI59/XI0/MM5_d N_XI59/XI0/NET33_XI59/XI0/MM5_g
+ N_VDD_XI59/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI0/MM4 N_XI59/XI0/NET33_XI59/XI0/MM4_d N_XI59/XI0/NET34_XI59/XI0/MM4_g
+ N_VDD_XI59/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI0/MM10 N_XI59/XI0/NET35_XI59/XI0/MM10_d N_XI59/XI0/NET36_XI59/XI0/MM10_g
+ N_VDD_XI59/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI0/MM11 N_XI59/XI0/NET36_XI59/XI0/MM11_d N_XI59/XI0/NET35_XI59/XI0/MM11_g
+ N_VDD_XI59/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI1/MM2 N_XI59/XI1/NET34_XI59/XI1/MM2_d N_XI59/XI1/NET33_XI59/XI1/MM2_g
+ N_VSS_XI59/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI1/MM3 N_XI59/XI1/NET33_XI59/XI1/MM3_d N_WL<114>_XI59/XI1/MM3_g
+ N_BLN<14>_XI59/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI1/MM0 N_XI59/XI1/NET34_XI59/XI1/MM0_d N_WL<114>_XI59/XI1/MM0_g
+ N_BL<14>_XI59/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI1/MM1 N_XI59/XI1/NET33_XI59/XI1/MM1_d N_XI59/XI1/NET34_XI59/XI1/MM1_g
+ N_VSS_XI59/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI1/MM9 N_XI59/XI1/NET36_XI59/XI1/MM9_d N_WL<115>_XI59/XI1/MM9_g
+ N_BL<14>_XI59/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI1/MM6 N_XI59/XI1/NET35_XI59/XI1/MM6_d N_XI59/XI1/NET36_XI59/XI1/MM6_g
+ N_VSS_XI59/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI1/MM7 N_XI59/XI1/NET36_XI59/XI1/MM7_d N_XI59/XI1/NET35_XI59/XI1/MM7_g
+ N_VSS_XI59/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI1/MM8 N_XI59/XI1/NET35_XI59/XI1/MM8_d N_WL<115>_XI59/XI1/MM8_g
+ N_BLN<14>_XI59/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI1/MM5 N_XI59/XI1/NET34_XI59/XI1/MM5_d N_XI59/XI1/NET33_XI59/XI1/MM5_g
+ N_VDD_XI59/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI1/MM4 N_XI59/XI1/NET33_XI59/XI1/MM4_d N_XI59/XI1/NET34_XI59/XI1/MM4_g
+ N_VDD_XI59/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI1/MM10 N_XI59/XI1/NET35_XI59/XI1/MM10_d N_XI59/XI1/NET36_XI59/XI1/MM10_g
+ N_VDD_XI59/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI1/MM11 N_XI59/XI1/NET36_XI59/XI1/MM11_d N_XI59/XI1/NET35_XI59/XI1/MM11_g
+ N_VDD_XI59/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI2/MM2 N_XI59/XI2/NET34_XI59/XI2/MM2_d N_XI59/XI2/NET33_XI59/XI2/MM2_g
+ N_VSS_XI59/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI2/MM3 N_XI59/XI2/NET33_XI59/XI2/MM3_d N_WL<114>_XI59/XI2/MM3_g
+ N_BLN<13>_XI59/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI2/MM0 N_XI59/XI2/NET34_XI59/XI2/MM0_d N_WL<114>_XI59/XI2/MM0_g
+ N_BL<13>_XI59/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI2/MM1 N_XI59/XI2/NET33_XI59/XI2/MM1_d N_XI59/XI2/NET34_XI59/XI2/MM1_g
+ N_VSS_XI59/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI2/MM9 N_XI59/XI2/NET36_XI59/XI2/MM9_d N_WL<115>_XI59/XI2/MM9_g
+ N_BL<13>_XI59/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI2/MM6 N_XI59/XI2/NET35_XI59/XI2/MM6_d N_XI59/XI2/NET36_XI59/XI2/MM6_g
+ N_VSS_XI59/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI2/MM7 N_XI59/XI2/NET36_XI59/XI2/MM7_d N_XI59/XI2/NET35_XI59/XI2/MM7_g
+ N_VSS_XI59/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI2/MM8 N_XI59/XI2/NET35_XI59/XI2/MM8_d N_WL<115>_XI59/XI2/MM8_g
+ N_BLN<13>_XI59/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI2/MM5 N_XI59/XI2/NET34_XI59/XI2/MM5_d N_XI59/XI2/NET33_XI59/XI2/MM5_g
+ N_VDD_XI59/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI2/MM4 N_XI59/XI2/NET33_XI59/XI2/MM4_d N_XI59/XI2/NET34_XI59/XI2/MM4_g
+ N_VDD_XI59/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI2/MM10 N_XI59/XI2/NET35_XI59/XI2/MM10_d N_XI59/XI2/NET36_XI59/XI2/MM10_g
+ N_VDD_XI59/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI2/MM11 N_XI59/XI2/NET36_XI59/XI2/MM11_d N_XI59/XI2/NET35_XI59/XI2/MM11_g
+ N_VDD_XI59/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI3/MM2 N_XI59/XI3/NET34_XI59/XI3/MM2_d N_XI59/XI3/NET33_XI59/XI3/MM2_g
+ N_VSS_XI59/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI3/MM3 N_XI59/XI3/NET33_XI59/XI3/MM3_d N_WL<114>_XI59/XI3/MM3_g
+ N_BLN<12>_XI59/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI3/MM0 N_XI59/XI3/NET34_XI59/XI3/MM0_d N_WL<114>_XI59/XI3/MM0_g
+ N_BL<12>_XI59/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI3/MM1 N_XI59/XI3/NET33_XI59/XI3/MM1_d N_XI59/XI3/NET34_XI59/XI3/MM1_g
+ N_VSS_XI59/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI3/MM9 N_XI59/XI3/NET36_XI59/XI3/MM9_d N_WL<115>_XI59/XI3/MM9_g
+ N_BL<12>_XI59/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI3/MM6 N_XI59/XI3/NET35_XI59/XI3/MM6_d N_XI59/XI3/NET36_XI59/XI3/MM6_g
+ N_VSS_XI59/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI3/MM7 N_XI59/XI3/NET36_XI59/XI3/MM7_d N_XI59/XI3/NET35_XI59/XI3/MM7_g
+ N_VSS_XI59/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI3/MM8 N_XI59/XI3/NET35_XI59/XI3/MM8_d N_WL<115>_XI59/XI3/MM8_g
+ N_BLN<12>_XI59/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI3/MM5 N_XI59/XI3/NET34_XI59/XI3/MM5_d N_XI59/XI3/NET33_XI59/XI3/MM5_g
+ N_VDD_XI59/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI3/MM4 N_XI59/XI3/NET33_XI59/XI3/MM4_d N_XI59/XI3/NET34_XI59/XI3/MM4_g
+ N_VDD_XI59/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI3/MM10 N_XI59/XI3/NET35_XI59/XI3/MM10_d N_XI59/XI3/NET36_XI59/XI3/MM10_g
+ N_VDD_XI59/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI3/MM11 N_XI59/XI3/NET36_XI59/XI3/MM11_d N_XI59/XI3/NET35_XI59/XI3/MM11_g
+ N_VDD_XI59/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI4/MM2 N_XI59/XI4/NET34_XI59/XI4/MM2_d N_XI59/XI4/NET33_XI59/XI4/MM2_g
+ N_VSS_XI59/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI4/MM3 N_XI59/XI4/NET33_XI59/XI4/MM3_d N_WL<114>_XI59/XI4/MM3_g
+ N_BLN<11>_XI59/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI4/MM0 N_XI59/XI4/NET34_XI59/XI4/MM0_d N_WL<114>_XI59/XI4/MM0_g
+ N_BL<11>_XI59/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI4/MM1 N_XI59/XI4/NET33_XI59/XI4/MM1_d N_XI59/XI4/NET34_XI59/XI4/MM1_g
+ N_VSS_XI59/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI4/MM9 N_XI59/XI4/NET36_XI59/XI4/MM9_d N_WL<115>_XI59/XI4/MM9_g
+ N_BL<11>_XI59/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI4/MM6 N_XI59/XI4/NET35_XI59/XI4/MM6_d N_XI59/XI4/NET36_XI59/XI4/MM6_g
+ N_VSS_XI59/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI4/MM7 N_XI59/XI4/NET36_XI59/XI4/MM7_d N_XI59/XI4/NET35_XI59/XI4/MM7_g
+ N_VSS_XI59/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI4/MM8 N_XI59/XI4/NET35_XI59/XI4/MM8_d N_WL<115>_XI59/XI4/MM8_g
+ N_BLN<11>_XI59/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI4/MM5 N_XI59/XI4/NET34_XI59/XI4/MM5_d N_XI59/XI4/NET33_XI59/XI4/MM5_g
+ N_VDD_XI59/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI4/MM4 N_XI59/XI4/NET33_XI59/XI4/MM4_d N_XI59/XI4/NET34_XI59/XI4/MM4_g
+ N_VDD_XI59/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI4/MM10 N_XI59/XI4/NET35_XI59/XI4/MM10_d N_XI59/XI4/NET36_XI59/XI4/MM10_g
+ N_VDD_XI59/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI4/MM11 N_XI59/XI4/NET36_XI59/XI4/MM11_d N_XI59/XI4/NET35_XI59/XI4/MM11_g
+ N_VDD_XI59/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI5/MM2 N_XI59/XI5/NET34_XI59/XI5/MM2_d N_XI59/XI5/NET33_XI59/XI5/MM2_g
+ N_VSS_XI59/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI5/MM3 N_XI59/XI5/NET33_XI59/XI5/MM3_d N_WL<114>_XI59/XI5/MM3_g
+ N_BLN<10>_XI59/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI5/MM0 N_XI59/XI5/NET34_XI59/XI5/MM0_d N_WL<114>_XI59/XI5/MM0_g
+ N_BL<10>_XI59/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI5/MM1 N_XI59/XI5/NET33_XI59/XI5/MM1_d N_XI59/XI5/NET34_XI59/XI5/MM1_g
+ N_VSS_XI59/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI5/MM9 N_XI59/XI5/NET36_XI59/XI5/MM9_d N_WL<115>_XI59/XI5/MM9_g
+ N_BL<10>_XI59/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI5/MM6 N_XI59/XI5/NET35_XI59/XI5/MM6_d N_XI59/XI5/NET36_XI59/XI5/MM6_g
+ N_VSS_XI59/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI5/MM7 N_XI59/XI5/NET36_XI59/XI5/MM7_d N_XI59/XI5/NET35_XI59/XI5/MM7_g
+ N_VSS_XI59/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI5/MM8 N_XI59/XI5/NET35_XI59/XI5/MM8_d N_WL<115>_XI59/XI5/MM8_g
+ N_BLN<10>_XI59/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI5/MM5 N_XI59/XI5/NET34_XI59/XI5/MM5_d N_XI59/XI5/NET33_XI59/XI5/MM5_g
+ N_VDD_XI59/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI5/MM4 N_XI59/XI5/NET33_XI59/XI5/MM4_d N_XI59/XI5/NET34_XI59/XI5/MM4_g
+ N_VDD_XI59/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI5/MM10 N_XI59/XI5/NET35_XI59/XI5/MM10_d N_XI59/XI5/NET36_XI59/XI5/MM10_g
+ N_VDD_XI59/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI5/MM11 N_XI59/XI5/NET36_XI59/XI5/MM11_d N_XI59/XI5/NET35_XI59/XI5/MM11_g
+ N_VDD_XI59/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI6/MM2 N_XI59/XI6/NET34_XI59/XI6/MM2_d N_XI59/XI6/NET33_XI59/XI6/MM2_g
+ N_VSS_XI59/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM3 N_XI59/XI6/NET33_XI59/XI6/MM3_d N_WL<114>_XI59/XI6/MM3_g
+ N_BLN<9>_XI59/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM0 N_XI59/XI6/NET34_XI59/XI6/MM0_d N_WL<114>_XI59/XI6/MM0_g
+ N_BL<9>_XI59/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM1 N_XI59/XI6/NET33_XI59/XI6/MM1_d N_XI59/XI6/NET34_XI59/XI6/MM1_g
+ N_VSS_XI59/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM9 N_XI59/XI6/NET36_XI59/XI6/MM9_d N_WL<115>_XI59/XI6/MM9_g
+ N_BL<9>_XI59/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM6 N_XI59/XI6/NET35_XI59/XI6/MM6_d N_XI59/XI6/NET36_XI59/XI6/MM6_g
+ N_VSS_XI59/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM7 N_XI59/XI6/NET36_XI59/XI6/MM7_d N_XI59/XI6/NET35_XI59/XI6/MM7_g
+ N_VSS_XI59/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM8 N_XI59/XI6/NET35_XI59/XI6/MM8_d N_WL<115>_XI59/XI6/MM8_g
+ N_BLN<9>_XI59/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI6/MM5 N_XI59/XI6/NET34_XI59/XI6/MM5_d N_XI59/XI6/NET33_XI59/XI6/MM5_g
+ N_VDD_XI59/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI6/MM4 N_XI59/XI6/NET33_XI59/XI6/MM4_d N_XI59/XI6/NET34_XI59/XI6/MM4_g
+ N_VDD_XI59/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI6/MM10 N_XI59/XI6/NET35_XI59/XI6/MM10_d N_XI59/XI6/NET36_XI59/XI6/MM10_g
+ N_VDD_XI59/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI6/MM11 N_XI59/XI6/NET36_XI59/XI6/MM11_d N_XI59/XI6/NET35_XI59/XI6/MM11_g
+ N_VDD_XI59/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI7/MM2 N_XI59/XI7/NET34_XI59/XI7/MM2_d N_XI59/XI7/NET33_XI59/XI7/MM2_g
+ N_VSS_XI59/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM3 N_XI59/XI7/NET33_XI59/XI7/MM3_d N_WL<114>_XI59/XI7/MM3_g
+ N_BLN<8>_XI59/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM0 N_XI59/XI7/NET34_XI59/XI7/MM0_d N_WL<114>_XI59/XI7/MM0_g
+ N_BL<8>_XI59/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM1 N_XI59/XI7/NET33_XI59/XI7/MM1_d N_XI59/XI7/NET34_XI59/XI7/MM1_g
+ N_VSS_XI59/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM9 N_XI59/XI7/NET36_XI59/XI7/MM9_d N_WL<115>_XI59/XI7/MM9_g
+ N_BL<8>_XI59/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM6 N_XI59/XI7/NET35_XI59/XI7/MM6_d N_XI59/XI7/NET36_XI59/XI7/MM6_g
+ N_VSS_XI59/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM7 N_XI59/XI7/NET36_XI59/XI7/MM7_d N_XI59/XI7/NET35_XI59/XI7/MM7_g
+ N_VSS_XI59/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM8 N_XI59/XI7/NET35_XI59/XI7/MM8_d N_WL<115>_XI59/XI7/MM8_g
+ N_BLN<8>_XI59/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI7/MM5 N_XI59/XI7/NET34_XI59/XI7/MM5_d N_XI59/XI7/NET33_XI59/XI7/MM5_g
+ N_VDD_XI59/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI7/MM4 N_XI59/XI7/NET33_XI59/XI7/MM4_d N_XI59/XI7/NET34_XI59/XI7/MM4_g
+ N_VDD_XI59/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI7/MM10 N_XI59/XI7/NET35_XI59/XI7/MM10_d N_XI59/XI7/NET36_XI59/XI7/MM10_g
+ N_VDD_XI59/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI7/MM11 N_XI59/XI7/NET36_XI59/XI7/MM11_d N_XI59/XI7/NET35_XI59/XI7/MM11_g
+ N_VDD_XI59/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI8/MM2 N_XI59/XI8/NET34_XI59/XI8/MM2_d N_XI59/XI8/NET33_XI59/XI8/MM2_g
+ N_VSS_XI59/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM3 N_XI59/XI8/NET33_XI59/XI8/MM3_d N_WL<114>_XI59/XI8/MM3_g
+ N_BLN<7>_XI59/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM0 N_XI59/XI8/NET34_XI59/XI8/MM0_d N_WL<114>_XI59/XI8/MM0_g
+ N_BL<7>_XI59/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM1 N_XI59/XI8/NET33_XI59/XI8/MM1_d N_XI59/XI8/NET34_XI59/XI8/MM1_g
+ N_VSS_XI59/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM9 N_XI59/XI8/NET36_XI59/XI8/MM9_d N_WL<115>_XI59/XI8/MM9_g
+ N_BL<7>_XI59/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM6 N_XI59/XI8/NET35_XI59/XI8/MM6_d N_XI59/XI8/NET36_XI59/XI8/MM6_g
+ N_VSS_XI59/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM7 N_XI59/XI8/NET36_XI59/XI8/MM7_d N_XI59/XI8/NET35_XI59/XI8/MM7_g
+ N_VSS_XI59/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM8 N_XI59/XI8/NET35_XI59/XI8/MM8_d N_WL<115>_XI59/XI8/MM8_g
+ N_BLN<7>_XI59/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI8/MM5 N_XI59/XI8/NET34_XI59/XI8/MM5_d N_XI59/XI8/NET33_XI59/XI8/MM5_g
+ N_VDD_XI59/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI8/MM4 N_XI59/XI8/NET33_XI59/XI8/MM4_d N_XI59/XI8/NET34_XI59/XI8/MM4_g
+ N_VDD_XI59/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI8/MM10 N_XI59/XI8/NET35_XI59/XI8/MM10_d N_XI59/XI8/NET36_XI59/XI8/MM10_g
+ N_VDD_XI59/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI8/MM11 N_XI59/XI8/NET36_XI59/XI8/MM11_d N_XI59/XI8/NET35_XI59/XI8/MM11_g
+ N_VDD_XI59/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI9/MM2 N_XI59/XI9/NET34_XI59/XI9/MM2_d N_XI59/XI9/NET33_XI59/XI9/MM2_g
+ N_VSS_XI59/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM3 N_XI59/XI9/NET33_XI59/XI9/MM3_d N_WL<114>_XI59/XI9/MM3_g
+ N_BLN<6>_XI59/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM0 N_XI59/XI9/NET34_XI59/XI9/MM0_d N_WL<114>_XI59/XI9/MM0_g
+ N_BL<6>_XI59/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM1 N_XI59/XI9/NET33_XI59/XI9/MM1_d N_XI59/XI9/NET34_XI59/XI9/MM1_g
+ N_VSS_XI59/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM9 N_XI59/XI9/NET36_XI59/XI9/MM9_d N_WL<115>_XI59/XI9/MM9_g
+ N_BL<6>_XI59/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM6 N_XI59/XI9/NET35_XI59/XI9/MM6_d N_XI59/XI9/NET36_XI59/XI9/MM6_g
+ N_VSS_XI59/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM7 N_XI59/XI9/NET36_XI59/XI9/MM7_d N_XI59/XI9/NET35_XI59/XI9/MM7_g
+ N_VSS_XI59/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM8 N_XI59/XI9/NET35_XI59/XI9/MM8_d N_WL<115>_XI59/XI9/MM8_g
+ N_BLN<6>_XI59/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI9/MM5 N_XI59/XI9/NET34_XI59/XI9/MM5_d N_XI59/XI9/NET33_XI59/XI9/MM5_g
+ N_VDD_XI59/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI9/MM4 N_XI59/XI9/NET33_XI59/XI9/MM4_d N_XI59/XI9/NET34_XI59/XI9/MM4_g
+ N_VDD_XI59/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI9/MM10 N_XI59/XI9/NET35_XI59/XI9/MM10_d N_XI59/XI9/NET36_XI59/XI9/MM10_g
+ N_VDD_XI59/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI9/MM11 N_XI59/XI9/NET36_XI59/XI9/MM11_d N_XI59/XI9/NET35_XI59/XI9/MM11_g
+ N_VDD_XI59/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI10/MM2 N_XI59/XI10/NET34_XI59/XI10/MM2_d
+ N_XI59/XI10/NET33_XI59/XI10/MM2_g N_VSS_XI59/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI10/MM3 N_XI59/XI10/NET33_XI59/XI10/MM3_d N_WL<114>_XI59/XI10/MM3_g
+ N_BLN<5>_XI59/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI10/MM0 N_XI59/XI10/NET34_XI59/XI10/MM0_d N_WL<114>_XI59/XI10/MM0_g
+ N_BL<5>_XI59/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI10/MM1 N_XI59/XI10/NET33_XI59/XI10/MM1_d
+ N_XI59/XI10/NET34_XI59/XI10/MM1_g N_VSS_XI59/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI10/MM9 N_XI59/XI10/NET36_XI59/XI10/MM9_d N_WL<115>_XI59/XI10/MM9_g
+ N_BL<5>_XI59/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI10/MM6 N_XI59/XI10/NET35_XI59/XI10/MM6_d
+ N_XI59/XI10/NET36_XI59/XI10/MM6_g N_VSS_XI59/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI10/MM7 N_XI59/XI10/NET36_XI59/XI10/MM7_d
+ N_XI59/XI10/NET35_XI59/XI10/MM7_g N_VSS_XI59/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI10/MM8 N_XI59/XI10/NET35_XI59/XI10/MM8_d N_WL<115>_XI59/XI10/MM8_g
+ N_BLN<5>_XI59/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI10/MM5 N_XI59/XI10/NET34_XI59/XI10/MM5_d
+ N_XI59/XI10/NET33_XI59/XI10/MM5_g N_VDD_XI59/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI10/MM4 N_XI59/XI10/NET33_XI59/XI10/MM4_d
+ N_XI59/XI10/NET34_XI59/XI10/MM4_g N_VDD_XI59/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI10/MM10 N_XI59/XI10/NET35_XI59/XI10/MM10_d
+ N_XI59/XI10/NET36_XI59/XI10/MM10_g N_VDD_XI59/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI10/MM11 N_XI59/XI10/NET36_XI59/XI10/MM11_d
+ N_XI59/XI10/NET35_XI59/XI10/MM11_g N_VDD_XI59/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI11/MM2 N_XI59/XI11/NET34_XI59/XI11/MM2_d
+ N_XI59/XI11/NET33_XI59/XI11/MM2_g N_VSS_XI59/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI11/MM3 N_XI59/XI11/NET33_XI59/XI11/MM3_d N_WL<114>_XI59/XI11/MM3_g
+ N_BLN<4>_XI59/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI11/MM0 N_XI59/XI11/NET34_XI59/XI11/MM0_d N_WL<114>_XI59/XI11/MM0_g
+ N_BL<4>_XI59/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI11/MM1 N_XI59/XI11/NET33_XI59/XI11/MM1_d
+ N_XI59/XI11/NET34_XI59/XI11/MM1_g N_VSS_XI59/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI11/MM9 N_XI59/XI11/NET36_XI59/XI11/MM9_d N_WL<115>_XI59/XI11/MM9_g
+ N_BL<4>_XI59/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI11/MM6 N_XI59/XI11/NET35_XI59/XI11/MM6_d
+ N_XI59/XI11/NET36_XI59/XI11/MM6_g N_VSS_XI59/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI11/MM7 N_XI59/XI11/NET36_XI59/XI11/MM7_d
+ N_XI59/XI11/NET35_XI59/XI11/MM7_g N_VSS_XI59/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI11/MM8 N_XI59/XI11/NET35_XI59/XI11/MM8_d N_WL<115>_XI59/XI11/MM8_g
+ N_BLN<4>_XI59/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI11/MM5 N_XI59/XI11/NET34_XI59/XI11/MM5_d
+ N_XI59/XI11/NET33_XI59/XI11/MM5_g N_VDD_XI59/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI11/MM4 N_XI59/XI11/NET33_XI59/XI11/MM4_d
+ N_XI59/XI11/NET34_XI59/XI11/MM4_g N_VDD_XI59/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI11/MM10 N_XI59/XI11/NET35_XI59/XI11/MM10_d
+ N_XI59/XI11/NET36_XI59/XI11/MM10_g N_VDD_XI59/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI11/MM11 N_XI59/XI11/NET36_XI59/XI11/MM11_d
+ N_XI59/XI11/NET35_XI59/XI11/MM11_g N_VDD_XI59/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI12/MM2 N_XI59/XI12/NET34_XI59/XI12/MM2_d
+ N_XI59/XI12/NET33_XI59/XI12/MM2_g N_VSS_XI59/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI12/MM3 N_XI59/XI12/NET33_XI59/XI12/MM3_d N_WL<114>_XI59/XI12/MM3_g
+ N_BLN<3>_XI59/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI12/MM0 N_XI59/XI12/NET34_XI59/XI12/MM0_d N_WL<114>_XI59/XI12/MM0_g
+ N_BL<3>_XI59/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI12/MM1 N_XI59/XI12/NET33_XI59/XI12/MM1_d
+ N_XI59/XI12/NET34_XI59/XI12/MM1_g N_VSS_XI59/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI12/MM9 N_XI59/XI12/NET36_XI59/XI12/MM9_d N_WL<115>_XI59/XI12/MM9_g
+ N_BL<3>_XI59/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI12/MM6 N_XI59/XI12/NET35_XI59/XI12/MM6_d
+ N_XI59/XI12/NET36_XI59/XI12/MM6_g N_VSS_XI59/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI12/MM7 N_XI59/XI12/NET36_XI59/XI12/MM7_d
+ N_XI59/XI12/NET35_XI59/XI12/MM7_g N_VSS_XI59/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI12/MM8 N_XI59/XI12/NET35_XI59/XI12/MM8_d N_WL<115>_XI59/XI12/MM8_g
+ N_BLN<3>_XI59/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI12/MM5 N_XI59/XI12/NET34_XI59/XI12/MM5_d
+ N_XI59/XI12/NET33_XI59/XI12/MM5_g N_VDD_XI59/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI12/MM4 N_XI59/XI12/NET33_XI59/XI12/MM4_d
+ N_XI59/XI12/NET34_XI59/XI12/MM4_g N_VDD_XI59/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI12/MM10 N_XI59/XI12/NET35_XI59/XI12/MM10_d
+ N_XI59/XI12/NET36_XI59/XI12/MM10_g N_VDD_XI59/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI12/MM11 N_XI59/XI12/NET36_XI59/XI12/MM11_d
+ N_XI59/XI12/NET35_XI59/XI12/MM11_g N_VDD_XI59/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI13/MM2 N_XI59/XI13/NET34_XI59/XI13/MM2_d
+ N_XI59/XI13/NET33_XI59/XI13/MM2_g N_VSS_XI59/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI13/MM3 N_XI59/XI13/NET33_XI59/XI13/MM3_d N_WL<114>_XI59/XI13/MM3_g
+ N_BLN<2>_XI59/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI13/MM0 N_XI59/XI13/NET34_XI59/XI13/MM0_d N_WL<114>_XI59/XI13/MM0_g
+ N_BL<2>_XI59/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI13/MM1 N_XI59/XI13/NET33_XI59/XI13/MM1_d
+ N_XI59/XI13/NET34_XI59/XI13/MM1_g N_VSS_XI59/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI13/MM9 N_XI59/XI13/NET36_XI59/XI13/MM9_d N_WL<115>_XI59/XI13/MM9_g
+ N_BL<2>_XI59/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI13/MM6 N_XI59/XI13/NET35_XI59/XI13/MM6_d
+ N_XI59/XI13/NET36_XI59/XI13/MM6_g N_VSS_XI59/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI13/MM7 N_XI59/XI13/NET36_XI59/XI13/MM7_d
+ N_XI59/XI13/NET35_XI59/XI13/MM7_g N_VSS_XI59/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI13/MM8 N_XI59/XI13/NET35_XI59/XI13/MM8_d N_WL<115>_XI59/XI13/MM8_g
+ N_BLN<2>_XI59/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI13/MM5 N_XI59/XI13/NET34_XI59/XI13/MM5_d
+ N_XI59/XI13/NET33_XI59/XI13/MM5_g N_VDD_XI59/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI13/MM4 N_XI59/XI13/NET33_XI59/XI13/MM4_d
+ N_XI59/XI13/NET34_XI59/XI13/MM4_g N_VDD_XI59/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI13/MM10 N_XI59/XI13/NET35_XI59/XI13/MM10_d
+ N_XI59/XI13/NET36_XI59/XI13/MM10_g N_VDD_XI59/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI13/MM11 N_XI59/XI13/NET36_XI59/XI13/MM11_d
+ N_XI59/XI13/NET35_XI59/XI13/MM11_g N_VDD_XI59/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI14/MM2 N_XI59/XI14/NET34_XI59/XI14/MM2_d
+ N_XI59/XI14/NET33_XI59/XI14/MM2_g N_VSS_XI59/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI14/MM3 N_XI59/XI14/NET33_XI59/XI14/MM3_d N_WL<114>_XI59/XI14/MM3_g
+ N_BLN<1>_XI59/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI14/MM0 N_XI59/XI14/NET34_XI59/XI14/MM0_d N_WL<114>_XI59/XI14/MM0_g
+ N_BL<1>_XI59/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI14/MM1 N_XI59/XI14/NET33_XI59/XI14/MM1_d
+ N_XI59/XI14/NET34_XI59/XI14/MM1_g N_VSS_XI59/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI14/MM9 N_XI59/XI14/NET36_XI59/XI14/MM9_d N_WL<115>_XI59/XI14/MM9_g
+ N_BL<1>_XI59/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI14/MM6 N_XI59/XI14/NET35_XI59/XI14/MM6_d
+ N_XI59/XI14/NET36_XI59/XI14/MM6_g N_VSS_XI59/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI14/MM7 N_XI59/XI14/NET36_XI59/XI14/MM7_d
+ N_XI59/XI14/NET35_XI59/XI14/MM7_g N_VSS_XI59/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI14/MM8 N_XI59/XI14/NET35_XI59/XI14/MM8_d N_WL<115>_XI59/XI14/MM8_g
+ N_BLN<1>_XI59/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI14/MM5 N_XI59/XI14/NET34_XI59/XI14/MM5_d
+ N_XI59/XI14/NET33_XI59/XI14/MM5_g N_VDD_XI59/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI14/MM4 N_XI59/XI14/NET33_XI59/XI14/MM4_d
+ N_XI59/XI14/NET34_XI59/XI14/MM4_g N_VDD_XI59/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI14/MM10 N_XI59/XI14/NET35_XI59/XI14/MM10_d
+ N_XI59/XI14/NET36_XI59/XI14/MM10_g N_VDD_XI59/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI14/MM11 N_XI59/XI14/NET36_XI59/XI14/MM11_d
+ N_XI59/XI14/NET35_XI59/XI14/MM11_g N_VDD_XI59/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI15/MM2 N_XI59/XI15/NET34_XI59/XI15/MM2_d
+ N_XI59/XI15/NET33_XI59/XI15/MM2_g N_VSS_XI59/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI15/MM3 N_XI59/XI15/NET33_XI59/XI15/MM3_d N_WL<114>_XI59/XI15/MM3_g
+ N_BLN<0>_XI59/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI15/MM0 N_XI59/XI15/NET34_XI59/XI15/MM0_d N_WL<114>_XI59/XI15/MM0_g
+ N_BL<0>_XI59/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI15/MM1 N_XI59/XI15/NET33_XI59/XI15/MM1_d
+ N_XI59/XI15/NET34_XI59/XI15/MM1_g N_VSS_XI59/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI15/MM9 N_XI59/XI15/NET36_XI59/XI15/MM9_d N_WL<115>_XI59/XI15/MM9_g
+ N_BL<0>_XI59/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI15/MM6 N_XI59/XI15/NET35_XI59/XI15/MM6_d
+ N_XI59/XI15/NET36_XI59/XI15/MM6_g N_VSS_XI59/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI15/MM7 N_XI59/XI15/NET36_XI59/XI15/MM7_d
+ N_XI59/XI15/NET35_XI59/XI15/MM7_g N_VSS_XI59/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI59/XI15/MM8 N_XI59/XI15/NET35_XI59/XI15/MM8_d N_WL<115>_XI59/XI15/MM8_g
+ N_BLN<0>_XI59/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI59/XI15/MM5 N_XI59/XI15/NET34_XI59/XI15/MM5_d
+ N_XI59/XI15/NET33_XI59/XI15/MM5_g N_VDD_XI59/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI15/MM4 N_XI59/XI15/NET33_XI59/XI15/MM4_d
+ N_XI59/XI15/NET34_XI59/XI15/MM4_g N_VDD_XI59/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI15/MM10 N_XI59/XI15/NET35_XI59/XI15/MM10_d
+ N_XI59/XI15/NET36_XI59/XI15/MM10_g N_VDD_XI59/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI59/XI15/MM11 N_XI59/XI15/NET36_XI59/XI15/MM11_d
+ N_XI59/XI15/NET35_XI59/XI15/MM11_g N_VDD_XI59/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI0/MM2 N_XI60/XI0/NET34_XI60/XI0/MM2_d N_XI60/XI0/NET33_XI60/XI0/MM2_g
+ N_VSS_XI60/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI0/MM3 N_XI60/XI0/NET33_XI60/XI0/MM3_d N_WL<116>_XI60/XI0/MM3_g
+ N_BLN<15>_XI60/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI0/MM0 N_XI60/XI0/NET34_XI60/XI0/MM0_d N_WL<116>_XI60/XI0/MM0_g
+ N_BL<15>_XI60/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI0/MM1 N_XI60/XI0/NET33_XI60/XI0/MM1_d N_XI60/XI0/NET34_XI60/XI0/MM1_g
+ N_VSS_XI60/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI0/MM9 N_XI60/XI0/NET36_XI60/XI0/MM9_d N_WL<117>_XI60/XI0/MM9_g
+ N_BL<15>_XI60/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI0/MM6 N_XI60/XI0/NET35_XI60/XI0/MM6_d N_XI60/XI0/NET36_XI60/XI0/MM6_g
+ N_VSS_XI60/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI0/MM7 N_XI60/XI0/NET36_XI60/XI0/MM7_d N_XI60/XI0/NET35_XI60/XI0/MM7_g
+ N_VSS_XI60/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI0/MM8 N_XI60/XI0/NET35_XI60/XI0/MM8_d N_WL<117>_XI60/XI0/MM8_g
+ N_BLN<15>_XI60/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI0/MM5 N_XI60/XI0/NET34_XI60/XI0/MM5_d N_XI60/XI0/NET33_XI60/XI0/MM5_g
+ N_VDD_XI60/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI0/MM4 N_XI60/XI0/NET33_XI60/XI0/MM4_d N_XI60/XI0/NET34_XI60/XI0/MM4_g
+ N_VDD_XI60/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI0/MM10 N_XI60/XI0/NET35_XI60/XI0/MM10_d N_XI60/XI0/NET36_XI60/XI0/MM10_g
+ N_VDD_XI60/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI0/MM11 N_XI60/XI0/NET36_XI60/XI0/MM11_d N_XI60/XI0/NET35_XI60/XI0/MM11_g
+ N_VDD_XI60/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI1/MM2 N_XI60/XI1/NET34_XI60/XI1/MM2_d N_XI60/XI1/NET33_XI60/XI1/MM2_g
+ N_VSS_XI60/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI1/MM3 N_XI60/XI1/NET33_XI60/XI1/MM3_d N_WL<116>_XI60/XI1/MM3_g
+ N_BLN<14>_XI60/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI1/MM0 N_XI60/XI1/NET34_XI60/XI1/MM0_d N_WL<116>_XI60/XI1/MM0_g
+ N_BL<14>_XI60/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI1/MM1 N_XI60/XI1/NET33_XI60/XI1/MM1_d N_XI60/XI1/NET34_XI60/XI1/MM1_g
+ N_VSS_XI60/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI1/MM9 N_XI60/XI1/NET36_XI60/XI1/MM9_d N_WL<117>_XI60/XI1/MM9_g
+ N_BL<14>_XI60/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI1/MM6 N_XI60/XI1/NET35_XI60/XI1/MM6_d N_XI60/XI1/NET36_XI60/XI1/MM6_g
+ N_VSS_XI60/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI1/MM7 N_XI60/XI1/NET36_XI60/XI1/MM7_d N_XI60/XI1/NET35_XI60/XI1/MM7_g
+ N_VSS_XI60/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI1/MM8 N_XI60/XI1/NET35_XI60/XI1/MM8_d N_WL<117>_XI60/XI1/MM8_g
+ N_BLN<14>_XI60/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI1/MM5 N_XI60/XI1/NET34_XI60/XI1/MM5_d N_XI60/XI1/NET33_XI60/XI1/MM5_g
+ N_VDD_XI60/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI1/MM4 N_XI60/XI1/NET33_XI60/XI1/MM4_d N_XI60/XI1/NET34_XI60/XI1/MM4_g
+ N_VDD_XI60/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI1/MM10 N_XI60/XI1/NET35_XI60/XI1/MM10_d N_XI60/XI1/NET36_XI60/XI1/MM10_g
+ N_VDD_XI60/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI1/MM11 N_XI60/XI1/NET36_XI60/XI1/MM11_d N_XI60/XI1/NET35_XI60/XI1/MM11_g
+ N_VDD_XI60/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI2/MM2 N_XI60/XI2/NET34_XI60/XI2/MM2_d N_XI60/XI2/NET33_XI60/XI2/MM2_g
+ N_VSS_XI60/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI2/MM3 N_XI60/XI2/NET33_XI60/XI2/MM3_d N_WL<116>_XI60/XI2/MM3_g
+ N_BLN<13>_XI60/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI2/MM0 N_XI60/XI2/NET34_XI60/XI2/MM0_d N_WL<116>_XI60/XI2/MM0_g
+ N_BL<13>_XI60/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI2/MM1 N_XI60/XI2/NET33_XI60/XI2/MM1_d N_XI60/XI2/NET34_XI60/XI2/MM1_g
+ N_VSS_XI60/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI2/MM9 N_XI60/XI2/NET36_XI60/XI2/MM9_d N_WL<117>_XI60/XI2/MM9_g
+ N_BL<13>_XI60/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI2/MM6 N_XI60/XI2/NET35_XI60/XI2/MM6_d N_XI60/XI2/NET36_XI60/XI2/MM6_g
+ N_VSS_XI60/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI2/MM7 N_XI60/XI2/NET36_XI60/XI2/MM7_d N_XI60/XI2/NET35_XI60/XI2/MM7_g
+ N_VSS_XI60/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI2/MM8 N_XI60/XI2/NET35_XI60/XI2/MM8_d N_WL<117>_XI60/XI2/MM8_g
+ N_BLN<13>_XI60/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI2/MM5 N_XI60/XI2/NET34_XI60/XI2/MM5_d N_XI60/XI2/NET33_XI60/XI2/MM5_g
+ N_VDD_XI60/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI2/MM4 N_XI60/XI2/NET33_XI60/XI2/MM4_d N_XI60/XI2/NET34_XI60/XI2/MM4_g
+ N_VDD_XI60/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI2/MM10 N_XI60/XI2/NET35_XI60/XI2/MM10_d N_XI60/XI2/NET36_XI60/XI2/MM10_g
+ N_VDD_XI60/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI2/MM11 N_XI60/XI2/NET36_XI60/XI2/MM11_d N_XI60/XI2/NET35_XI60/XI2/MM11_g
+ N_VDD_XI60/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI3/MM2 N_XI60/XI3/NET34_XI60/XI3/MM2_d N_XI60/XI3/NET33_XI60/XI3/MM2_g
+ N_VSS_XI60/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI3/MM3 N_XI60/XI3/NET33_XI60/XI3/MM3_d N_WL<116>_XI60/XI3/MM3_g
+ N_BLN<12>_XI60/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI3/MM0 N_XI60/XI3/NET34_XI60/XI3/MM0_d N_WL<116>_XI60/XI3/MM0_g
+ N_BL<12>_XI60/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI3/MM1 N_XI60/XI3/NET33_XI60/XI3/MM1_d N_XI60/XI3/NET34_XI60/XI3/MM1_g
+ N_VSS_XI60/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI3/MM9 N_XI60/XI3/NET36_XI60/XI3/MM9_d N_WL<117>_XI60/XI3/MM9_g
+ N_BL<12>_XI60/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI3/MM6 N_XI60/XI3/NET35_XI60/XI3/MM6_d N_XI60/XI3/NET36_XI60/XI3/MM6_g
+ N_VSS_XI60/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI3/MM7 N_XI60/XI3/NET36_XI60/XI3/MM7_d N_XI60/XI3/NET35_XI60/XI3/MM7_g
+ N_VSS_XI60/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI3/MM8 N_XI60/XI3/NET35_XI60/XI3/MM8_d N_WL<117>_XI60/XI3/MM8_g
+ N_BLN<12>_XI60/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI3/MM5 N_XI60/XI3/NET34_XI60/XI3/MM5_d N_XI60/XI3/NET33_XI60/XI3/MM5_g
+ N_VDD_XI60/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI3/MM4 N_XI60/XI3/NET33_XI60/XI3/MM4_d N_XI60/XI3/NET34_XI60/XI3/MM4_g
+ N_VDD_XI60/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI3/MM10 N_XI60/XI3/NET35_XI60/XI3/MM10_d N_XI60/XI3/NET36_XI60/XI3/MM10_g
+ N_VDD_XI60/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI3/MM11 N_XI60/XI3/NET36_XI60/XI3/MM11_d N_XI60/XI3/NET35_XI60/XI3/MM11_g
+ N_VDD_XI60/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI4/MM2 N_XI60/XI4/NET34_XI60/XI4/MM2_d N_XI60/XI4/NET33_XI60/XI4/MM2_g
+ N_VSS_XI60/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI4/MM3 N_XI60/XI4/NET33_XI60/XI4/MM3_d N_WL<116>_XI60/XI4/MM3_g
+ N_BLN<11>_XI60/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI4/MM0 N_XI60/XI4/NET34_XI60/XI4/MM0_d N_WL<116>_XI60/XI4/MM0_g
+ N_BL<11>_XI60/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI4/MM1 N_XI60/XI4/NET33_XI60/XI4/MM1_d N_XI60/XI4/NET34_XI60/XI4/MM1_g
+ N_VSS_XI60/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI4/MM9 N_XI60/XI4/NET36_XI60/XI4/MM9_d N_WL<117>_XI60/XI4/MM9_g
+ N_BL<11>_XI60/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI4/MM6 N_XI60/XI4/NET35_XI60/XI4/MM6_d N_XI60/XI4/NET36_XI60/XI4/MM6_g
+ N_VSS_XI60/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI4/MM7 N_XI60/XI4/NET36_XI60/XI4/MM7_d N_XI60/XI4/NET35_XI60/XI4/MM7_g
+ N_VSS_XI60/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI4/MM8 N_XI60/XI4/NET35_XI60/XI4/MM8_d N_WL<117>_XI60/XI4/MM8_g
+ N_BLN<11>_XI60/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI4/MM5 N_XI60/XI4/NET34_XI60/XI4/MM5_d N_XI60/XI4/NET33_XI60/XI4/MM5_g
+ N_VDD_XI60/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI4/MM4 N_XI60/XI4/NET33_XI60/XI4/MM4_d N_XI60/XI4/NET34_XI60/XI4/MM4_g
+ N_VDD_XI60/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI4/MM10 N_XI60/XI4/NET35_XI60/XI4/MM10_d N_XI60/XI4/NET36_XI60/XI4/MM10_g
+ N_VDD_XI60/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI4/MM11 N_XI60/XI4/NET36_XI60/XI4/MM11_d N_XI60/XI4/NET35_XI60/XI4/MM11_g
+ N_VDD_XI60/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI5/MM2 N_XI60/XI5/NET34_XI60/XI5/MM2_d N_XI60/XI5/NET33_XI60/XI5/MM2_g
+ N_VSS_XI60/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI5/MM3 N_XI60/XI5/NET33_XI60/XI5/MM3_d N_WL<116>_XI60/XI5/MM3_g
+ N_BLN<10>_XI60/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI5/MM0 N_XI60/XI5/NET34_XI60/XI5/MM0_d N_WL<116>_XI60/XI5/MM0_g
+ N_BL<10>_XI60/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI5/MM1 N_XI60/XI5/NET33_XI60/XI5/MM1_d N_XI60/XI5/NET34_XI60/XI5/MM1_g
+ N_VSS_XI60/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI5/MM9 N_XI60/XI5/NET36_XI60/XI5/MM9_d N_WL<117>_XI60/XI5/MM9_g
+ N_BL<10>_XI60/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI5/MM6 N_XI60/XI5/NET35_XI60/XI5/MM6_d N_XI60/XI5/NET36_XI60/XI5/MM6_g
+ N_VSS_XI60/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI5/MM7 N_XI60/XI5/NET36_XI60/XI5/MM7_d N_XI60/XI5/NET35_XI60/XI5/MM7_g
+ N_VSS_XI60/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI5/MM8 N_XI60/XI5/NET35_XI60/XI5/MM8_d N_WL<117>_XI60/XI5/MM8_g
+ N_BLN<10>_XI60/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI5/MM5 N_XI60/XI5/NET34_XI60/XI5/MM5_d N_XI60/XI5/NET33_XI60/XI5/MM5_g
+ N_VDD_XI60/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI5/MM4 N_XI60/XI5/NET33_XI60/XI5/MM4_d N_XI60/XI5/NET34_XI60/XI5/MM4_g
+ N_VDD_XI60/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI5/MM10 N_XI60/XI5/NET35_XI60/XI5/MM10_d N_XI60/XI5/NET36_XI60/XI5/MM10_g
+ N_VDD_XI60/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI5/MM11 N_XI60/XI5/NET36_XI60/XI5/MM11_d N_XI60/XI5/NET35_XI60/XI5/MM11_g
+ N_VDD_XI60/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI6/MM2 N_XI60/XI6/NET34_XI60/XI6/MM2_d N_XI60/XI6/NET33_XI60/XI6/MM2_g
+ N_VSS_XI60/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM3 N_XI60/XI6/NET33_XI60/XI6/MM3_d N_WL<116>_XI60/XI6/MM3_g
+ N_BLN<9>_XI60/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM0 N_XI60/XI6/NET34_XI60/XI6/MM0_d N_WL<116>_XI60/XI6/MM0_g
+ N_BL<9>_XI60/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM1 N_XI60/XI6/NET33_XI60/XI6/MM1_d N_XI60/XI6/NET34_XI60/XI6/MM1_g
+ N_VSS_XI60/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM9 N_XI60/XI6/NET36_XI60/XI6/MM9_d N_WL<117>_XI60/XI6/MM9_g
+ N_BL<9>_XI60/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM6 N_XI60/XI6/NET35_XI60/XI6/MM6_d N_XI60/XI6/NET36_XI60/XI6/MM6_g
+ N_VSS_XI60/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM7 N_XI60/XI6/NET36_XI60/XI6/MM7_d N_XI60/XI6/NET35_XI60/XI6/MM7_g
+ N_VSS_XI60/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM8 N_XI60/XI6/NET35_XI60/XI6/MM8_d N_WL<117>_XI60/XI6/MM8_g
+ N_BLN<9>_XI60/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI6/MM5 N_XI60/XI6/NET34_XI60/XI6/MM5_d N_XI60/XI6/NET33_XI60/XI6/MM5_g
+ N_VDD_XI60/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI6/MM4 N_XI60/XI6/NET33_XI60/XI6/MM4_d N_XI60/XI6/NET34_XI60/XI6/MM4_g
+ N_VDD_XI60/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI6/MM10 N_XI60/XI6/NET35_XI60/XI6/MM10_d N_XI60/XI6/NET36_XI60/XI6/MM10_g
+ N_VDD_XI60/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI6/MM11 N_XI60/XI6/NET36_XI60/XI6/MM11_d N_XI60/XI6/NET35_XI60/XI6/MM11_g
+ N_VDD_XI60/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI7/MM2 N_XI60/XI7/NET34_XI60/XI7/MM2_d N_XI60/XI7/NET33_XI60/XI7/MM2_g
+ N_VSS_XI60/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM3 N_XI60/XI7/NET33_XI60/XI7/MM3_d N_WL<116>_XI60/XI7/MM3_g
+ N_BLN<8>_XI60/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM0 N_XI60/XI7/NET34_XI60/XI7/MM0_d N_WL<116>_XI60/XI7/MM0_g
+ N_BL<8>_XI60/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM1 N_XI60/XI7/NET33_XI60/XI7/MM1_d N_XI60/XI7/NET34_XI60/XI7/MM1_g
+ N_VSS_XI60/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM9 N_XI60/XI7/NET36_XI60/XI7/MM9_d N_WL<117>_XI60/XI7/MM9_g
+ N_BL<8>_XI60/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM6 N_XI60/XI7/NET35_XI60/XI7/MM6_d N_XI60/XI7/NET36_XI60/XI7/MM6_g
+ N_VSS_XI60/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM7 N_XI60/XI7/NET36_XI60/XI7/MM7_d N_XI60/XI7/NET35_XI60/XI7/MM7_g
+ N_VSS_XI60/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM8 N_XI60/XI7/NET35_XI60/XI7/MM8_d N_WL<117>_XI60/XI7/MM8_g
+ N_BLN<8>_XI60/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI7/MM5 N_XI60/XI7/NET34_XI60/XI7/MM5_d N_XI60/XI7/NET33_XI60/XI7/MM5_g
+ N_VDD_XI60/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI7/MM4 N_XI60/XI7/NET33_XI60/XI7/MM4_d N_XI60/XI7/NET34_XI60/XI7/MM4_g
+ N_VDD_XI60/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI7/MM10 N_XI60/XI7/NET35_XI60/XI7/MM10_d N_XI60/XI7/NET36_XI60/XI7/MM10_g
+ N_VDD_XI60/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI7/MM11 N_XI60/XI7/NET36_XI60/XI7/MM11_d N_XI60/XI7/NET35_XI60/XI7/MM11_g
+ N_VDD_XI60/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI8/MM2 N_XI60/XI8/NET34_XI60/XI8/MM2_d N_XI60/XI8/NET33_XI60/XI8/MM2_g
+ N_VSS_XI60/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM3 N_XI60/XI8/NET33_XI60/XI8/MM3_d N_WL<116>_XI60/XI8/MM3_g
+ N_BLN<7>_XI60/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM0 N_XI60/XI8/NET34_XI60/XI8/MM0_d N_WL<116>_XI60/XI8/MM0_g
+ N_BL<7>_XI60/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM1 N_XI60/XI8/NET33_XI60/XI8/MM1_d N_XI60/XI8/NET34_XI60/XI8/MM1_g
+ N_VSS_XI60/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM9 N_XI60/XI8/NET36_XI60/XI8/MM9_d N_WL<117>_XI60/XI8/MM9_g
+ N_BL<7>_XI60/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM6 N_XI60/XI8/NET35_XI60/XI8/MM6_d N_XI60/XI8/NET36_XI60/XI8/MM6_g
+ N_VSS_XI60/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM7 N_XI60/XI8/NET36_XI60/XI8/MM7_d N_XI60/XI8/NET35_XI60/XI8/MM7_g
+ N_VSS_XI60/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM8 N_XI60/XI8/NET35_XI60/XI8/MM8_d N_WL<117>_XI60/XI8/MM8_g
+ N_BLN<7>_XI60/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI8/MM5 N_XI60/XI8/NET34_XI60/XI8/MM5_d N_XI60/XI8/NET33_XI60/XI8/MM5_g
+ N_VDD_XI60/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI8/MM4 N_XI60/XI8/NET33_XI60/XI8/MM4_d N_XI60/XI8/NET34_XI60/XI8/MM4_g
+ N_VDD_XI60/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI8/MM10 N_XI60/XI8/NET35_XI60/XI8/MM10_d N_XI60/XI8/NET36_XI60/XI8/MM10_g
+ N_VDD_XI60/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI8/MM11 N_XI60/XI8/NET36_XI60/XI8/MM11_d N_XI60/XI8/NET35_XI60/XI8/MM11_g
+ N_VDD_XI60/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI9/MM2 N_XI60/XI9/NET34_XI60/XI9/MM2_d N_XI60/XI9/NET33_XI60/XI9/MM2_g
+ N_VSS_XI60/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM3 N_XI60/XI9/NET33_XI60/XI9/MM3_d N_WL<116>_XI60/XI9/MM3_g
+ N_BLN<6>_XI60/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM0 N_XI60/XI9/NET34_XI60/XI9/MM0_d N_WL<116>_XI60/XI9/MM0_g
+ N_BL<6>_XI60/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM1 N_XI60/XI9/NET33_XI60/XI9/MM1_d N_XI60/XI9/NET34_XI60/XI9/MM1_g
+ N_VSS_XI60/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM9 N_XI60/XI9/NET36_XI60/XI9/MM9_d N_WL<117>_XI60/XI9/MM9_g
+ N_BL<6>_XI60/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM6 N_XI60/XI9/NET35_XI60/XI9/MM6_d N_XI60/XI9/NET36_XI60/XI9/MM6_g
+ N_VSS_XI60/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM7 N_XI60/XI9/NET36_XI60/XI9/MM7_d N_XI60/XI9/NET35_XI60/XI9/MM7_g
+ N_VSS_XI60/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM8 N_XI60/XI9/NET35_XI60/XI9/MM8_d N_WL<117>_XI60/XI9/MM8_g
+ N_BLN<6>_XI60/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI9/MM5 N_XI60/XI9/NET34_XI60/XI9/MM5_d N_XI60/XI9/NET33_XI60/XI9/MM5_g
+ N_VDD_XI60/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI9/MM4 N_XI60/XI9/NET33_XI60/XI9/MM4_d N_XI60/XI9/NET34_XI60/XI9/MM4_g
+ N_VDD_XI60/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI9/MM10 N_XI60/XI9/NET35_XI60/XI9/MM10_d N_XI60/XI9/NET36_XI60/XI9/MM10_g
+ N_VDD_XI60/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI9/MM11 N_XI60/XI9/NET36_XI60/XI9/MM11_d N_XI60/XI9/NET35_XI60/XI9/MM11_g
+ N_VDD_XI60/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI10/MM2 N_XI60/XI10/NET34_XI60/XI10/MM2_d
+ N_XI60/XI10/NET33_XI60/XI10/MM2_g N_VSS_XI60/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI10/MM3 N_XI60/XI10/NET33_XI60/XI10/MM3_d N_WL<116>_XI60/XI10/MM3_g
+ N_BLN<5>_XI60/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI10/MM0 N_XI60/XI10/NET34_XI60/XI10/MM0_d N_WL<116>_XI60/XI10/MM0_g
+ N_BL<5>_XI60/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI10/MM1 N_XI60/XI10/NET33_XI60/XI10/MM1_d
+ N_XI60/XI10/NET34_XI60/XI10/MM1_g N_VSS_XI60/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI10/MM9 N_XI60/XI10/NET36_XI60/XI10/MM9_d N_WL<117>_XI60/XI10/MM9_g
+ N_BL<5>_XI60/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI10/MM6 N_XI60/XI10/NET35_XI60/XI10/MM6_d
+ N_XI60/XI10/NET36_XI60/XI10/MM6_g N_VSS_XI60/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI10/MM7 N_XI60/XI10/NET36_XI60/XI10/MM7_d
+ N_XI60/XI10/NET35_XI60/XI10/MM7_g N_VSS_XI60/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI10/MM8 N_XI60/XI10/NET35_XI60/XI10/MM8_d N_WL<117>_XI60/XI10/MM8_g
+ N_BLN<5>_XI60/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI10/MM5 N_XI60/XI10/NET34_XI60/XI10/MM5_d
+ N_XI60/XI10/NET33_XI60/XI10/MM5_g N_VDD_XI60/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI10/MM4 N_XI60/XI10/NET33_XI60/XI10/MM4_d
+ N_XI60/XI10/NET34_XI60/XI10/MM4_g N_VDD_XI60/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI10/MM10 N_XI60/XI10/NET35_XI60/XI10/MM10_d
+ N_XI60/XI10/NET36_XI60/XI10/MM10_g N_VDD_XI60/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI10/MM11 N_XI60/XI10/NET36_XI60/XI10/MM11_d
+ N_XI60/XI10/NET35_XI60/XI10/MM11_g N_VDD_XI60/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI11/MM2 N_XI60/XI11/NET34_XI60/XI11/MM2_d
+ N_XI60/XI11/NET33_XI60/XI11/MM2_g N_VSS_XI60/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI11/MM3 N_XI60/XI11/NET33_XI60/XI11/MM3_d N_WL<116>_XI60/XI11/MM3_g
+ N_BLN<4>_XI60/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI11/MM0 N_XI60/XI11/NET34_XI60/XI11/MM0_d N_WL<116>_XI60/XI11/MM0_g
+ N_BL<4>_XI60/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI11/MM1 N_XI60/XI11/NET33_XI60/XI11/MM1_d
+ N_XI60/XI11/NET34_XI60/XI11/MM1_g N_VSS_XI60/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI11/MM9 N_XI60/XI11/NET36_XI60/XI11/MM9_d N_WL<117>_XI60/XI11/MM9_g
+ N_BL<4>_XI60/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI11/MM6 N_XI60/XI11/NET35_XI60/XI11/MM6_d
+ N_XI60/XI11/NET36_XI60/XI11/MM6_g N_VSS_XI60/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI11/MM7 N_XI60/XI11/NET36_XI60/XI11/MM7_d
+ N_XI60/XI11/NET35_XI60/XI11/MM7_g N_VSS_XI60/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI11/MM8 N_XI60/XI11/NET35_XI60/XI11/MM8_d N_WL<117>_XI60/XI11/MM8_g
+ N_BLN<4>_XI60/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI11/MM5 N_XI60/XI11/NET34_XI60/XI11/MM5_d
+ N_XI60/XI11/NET33_XI60/XI11/MM5_g N_VDD_XI60/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI11/MM4 N_XI60/XI11/NET33_XI60/XI11/MM4_d
+ N_XI60/XI11/NET34_XI60/XI11/MM4_g N_VDD_XI60/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI11/MM10 N_XI60/XI11/NET35_XI60/XI11/MM10_d
+ N_XI60/XI11/NET36_XI60/XI11/MM10_g N_VDD_XI60/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI11/MM11 N_XI60/XI11/NET36_XI60/XI11/MM11_d
+ N_XI60/XI11/NET35_XI60/XI11/MM11_g N_VDD_XI60/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI12/MM2 N_XI60/XI12/NET34_XI60/XI12/MM2_d
+ N_XI60/XI12/NET33_XI60/XI12/MM2_g N_VSS_XI60/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI12/MM3 N_XI60/XI12/NET33_XI60/XI12/MM3_d N_WL<116>_XI60/XI12/MM3_g
+ N_BLN<3>_XI60/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI12/MM0 N_XI60/XI12/NET34_XI60/XI12/MM0_d N_WL<116>_XI60/XI12/MM0_g
+ N_BL<3>_XI60/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI12/MM1 N_XI60/XI12/NET33_XI60/XI12/MM1_d
+ N_XI60/XI12/NET34_XI60/XI12/MM1_g N_VSS_XI60/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI12/MM9 N_XI60/XI12/NET36_XI60/XI12/MM9_d N_WL<117>_XI60/XI12/MM9_g
+ N_BL<3>_XI60/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI12/MM6 N_XI60/XI12/NET35_XI60/XI12/MM6_d
+ N_XI60/XI12/NET36_XI60/XI12/MM6_g N_VSS_XI60/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI12/MM7 N_XI60/XI12/NET36_XI60/XI12/MM7_d
+ N_XI60/XI12/NET35_XI60/XI12/MM7_g N_VSS_XI60/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI12/MM8 N_XI60/XI12/NET35_XI60/XI12/MM8_d N_WL<117>_XI60/XI12/MM8_g
+ N_BLN<3>_XI60/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI12/MM5 N_XI60/XI12/NET34_XI60/XI12/MM5_d
+ N_XI60/XI12/NET33_XI60/XI12/MM5_g N_VDD_XI60/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI12/MM4 N_XI60/XI12/NET33_XI60/XI12/MM4_d
+ N_XI60/XI12/NET34_XI60/XI12/MM4_g N_VDD_XI60/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI12/MM10 N_XI60/XI12/NET35_XI60/XI12/MM10_d
+ N_XI60/XI12/NET36_XI60/XI12/MM10_g N_VDD_XI60/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI12/MM11 N_XI60/XI12/NET36_XI60/XI12/MM11_d
+ N_XI60/XI12/NET35_XI60/XI12/MM11_g N_VDD_XI60/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI13/MM2 N_XI60/XI13/NET34_XI60/XI13/MM2_d
+ N_XI60/XI13/NET33_XI60/XI13/MM2_g N_VSS_XI60/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI13/MM3 N_XI60/XI13/NET33_XI60/XI13/MM3_d N_WL<116>_XI60/XI13/MM3_g
+ N_BLN<2>_XI60/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI13/MM0 N_XI60/XI13/NET34_XI60/XI13/MM0_d N_WL<116>_XI60/XI13/MM0_g
+ N_BL<2>_XI60/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI13/MM1 N_XI60/XI13/NET33_XI60/XI13/MM1_d
+ N_XI60/XI13/NET34_XI60/XI13/MM1_g N_VSS_XI60/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI13/MM9 N_XI60/XI13/NET36_XI60/XI13/MM9_d N_WL<117>_XI60/XI13/MM9_g
+ N_BL<2>_XI60/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI13/MM6 N_XI60/XI13/NET35_XI60/XI13/MM6_d
+ N_XI60/XI13/NET36_XI60/XI13/MM6_g N_VSS_XI60/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI13/MM7 N_XI60/XI13/NET36_XI60/XI13/MM7_d
+ N_XI60/XI13/NET35_XI60/XI13/MM7_g N_VSS_XI60/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI13/MM8 N_XI60/XI13/NET35_XI60/XI13/MM8_d N_WL<117>_XI60/XI13/MM8_g
+ N_BLN<2>_XI60/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI13/MM5 N_XI60/XI13/NET34_XI60/XI13/MM5_d
+ N_XI60/XI13/NET33_XI60/XI13/MM5_g N_VDD_XI60/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI13/MM4 N_XI60/XI13/NET33_XI60/XI13/MM4_d
+ N_XI60/XI13/NET34_XI60/XI13/MM4_g N_VDD_XI60/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI13/MM10 N_XI60/XI13/NET35_XI60/XI13/MM10_d
+ N_XI60/XI13/NET36_XI60/XI13/MM10_g N_VDD_XI60/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI13/MM11 N_XI60/XI13/NET36_XI60/XI13/MM11_d
+ N_XI60/XI13/NET35_XI60/XI13/MM11_g N_VDD_XI60/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI14/MM2 N_XI60/XI14/NET34_XI60/XI14/MM2_d
+ N_XI60/XI14/NET33_XI60/XI14/MM2_g N_VSS_XI60/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI14/MM3 N_XI60/XI14/NET33_XI60/XI14/MM3_d N_WL<116>_XI60/XI14/MM3_g
+ N_BLN<1>_XI60/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI14/MM0 N_XI60/XI14/NET34_XI60/XI14/MM0_d N_WL<116>_XI60/XI14/MM0_g
+ N_BL<1>_XI60/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI14/MM1 N_XI60/XI14/NET33_XI60/XI14/MM1_d
+ N_XI60/XI14/NET34_XI60/XI14/MM1_g N_VSS_XI60/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI14/MM9 N_XI60/XI14/NET36_XI60/XI14/MM9_d N_WL<117>_XI60/XI14/MM9_g
+ N_BL<1>_XI60/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI14/MM6 N_XI60/XI14/NET35_XI60/XI14/MM6_d
+ N_XI60/XI14/NET36_XI60/XI14/MM6_g N_VSS_XI60/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI14/MM7 N_XI60/XI14/NET36_XI60/XI14/MM7_d
+ N_XI60/XI14/NET35_XI60/XI14/MM7_g N_VSS_XI60/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI14/MM8 N_XI60/XI14/NET35_XI60/XI14/MM8_d N_WL<117>_XI60/XI14/MM8_g
+ N_BLN<1>_XI60/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI14/MM5 N_XI60/XI14/NET34_XI60/XI14/MM5_d
+ N_XI60/XI14/NET33_XI60/XI14/MM5_g N_VDD_XI60/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI14/MM4 N_XI60/XI14/NET33_XI60/XI14/MM4_d
+ N_XI60/XI14/NET34_XI60/XI14/MM4_g N_VDD_XI60/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI14/MM10 N_XI60/XI14/NET35_XI60/XI14/MM10_d
+ N_XI60/XI14/NET36_XI60/XI14/MM10_g N_VDD_XI60/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI14/MM11 N_XI60/XI14/NET36_XI60/XI14/MM11_d
+ N_XI60/XI14/NET35_XI60/XI14/MM11_g N_VDD_XI60/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI15/MM2 N_XI60/XI15/NET34_XI60/XI15/MM2_d
+ N_XI60/XI15/NET33_XI60/XI15/MM2_g N_VSS_XI60/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI15/MM3 N_XI60/XI15/NET33_XI60/XI15/MM3_d N_WL<116>_XI60/XI15/MM3_g
+ N_BLN<0>_XI60/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI15/MM0 N_XI60/XI15/NET34_XI60/XI15/MM0_d N_WL<116>_XI60/XI15/MM0_g
+ N_BL<0>_XI60/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI15/MM1 N_XI60/XI15/NET33_XI60/XI15/MM1_d
+ N_XI60/XI15/NET34_XI60/XI15/MM1_g N_VSS_XI60/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI15/MM9 N_XI60/XI15/NET36_XI60/XI15/MM9_d N_WL<117>_XI60/XI15/MM9_g
+ N_BL<0>_XI60/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI15/MM6 N_XI60/XI15/NET35_XI60/XI15/MM6_d
+ N_XI60/XI15/NET36_XI60/XI15/MM6_g N_VSS_XI60/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI15/MM7 N_XI60/XI15/NET36_XI60/XI15/MM7_d
+ N_XI60/XI15/NET35_XI60/XI15/MM7_g N_VSS_XI60/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI60/XI15/MM8 N_XI60/XI15/NET35_XI60/XI15/MM8_d N_WL<117>_XI60/XI15/MM8_g
+ N_BLN<0>_XI60/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI60/XI15/MM5 N_XI60/XI15/NET34_XI60/XI15/MM5_d
+ N_XI60/XI15/NET33_XI60/XI15/MM5_g N_VDD_XI60/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI15/MM4 N_XI60/XI15/NET33_XI60/XI15/MM4_d
+ N_XI60/XI15/NET34_XI60/XI15/MM4_g N_VDD_XI60/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI15/MM10 N_XI60/XI15/NET35_XI60/XI15/MM10_d
+ N_XI60/XI15/NET36_XI60/XI15/MM10_g N_VDD_XI60/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI60/XI15/MM11 N_XI60/XI15/NET36_XI60/XI15/MM11_d
+ N_XI60/XI15/NET35_XI60/XI15/MM11_g N_VDD_XI60/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI0/MM2 N_XI61/XI0/NET34_XI61/XI0/MM2_d N_XI61/XI0/NET33_XI61/XI0/MM2_g
+ N_VSS_XI61/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI0/MM3 N_XI61/XI0/NET33_XI61/XI0/MM3_d N_WL<118>_XI61/XI0/MM3_g
+ N_BLN<15>_XI61/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI0/MM0 N_XI61/XI0/NET34_XI61/XI0/MM0_d N_WL<118>_XI61/XI0/MM0_g
+ N_BL<15>_XI61/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI0/MM1 N_XI61/XI0/NET33_XI61/XI0/MM1_d N_XI61/XI0/NET34_XI61/XI0/MM1_g
+ N_VSS_XI61/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI0/MM9 N_XI61/XI0/NET36_XI61/XI0/MM9_d N_WL<119>_XI61/XI0/MM9_g
+ N_BL<15>_XI61/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI0/MM6 N_XI61/XI0/NET35_XI61/XI0/MM6_d N_XI61/XI0/NET36_XI61/XI0/MM6_g
+ N_VSS_XI61/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI0/MM7 N_XI61/XI0/NET36_XI61/XI0/MM7_d N_XI61/XI0/NET35_XI61/XI0/MM7_g
+ N_VSS_XI61/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI0/MM8 N_XI61/XI0/NET35_XI61/XI0/MM8_d N_WL<119>_XI61/XI0/MM8_g
+ N_BLN<15>_XI61/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI0/MM5 N_XI61/XI0/NET34_XI61/XI0/MM5_d N_XI61/XI0/NET33_XI61/XI0/MM5_g
+ N_VDD_XI61/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI0/MM4 N_XI61/XI0/NET33_XI61/XI0/MM4_d N_XI61/XI0/NET34_XI61/XI0/MM4_g
+ N_VDD_XI61/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI0/MM10 N_XI61/XI0/NET35_XI61/XI0/MM10_d N_XI61/XI0/NET36_XI61/XI0/MM10_g
+ N_VDD_XI61/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI0/MM11 N_XI61/XI0/NET36_XI61/XI0/MM11_d N_XI61/XI0/NET35_XI61/XI0/MM11_g
+ N_VDD_XI61/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI1/MM2 N_XI61/XI1/NET34_XI61/XI1/MM2_d N_XI61/XI1/NET33_XI61/XI1/MM2_g
+ N_VSS_XI61/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI1/MM3 N_XI61/XI1/NET33_XI61/XI1/MM3_d N_WL<118>_XI61/XI1/MM3_g
+ N_BLN<14>_XI61/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI1/MM0 N_XI61/XI1/NET34_XI61/XI1/MM0_d N_WL<118>_XI61/XI1/MM0_g
+ N_BL<14>_XI61/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI1/MM1 N_XI61/XI1/NET33_XI61/XI1/MM1_d N_XI61/XI1/NET34_XI61/XI1/MM1_g
+ N_VSS_XI61/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI1/MM9 N_XI61/XI1/NET36_XI61/XI1/MM9_d N_WL<119>_XI61/XI1/MM9_g
+ N_BL<14>_XI61/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI1/MM6 N_XI61/XI1/NET35_XI61/XI1/MM6_d N_XI61/XI1/NET36_XI61/XI1/MM6_g
+ N_VSS_XI61/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI1/MM7 N_XI61/XI1/NET36_XI61/XI1/MM7_d N_XI61/XI1/NET35_XI61/XI1/MM7_g
+ N_VSS_XI61/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI1/MM8 N_XI61/XI1/NET35_XI61/XI1/MM8_d N_WL<119>_XI61/XI1/MM8_g
+ N_BLN<14>_XI61/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI1/MM5 N_XI61/XI1/NET34_XI61/XI1/MM5_d N_XI61/XI1/NET33_XI61/XI1/MM5_g
+ N_VDD_XI61/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI1/MM4 N_XI61/XI1/NET33_XI61/XI1/MM4_d N_XI61/XI1/NET34_XI61/XI1/MM4_g
+ N_VDD_XI61/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI1/MM10 N_XI61/XI1/NET35_XI61/XI1/MM10_d N_XI61/XI1/NET36_XI61/XI1/MM10_g
+ N_VDD_XI61/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI1/MM11 N_XI61/XI1/NET36_XI61/XI1/MM11_d N_XI61/XI1/NET35_XI61/XI1/MM11_g
+ N_VDD_XI61/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI2/MM2 N_XI61/XI2/NET34_XI61/XI2/MM2_d N_XI61/XI2/NET33_XI61/XI2/MM2_g
+ N_VSS_XI61/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI2/MM3 N_XI61/XI2/NET33_XI61/XI2/MM3_d N_WL<118>_XI61/XI2/MM3_g
+ N_BLN<13>_XI61/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI2/MM0 N_XI61/XI2/NET34_XI61/XI2/MM0_d N_WL<118>_XI61/XI2/MM0_g
+ N_BL<13>_XI61/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI2/MM1 N_XI61/XI2/NET33_XI61/XI2/MM1_d N_XI61/XI2/NET34_XI61/XI2/MM1_g
+ N_VSS_XI61/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI2/MM9 N_XI61/XI2/NET36_XI61/XI2/MM9_d N_WL<119>_XI61/XI2/MM9_g
+ N_BL<13>_XI61/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI2/MM6 N_XI61/XI2/NET35_XI61/XI2/MM6_d N_XI61/XI2/NET36_XI61/XI2/MM6_g
+ N_VSS_XI61/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI2/MM7 N_XI61/XI2/NET36_XI61/XI2/MM7_d N_XI61/XI2/NET35_XI61/XI2/MM7_g
+ N_VSS_XI61/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI2/MM8 N_XI61/XI2/NET35_XI61/XI2/MM8_d N_WL<119>_XI61/XI2/MM8_g
+ N_BLN<13>_XI61/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI2/MM5 N_XI61/XI2/NET34_XI61/XI2/MM5_d N_XI61/XI2/NET33_XI61/XI2/MM5_g
+ N_VDD_XI61/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI2/MM4 N_XI61/XI2/NET33_XI61/XI2/MM4_d N_XI61/XI2/NET34_XI61/XI2/MM4_g
+ N_VDD_XI61/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI2/MM10 N_XI61/XI2/NET35_XI61/XI2/MM10_d N_XI61/XI2/NET36_XI61/XI2/MM10_g
+ N_VDD_XI61/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI2/MM11 N_XI61/XI2/NET36_XI61/XI2/MM11_d N_XI61/XI2/NET35_XI61/XI2/MM11_g
+ N_VDD_XI61/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI3/MM2 N_XI61/XI3/NET34_XI61/XI3/MM2_d N_XI61/XI3/NET33_XI61/XI3/MM2_g
+ N_VSS_XI61/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI3/MM3 N_XI61/XI3/NET33_XI61/XI3/MM3_d N_WL<118>_XI61/XI3/MM3_g
+ N_BLN<12>_XI61/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI3/MM0 N_XI61/XI3/NET34_XI61/XI3/MM0_d N_WL<118>_XI61/XI3/MM0_g
+ N_BL<12>_XI61/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI3/MM1 N_XI61/XI3/NET33_XI61/XI3/MM1_d N_XI61/XI3/NET34_XI61/XI3/MM1_g
+ N_VSS_XI61/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI3/MM9 N_XI61/XI3/NET36_XI61/XI3/MM9_d N_WL<119>_XI61/XI3/MM9_g
+ N_BL<12>_XI61/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI3/MM6 N_XI61/XI3/NET35_XI61/XI3/MM6_d N_XI61/XI3/NET36_XI61/XI3/MM6_g
+ N_VSS_XI61/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI3/MM7 N_XI61/XI3/NET36_XI61/XI3/MM7_d N_XI61/XI3/NET35_XI61/XI3/MM7_g
+ N_VSS_XI61/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI3/MM8 N_XI61/XI3/NET35_XI61/XI3/MM8_d N_WL<119>_XI61/XI3/MM8_g
+ N_BLN<12>_XI61/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI3/MM5 N_XI61/XI3/NET34_XI61/XI3/MM5_d N_XI61/XI3/NET33_XI61/XI3/MM5_g
+ N_VDD_XI61/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI3/MM4 N_XI61/XI3/NET33_XI61/XI3/MM4_d N_XI61/XI3/NET34_XI61/XI3/MM4_g
+ N_VDD_XI61/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI3/MM10 N_XI61/XI3/NET35_XI61/XI3/MM10_d N_XI61/XI3/NET36_XI61/XI3/MM10_g
+ N_VDD_XI61/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI3/MM11 N_XI61/XI3/NET36_XI61/XI3/MM11_d N_XI61/XI3/NET35_XI61/XI3/MM11_g
+ N_VDD_XI61/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI4/MM2 N_XI61/XI4/NET34_XI61/XI4/MM2_d N_XI61/XI4/NET33_XI61/XI4/MM2_g
+ N_VSS_XI61/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI4/MM3 N_XI61/XI4/NET33_XI61/XI4/MM3_d N_WL<118>_XI61/XI4/MM3_g
+ N_BLN<11>_XI61/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI4/MM0 N_XI61/XI4/NET34_XI61/XI4/MM0_d N_WL<118>_XI61/XI4/MM0_g
+ N_BL<11>_XI61/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI4/MM1 N_XI61/XI4/NET33_XI61/XI4/MM1_d N_XI61/XI4/NET34_XI61/XI4/MM1_g
+ N_VSS_XI61/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI4/MM9 N_XI61/XI4/NET36_XI61/XI4/MM9_d N_WL<119>_XI61/XI4/MM9_g
+ N_BL<11>_XI61/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI4/MM6 N_XI61/XI4/NET35_XI61/XI4/MM6_d N_XI61/XI4/NET36_XI61/XI4/MM6_g
+ N_VSS_XI61/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI4/MM7 N_XI61/XI4/NET36_XI61/XI4/MM7_d N_XI61/XI4/NET35_XI61/XI4/MM7_g
+ N_VSS_XI61/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI4/MM8 N_XI61/XI4/NET35_XI61/XI4/MM8_d N_WL<119>_XI61/XI4/MM8_g
+ N_BLN<11>_XI61/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI4/MM5 N_XI61/XI4/NET34_XI61/XI4/MM5_d N_XI61/XI4/NET33_XI61/XI4/MM5_g
+ N_VDD_XI61/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI4/MM4 N_XI61/XI4/NET33_XI61/XI4/MM4_d N_XI61/XI4/NET34_XI61/XI4/MM4_g
+ N_VDD_XI61/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI4/MM10 N_XI61/XI4/NET35_XI61/XI4/MM10_d N_XI61/XI4/NET36_XI61/XI4/MM10_g
+ N_VDD_XI61/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI4/MM11 N_XI61/XI4/NET36_XI61/XI4/MM11_d N_XI61/XI4/NET35_XI61/XI4/MM11_g
+ N_VDD_XI61/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI5/MM2 N_XI61/XI5/NET34_XI61/XI5/MM2_d N_XI61/XI5/NET33_XI61/XI5/MM2_g
+ N_VSS_XI61/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI5/MM3 N_XI61/XI5/NET33_XI61/XI5/MM3_d N_WL<118>_XI61/XI5/MM3_g
+ N_BLN<10>_XI61/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI5/MM0 N_XI61/XI5/NET34_XI61/XI5/MM0_d N_WL<118>_XI61/XI5/MM0_g
+ N_BL<10>_XI61/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI5/MM1 N_XI61/XI5/NET33_XI61/XI5/MM1_d N_XI61/XI5/NET34_XI61/XI5/MM1_g
+ N_VSS_XI61/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI5/MM9 N_XI61/XI5/NET36_XI61/XI5/MM9_d N_WL<119>_XI61/XI5/MM9_g
+ N_BL<10>_XI61/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI5/MM6 N_XI61/XI5/NET35_XI61/XI5/MM6_d N_XI61/XI5/NET36_XI61/XI5/MM6_g
+ N_VSS_XI61/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI5/MM7 N_XI61/XI5/NET36_XI61/XI5/MM7_d N_XI61/XI5/NET35_XI61/XI5/MM7_g
+ N_VSS_XI61/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI5/MM8 N_XI61/XI5/NET35_XI61/XI5/MM8_d N_WL<119>_XI61/XI5/MM8_g
+ N_BLN<10>_XI61/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI5/MM5 N_XI61/XI5/NET34_XI61/XI5/MM5_d N_XI61/XI5/NET33_XI61/XI5/MM5_g
+ N_VDD_XI61/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI5/MM4 N_XI61/XI5/NET33_XI61/XI5/MM4_d N_XI61/XI5/NET34_XI61/XI5/MM4_g
+ N_VDD_XI61/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI5/MM10 N_XI61/XI5/NET35_XI61/XI5/MM10_d N_XI61/XI5/NET36_XI61/XI5/MM10_g
+ N_VDD_XI61/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI5/MM11 N_XI61/XI5/NET36_XI61/XI5/MM11_d N_XI61/XI5/NET35_XI61/XI5/MM11_g
+ N_VDD_XI61/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI6/MM2 N_XI61/XI6/NET34_XI61/XI6/MM2_d N_XI61/XI6/NET33_XI61/XI6/MM2_g
+ N_VSS_XI61/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM3 N_XI61/XI6/NET33_XI61/XI6/MM3_d N_WL<118>_XI61/XI6/MM3_g
+ N_BLN<9>_XI61/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM0 N_XI61/XI6/NET34_XI61/XI6/MM0_d N_WL<118>_XI61/XI6/MM0_g
+ N_BL<9>_XI61/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM1 N_XI61/XI6/NET33_XI61/XI6/MM1_d N_XI61/XI6/NET34_XI61/XI6/MM1_g
+ N_VSS_XI61/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM9 N_XI61/XI6/NET36_XI61/XI6/MM9_d N_WL<119>_XI61/XI6/MM9_g
+ N_BL<9>_XI61/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM6 N_XI61/XI6/NET35_XI61/XI6/MM6_d N_XI61/XI6/NET36_XI61/XI6/MM6_g
+ N_VSS_XI61/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM7 N_XI61/XI6/NET36_XI61/XI6/MM7_d N_XI61/XI6/NET35_XI61/XI6/MM7_g
+ N_VSS_XI61/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM8 N_XI61/XI6/NET35_XI61/XI6/MM8_d N_WL<119>_XI61/XI6/MM8_g
+ N_BLN<9>_XI61/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI6/MM5 N_XI61/XI6/NET34_XI61/XI6/MM5_d N_XI61/XI6/NET33_XI61/XI6/MM5_g
+ N_VDD_XI61/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI6/MM4 N_XI61/XI6/NET33_XI61/XI6/MM4_d N_XI61/XI6/NET34_XI61/XI6/MM4_g
+ N_VDD_XI61/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI6/MM10 N_XI61/XI6/NET35_XI61/XI6/MM10_d N_XI61/XI6/NET36_XI61/XI6/MM10_g
+ N_VDD_XI61/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI6/MM11 N_XI61/XI6/NET36_XI61/XI6/MM11_d N_XI61/XI6/NET35_XI61/XI6/MM11_g
+ N_VDD_XI61/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI7/MM2 N_XI61/XI7/NET34_XI61/XI7/MM2_d N_XI61/XI7/NET33_XI61/XI7/MM2_g
+ N_VSS_XI61/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM3 N_XI61/XI7/NET33_XI61/XI7/MM3_d N_WL<118>_XI61/XI7/MM3_g
+ N_BLN<8>_XI61/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM0 N_XI61/XI7/NET34_XI61/XI7/MM0_d N_WL<118>_XI61/XI7/MM0_g
+ N_BL<8>_XI61/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM1 N_XI61/XI7/NET33_XI61/XI7/MM1_d N_XI61/XI7/NET34_XI61/XI7/MM1_g
+ N_VSS_XI61/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM9 N_XI61/XI7/NET36_XI61/XI7/MM9_d N_WL<119>_XI61/XI7/MM9_g
+ N_BL<8>_XI61/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM6 N_XI61/XI7/NET35_XI61/XI7/MM6_d N_XI61/XI7/NET36_XI61/XI7/MM6_g
+ N_VSS_XI61/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM7 N_XI61/XI7/NET36_XI61/XI7/MM7_d N_XI61/XI7/NET35_XI61/XI7/MM7_g
+ N_VSS_XI61/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM8 N_XI61/XI7/NET35_XI61/XI7/MM8_d N_WL<119>_XI61/XI7/MM8_g
+ N_BLN<8>_XI61/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI7/MM5 N_XI61/XI7/NET34_XI61/XI7/MM5_d N_XI61/XI7/NET33_XI61/XI7/MM5_g
+ N_VDD_XI61/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI7/MM4 N_XI61/XI7/NET33_XI61/XI7/MM4_d N_XI61/XI7/NET34_XI61/XI7/MM4_g
+ N_VDD_XI61/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI7/MM10 N_XI61/XI7/NET35_XI61/XI7/MM10_d N_XI61/XI7/NET36_XI61/XI7/MM10_g
+ N_VDD_XI61/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI7/MM11 N_XI61/XI7/NET36_XI61/XI7/MM11_d N_XI61/XI7/NET35_XI61/XI7/MM11_g
+ N_VDD_XI61/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI8/MM2 N_XI61/XI8/NET34_XI61/XI8/MM2_d N_XI61/XI8/NET33_XI61/XI8/MM2_g
+ N_VSS_XI61/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM3 N_XI61/XI8/NET33_XI61/XI8/MM3_d N_WL<118>_XI61/XI8/MM3_g
+ N_BLN<7>_XI61/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM0 N_XI61/XI8/NET34_XI61/XI8/MM0_d N_WL<118>_XI61/XI8/MM0_g
+ N_BL<7>_XI61/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM1 N_XI61/XI8/NET33_XI61/XI8/MM1_d N_XI61/XI8/NET34_XI61/XI8/MM1_g
+ N_VSS_XI61/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM9 N_XI61/XI8/NET36_XI61/XI8/MM9_d N_WL<119>_XI61/XI8/MM9_g
+ N_BL<7>_XI61/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM6 N_XI61/XI8/NET35_XI61/XI8/MM6_d N_XI61/XI8/NET36_XI61/XI8/MM6_g
+ N_VSS_XI61/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM7 N_XI61/XI8/NET36_XI61/XI8/MM7_d N_XI61/XI8/NET35_XI61/XI8/MM7_g
+ N_VSS_XI61/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM8 N_XI61/XI8/NET35_XI61/XI8/MM8_d N_WL<119>_XI61/XI8/MM8_g
+ N_BLN<7>_XI61/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI8/MM5 N_XI61/XI8/NET34_XI61/XI8/MM5_d N_XI61/XI8/NET33_XI61/XI8/MM5_g
+ N_VDD_XI61/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI8/MM4 N_XI61/XI8/NET33_XI61/XI8/MM4_d N_XI61/XI8/NET34_XI61/XI8/MM4_g
+ N_VDD_XI61/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI8/MM10 N_XI61/XI8/NET35_XI61/XI8/MM10_d N_XI61/XI8/NET36_XI61/XI8/MM10_g
+ N_VDD_XI61/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI8/MM11 N_XI61/XI8/NET36_XI61/XI8/MM11_d N_XI61/XI8/NET35_XI61/XI8/MM11_g
+ N_VDD_XI61/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI9/MM2 N_XI61/XI9/NET34_XI61/XI9/MM2_d N_XI61/XI9/NET33_XI61/XI9/MM2_g
+ N_VSS_XI61/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM3 N_XI61/XI9/NET33_XI61/XI9/MM3_d N_WL<118>_XI61/XI9/MM3_g
+ N_BLN<6>_XI61/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM0 N_XI61/XI9/NET34_XI61/XI9/MM0_d N_WL<118>_XI61/XI9/MM0_g
+ N_BL<6>_XI61/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM1 N_XI61/XI9/NET33_XI61/XI9/MM1_d N_XI61/XI9/NET34_XI61/XI9/MM1_g
+ N_VSS_XI61/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM9 N_XI61/XI9/NET36_XI61/XI9/MM9_d N_WL<119>_XI61/XI9/MM9_g
+ N_BL<6>_XI61/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM6 N_XI61/XI9/NET35_XI61/XI9/MM6_d N_XI61/XI9/NET36_XI61/XI9/MM6_g
+ N_VSS_XI61/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM7 N_XI61/XI9/NET36_XI61/XI9/MM7_d N_XI61/XI9/NET35_XI61/XI9/MM7_g
+ N_VSS_XI61/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM8 N_XI61/XI9/NET35_XI61/XI9/MM8_d N_WL<119>_XI61/XI9/MM8_g
+ N_BLN<6>_XI61/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI9/MM5 N_XI61/XI9/NET34_XI61/XI9/MM5_d N_XI61/XI9/NET33_XI61/XI9/MM5_g
+ N_VDD_XI61/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI9/MM4 N_XI61/XI9/NET33_XI61/XI9/MM4_d N_XI61/XI9/NET34_XI61/XI9/MM4_g
+ N_VDD_XI61/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI9/MM10 N_XI61/XI9/NET35_XI61/XI9/MM10_d N_XI61/XI9/NET36_XI61/XI9/MM10_g
+ N_VDD_XI61/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI9/MM11 N_XI61/XI9/NET36_XI61/XI9/MM11_d N_XI61/XI9/NET35_XI61/XI9/MM11_g
+ N_VDD_XI61/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI10/MM2 N_XI61/XI10/NET34_XI61/XI10/MM2_d
+ N_XI61/XI10/NET33_XI61/XI10/MM2_g N_VSS_XI61/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI10/MM3 N_XI61/XI10/NET33_XI61/XI10/MM3_d N_WL<118>_XI61/XI10/MM3_g
+ N_BLN<5>_XI61/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI10/MM0 N_XI61/XI10/NET34_XI61/XI10/MM0_d N_WL<118>_XI61/XI10/MM0_g
+ N_BL<5>_XI61/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI10/MM1 N_XI61/XI10/NET33_XI61/XI10/MM1_d
+ N_XI61/XI10/NET34_XI61/XI10/MM1_g N_VSS_XI61/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI10/MM9 N_XI61/XI10/NET36_XI61/XI10/MM9_d N_WL<119>_XI61/XI10/MM9_g
+ N_BL<5>_XI61/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI10/MM6 N_XI61/XI10/NET35_XI61/XI10/MM6_d
+ N_XI61/XI10/NET36_XI61/XI10/MM6_g N_VSS_XI61/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI10/MM7 N_XI61/XI10/NET36_XI61/XI10/MM7_d
+ N_XI61/XI10/NET35_XI61/XI10/MM7_g N_VSS_XI61/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI10/MM8 N_XI61/XI10/NET35_XI61/XI10/MM8_d N_WL<119>_XI61/XI10/MM8_g
+ N_BLN<5>_XI61/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI10/MM5 N_XI61/XI10/NET34_XI61/XI10/MM5_d
+ N_XI61/XI10/NET33_XI61/XI10/MM5_g N_VDD_XI61/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI10/MM4 N_XI61/XI10/NET33_XI61/XI10/MM4_d
+ N_XI61/XI10/NET34_XI61/XI10/MM4_g N_VDD_XI61/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI10/MM10 N_XI61/XI10/NET35_XI61/XI10/MM10_d
+ N_XI61/XI10/NET36_XI61/XI10/MM10_g N_VDD_XI61/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI10/MM11 N_XI61/XI10/NET36_XI61/XI10/MM11_d
+ N_XI61/XI10/NET35_XI61/XI10/MM11_g N_VDD_XI61/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI11/MM2 N_XI61/XI11/NET34_XI61/XI11/MM2_d
+ N_XI61/XI11/NET33_XI61/XI11/MM2_g N_VSS_XI61/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI11/MM3 N_XI61/XI11/NET33_XI61/XI11/MM3_d N_WL<118>_XI61/XI11/MM3_g
+ N_BLN<4>_XI61/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI11/MM0 N_XI61/XI11/NET34_XI61/XI11/MM0_d N_WL<118>_XI61/XI11/MM0_g
+ N_BL<4>_XI61/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI11/MM1 N_XI61/XI11/NET33_XI61/XI11/MM1_d
+ N_XI61/XI11/NET34_XI61/XI11/MM1_g N_VSS_XI61/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI11/MM9 N_XI61/XI11/NET36_XI61/XI11/MM9_d N_WL<119>_XI61/XI11/MM9_g
+ N_BL<4>_XI61/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI11/MM6 N_XI61/XI11/NET35_XI61/XI11/MM6_d
+ N_XI61/XI11/NET36_XI61/XI11/MM6_g N_VSS_XI61/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI11/MM7 N_XI61/XI11/NET36_XI61/XI11/MM7_d
+ N_XI61/XI11/NET35_XI61/XI11/MM7_g N_VSS_XI61/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI11/MM8 N_XI61/XI11/NET35_XI61/XI11/MM8_d N_WL<119>_XI61/XI11/MM8_g
+ N_BLN<4>_XI61/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI11/MM5 N_XI61/XI11/NET34_XI61/XI11/MM5_d
+ N_XI61/XI11/NET33_XI61/XI11/MM5_g N_VDD_XI61/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI11/MM4 N_XI61/XI11/NET33_XI61/XI11/MM4_d
+ N_XI61/XI11/NET34_XI61/XI11/MM4_g N_VDD_XI61/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI11/MM10 N_XI61/XI11/NET35_XI61/XI11/MM10_d
+ N_XI61/XI11/NET36_XI61/XI11/MM10_g N_VDD_XI61/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI11/MM11 N_XI61/XI11/NET36_XI61/XI11/MM11_d
+ N_XI61/XI11/NET35_XI61/XI11/MM11_g N_VDD_XI61/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI12/MM2 N_XI61/XI12/NET34_XI61/XI12/MM2_d
+ N_XI61/XI12/NET33_XI61/XI12/MM2_g N_VSS_XI61/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI12/MM3 N_XI61/XI12/NET33_XI61/XI12/MM3_d N_WL<118>_XI61/XI12/MM3_g
+ N_BLN<3>_XI61/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI12/MM0 N_XI61/XI12/NET34_XI61/XI12/MM0_d N_WL<118>_XI61/XI12/MM0_g
+ N_BL<3>_XI61/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI12/MM1 N_XI61/XI12/NET33_XI61/XI12/MM1_d
+ N_XI61/XI12/NET34_XI61/XI12/MM1_g N_VSS_XI61/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI12/MM9 N_XI61/XI12/NET36_XI61/XI12/MM9_d N_WL<119>_XI61/XI12/MM9_g
+ N_BL<3>_XI61/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI12/MM6 N_XI61/XI12/NET35_XI61/XI12/MM6_d
+ N_XI61/XI12/NET36_XI61/XI12/MM6_g N_VSS_XI61/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI12/MM7 N_XI61/XI12/NET36_XI61/XI12/MM7_d
+ N_XI61/XI12/NET35_XI61/XI12/MM7_g N_VSS_XI61/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI12/MM8 N_XI61/XI12/NET35_XI61/XI12/MM8_d N_WL<119>_XI61/XI12/MM8_g
+ N_BLN<3>_XI61/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI12/MM5 N_XI61/XI12/NET34_XI61/XI12/MM5_d
+ N_XI61/XI12/NET33_XI61/XI12/MM5_g N_VDD_XI61/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI12/MM4 N_XI61/XI12/NET33_XI61/XI12/MM4_d
+ N_XI61/XI12/NET34_XI61/XI12/MM4_g N_VDD_XI61/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI12/MM10 N_XI61/XI12/NET35_XI61/XI12/MM10_d
+ N_XI61/XI12/NET36_XI61/XI12/MM10_g N_VDD_XI61/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI12/MM11 N_XI61/XI12/NET36_XI61/XI12/MM11_d
+ N_XI61/XI12/NET35_XI61/XI12/MM11_g N_VDD_XI61/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI13/MM2 N_XI61/XI13/NET34_XI61/XI13/MM2_d
+ N_XI61/XI13/NET33_XI61/XI13/MM2_g N_VSS_XI61/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI13/MM3 N_XI61/XI13/NET33_XI61/XI13/MM3_d N_WL<118>_XI61/XI13/MM3_g
+ N_BLN<2>_XI61/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI13/MM0 N_XI61/XI13/NET34_XI61/XI13/MM0_d N_WL<118>_XI61/XI13/MM0_g
+ N_BL<2>_XI61/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI13/MM1 N_XI61/XI13/NET33_XI61/XI13/MM1_d
+ N_XI61/XI13/NET34_XI61/XI13/MM1_g N_VSS_XI61/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI13/MM9 N_XI61/XI13/NET36_XI61/XI13/MM9_d N_WL<119>_XI61/XI13/MM9_g
+ N_BL<2>_XI61/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI13/MM6 N_XI61/XI13/NET35_XI61/XI13/MM6_d
+ N_XI61/XI13/NET36_XI61/XI13/MM6_g N_VSS_XI61/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI13/MM7 N_XI61/XI13/NET36_XI61/XI13/MM7_d
+ N_XI61/XI13/NET35_XI61/XI13/MM7_g N_VSS_XI61/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI13/MM8 N_XI61/XI13/NET35_XI61/XI13/MM8_d N_WL<119>_XI61/XI13/MM8_g
+ N_BLN<2>_XI61/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI13/MM5 N_XI61/XI13/NET34_XI61/XI13/MM5_d
+ N_XI61/XI13/NET33_XI61/XI13/MM5_g N_VDD_XI61/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI13/MM4 N_XI61/XI13/NET33_XI61/XI13/MM4_d
+ N_XI61/XI13/NET34_XI61/XI13/MM4_g N_VDD_XI61/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI13/MM10 N_XI61/XI13/NET35_XI61/XI13/MM10_d
+ N_XI61/XI13/NET36_XI61/XI13/MM10_g N_VDD_XI61/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI13/MM11 N_XI61/XI13/NET36_XI61/XI13/MM11_d
+ N_XI61/XI13/NET35_XI61/XI13/MM11_g N_VDD_XI61/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI14/MM2 N_XI61/XI14/NET34_XI61/XI14/MM2_d
+ N_XI61/XI14/NET33_XI61/XI14/MM2_g N_VSS_XI61/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI14/MM3 N_XI61/XI14/NET33_XI61/XI14/MM3_d N_WL<118>_XI61/XI14/MM3_g
+ N_BLN<1>_XI61/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI14/MM0 N_XI61/XI14/NET34_XI61/XI14/MM0_d N_WL<118>_XI61/XI14/MM0_g
+ N_BL<1>_XI61/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI14/MM1 N_XI61/XI14/NET33_XI61/XI14/MM1_d
+ N_XI61/XI14/NET34_XI61/XI14/MM1_g N_VSS_XI61/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI14/MM9 N_XI61/XI14/NET36_XI61/XI14/MM9_d N_WL<119>_XI61/XI14/MM9_g
+ N_BL<1>_XI61/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI14/MM6 N_XI61/XI14/NET35_XI61/XI14/MM6_d
+ N_XI61/XI14/NET36_XI61/XI14/MM6_g N_VSS_XI61/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI14/MM7 N_XI61/XI14/NET36_XI61/XI14/MM7_d
+ N_XI61/XI14/NET35_XI61/XI14/MM7_g N_VSS_XI61/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI14/MM8 N_XI61/XI14/NET35_XI61/XI14/MM8_d N_WL<119>_XI61/XI14/MM8_g
+ N_BLN<1>_XI61/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI14/MM5 N_XI61/XI14/NET34_XI61/XI14/MM5_d
+ N_XI61/XI14/NET33_XI61/XI14/MM5_g N_VDD_XI61/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI14/MM4 N_XI61/XI14/NET33_XI61/XI14/MM4_d
+ N_XI61/XI14/NET34_XI61/XI14/MM4_g N_VDD_XI61/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI14/MM10 N_XI61/XI14/NET35_XI61/XI14/MM10_d
+ N_XI61/XI14/NET36_XI61/XI14/MM10_g N_VDD_XI61/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI14/MM11 N_XI61/XI14/NET36_XI61/XI14/MM11_d
+ N_XI61/XI14/NET35_XI61/XI14/MM11_g N_VDD_XI61/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI15/MM2 N_XI61/XI15/NET34_XI61/XI15/MM2_d
+ N_XI61/XI15/NET33_XI61/XI15/MM2_g N_VSS_XI61/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI15/MM3 N_XI61/XI15/NET33_XI61/XI15/MM3_d N_WL<118>_XI61/XI15/MM3_g
+ N_BLN<0>_XI61/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI15/MM0 N_XI61/XI15/NET34_XI61/XI15/MM0_d N_WL<118>_XI61/XI15/MM0_g
+ N_BL<0>_XI61/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI15/MM1 N_XI61/XI15/NET33_XI61/XI15/MM1_d
+ N_XI61/XI15/NET34_XI61/XI15/MM1_g N_VSS_XI61/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI15/MM9 N_XI61/XI15/NET36_XI61/XI15/MM9_d N_WL<119>_XI61/XI15/MM9_g
+ N_BL<0>_XI61/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI15/MM6 N_XI61/XI15/NET35_XI61/XI15/MM6_d
+ N_XI61/XI15/NET36_XI61/XI15/MM6_g N_VSS_XI61/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI15/MM7 N_XI61/XI15/NET36_XI61/XI15/MM7_d
+ N_XI61/XI15/NET35_XI61/XI15/MM7_g N_VSS_XI61/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI61/XI15/MM8 N_XI61/XI15/NET35_XI61/XI15/MM8_d N_WL<119>_XI61/XI15/MM8_g
+ N_BLN<0>_XI61/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI61/XI15/MM5 N_XI61/XI15/NET34_XI61/XI15/MM5_d
+ N_XI61/XI15/NET33_XI61/XI15/MM5_g N_VDD_XI61/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI15/MM4 N_XI61/XI15/NET33_XI61/XI15/MM4_d
+ N_XI61/XI15/NET34_XI61/XI15/MM4_g N_VDD_XI61/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI15/MM10 N_XI61/XI15/NET35_XI61/XI15/MM10_d
+ N_XI61/XI15/NET36_XI61/XI15/MM10_g N_VDD_XI61/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI61/XI15/MM11 N_XI61/XI15/NET36_XI61/XI15/MM11_d
+ N_XI61/XI15/NET35_XI61/XI15/MM11_g N_VDD_XI61/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI0/MM2 N_XI62/XI0/NET34_XI62/XI0/MM2_d N_XI62/XI0/NET33_XI62/XI0/MM2_g
+ N_VSS_XI62/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI0/MM3 N_XI62/XI0/NET33_XI62/XI0/MM3_d N_WL<120>_XI62/XI0/MM3_g
+ N_BLN<15>_XI62/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI0/MM0 N_XI62/XI0/NET34_XI62/XI0/MM0_d N_WL<120>_XI62/XI0/MM0_g
+ N_BL<15>_XI62/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI0/MM1 N_XI62/XI0/NET33_XI62/XI0/MM1_d N_XI62/XI0/NET34_XI62/XI0/MM1_g
+ N_VSS_XI62/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI0/MM9 N_XI62/XI0/NET36_XI62/XI0/MM9_d N_WL<121>_XI62/XI0/MM9_g
+ N_BL<15>_XI62/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI0/MM6 N_XI62/XI0/NET35_XI62/XI0/MM6_d N_XI62/XI0/NET36_XI62/XI0/MM6_g
+ N_VSS_XI62/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI0/MM7 N_XI62/XI0/NET36_XI62/XI0/MM7_d N_XI62/XI0/NET35_XI62/XI0/MM7_g
+ N_VSS_XI62/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI0/MM8 N_XI62/XI0/NET35_XI62/XI0/MM8_d N_WL<121>_XI62/XI0/MM8_g
+ N_BLN<15>_XI62/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI0/MM5 N_XI62/XI0/NET34_XI62/XI0/MM5_d N_XI62/XI0/NET33_XI62/XI0/MM5_g
+ N_VDD_XI62/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI0/MM4 N_XI62/XI0/NET33_XI62/XI0/MM4_d N_XI62/XI0/NET34_XI62/XI0/MM4_g
+ N_VDD_XI62/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI0/MM10 N_XI62/XI0/NET35_XI62/XI0/MM10_d N_XI62/XI0/NET36_XI62/XI0/MM10_g
+ N_VDD_XI62/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI0/MM11 N_XI62/XI0/NET36_XI62/XI0/MM11_d N_XI62/XI0/NET35_XI62/XI0/MM11_g
+ N_VDD_XI62/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI1/MM2 N_XI62/XI1/NET34_XI62/XI1/MM2_d N_XI62/XI1/NET33_XI62/XI1/MM2_g
+ N_VSS_XI62/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI1/MM3 N_XI62/XI1/NET33_XI62/XI1/MM3_d N_WL<120>_XI62/XI1/MM3_g
+ N_BLN<14>_XI62/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI1/MM0 N_XI62/XI1/NET34_XI62/XI1/MM0_d N_WL<120>_XI62/XI1/MM0_g
+ N_BL<14>_XI62/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI1/MM1 N_XI62/XI1/NET33_XI62/XI1/MM1_d N_XI62/XI1/NET34_XI62/XI1/MM1_g
+ N_VSS_XI62/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI1/MM9 N_XI62/XI1/NET36_XI62/XI1/MM9_d N_WL<121>_XI62/XI1/MM9_g
+ N_BL<14>_XI62/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI1/MM6 N_XI62/XI1/NET35_XI62/XI1/MM6_d N_XI62/XI1/NET36_XI62/XI1/MM6_g
+ N_VSS_XI62/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI1/MM7 N_XI62/XI1/NET36_XI62/XI1/MM7_d N_XI62/XI1/NET35_XI62/XI1/MM7_g
+ N_VSS_XI62/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI1/MM8 N_XI62/XI1/NET35_XI62/XI1/MM8_d N_WL<121>_XI62/XI1/MM8_g
+ N_BLN<14>_XI62/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI1/MM5 N_XI62/XI1/NET34_XI62/XI1/MM5_d N_XI62/XI1/NET33_XI62/XI1/MM5_g
+ N_VDD_XI62/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI1/MM4 N_XI62/XI1/NET33_XI62/XI1/MM4_d N_XI62/XI1/NET34_XI62/XI1/MM4_g
+ N_VDD_XI62/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI1/MM10 N_XI62/XI1/NET35_XI62/XI1/MM10_d N_XI62/XI1/NET36_XI62/XI1/MM10_g
+ N_VDD_XI62/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI1/MM11 N_XI62/XI1/NET36_XI62/XI1/MM11_d N_XI62/XI1/NET35_XI62/XI1/MM11_g
+ N_VDD_XI62/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI2/MM2 N_XI62/XI2/NET34_XI62/XI2/MM2_d N_XI62/XI2/NET33_XI62/XI2/MM2_g
+ N_VSS_XI62/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI2/MM3 N_XI62/XI2/NET33_XI62/XI2/MM3_d N_WL<120>_XI62/XI2/MM3_g
+ N_BLN<13>_XI62/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI2/MM0 N_XI62/XI2/NET34_XI62/XI2/MM0_d N_WL<120>_XI62/XI2/MM0_g
+ N_BL<13>_XI62/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI2/MM1 N_XI62/XI2/NET33_XI62/XI2/MM1_d N_XI62/XI2/NET34_XI62/XI2/MM1_g
+ N_VSS_XI62/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI2/MM9 N_XI62/XI2/NET36_XI62/XI2/MM9_d N_WL<121>_XI62/XI2/MM9_g
+ N_BL<13>_XI62/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI2/MM6 N_XI62/XI2/NET35_XI62/XI2/MM6_d N_XI62/XI2/NET36_XI62/XI2/MM6_g
+ N_VSS_XI62/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI2/MM7 N_XI62/XI2/NET36_XI62/XI2/MM7_d N_XI62/XI2/NET35_XI62/XI2/MM7_g
+ N_VSS_XI62/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI2/MM8 N_XI62/XI2/NET35_XI62/XI2/MM8_d N_WL<121>_XI62/XI2/MM8_g
+ N_BLN<13>_XI62/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI2/MM5 N_XI62/XI2/NET34_XI62/XI2/MM5_d N_XI62/XI2/NET33_XI62/XI2/MM5_g
+ N_VDD_XI62/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI2/MM4 N_XI62/XI2/NET33_XI62/XI2/MM4_d N_XI62/XI2/NET34_XI62/XI2/MM4_g
+ N_VDD_XI62/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI2/MM10 N_XI62/XI2/NET35_XI62/XI2/MM10_d N_XI62/XI2/NET36_XI62/XI2/MM10_g
+ N_VDD_XI62/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI2/MM11 N_XI62/XI2/NET36_XI62/XI2/MM11_d N_XI62/XI2/NET35_XI62/XI2/MM11_g
+ N_VDD_XI62/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI3/MM2 N_XI62/XI3/NET34_XI62/XI3/MM2_d N_XI62/XI3/NET33_XI62/XI3/MM2_g
+ N_VSS_XI62/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI3/MM3 N_XI62/XI3/NET33_XI62/XI3/MM3_d N_WL<120>_XI62/XI3/MM3_g
+ N_BLN<12>_XI62/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI3/MM0 N_XI62/XI3/NET34_XI62/XI3/MM0_d N_WL<120>_XI62/XI3/MM0_g
+ N_BL<12>_XI62/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI3/MM1 N_XI62/XI3/NET33_XI62/XI3/MM1_d N_XI62/XI3/NET34_XI62/XI3/MM1_g
+ N_VSS_XI62/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI3/MM9 N_XI62/XI3/NET36_XI62/XI3/MM9_d N_WL<121>_XI62/XI3/MM9_g
+ N_BL<12>_XI62/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI3/MM6 N_XI62/XI3/NET35_XI62/XI3/MM6_d N_XI62/XI3/NET36_XI62/XI3/MM6_g
+ N_VSS_XI62/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI3/MM7 N_XI62/XI3/NET36_XI62/XI3/MM7_d N_XI62/XI3/NET35_XI62/XI3/MM7_g
+ N_VSS_XI62/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI3/MM8 N_XI62/XI3/NET35_XI62/XI3/MM8_d N_WL<121>_XI62/XI3/MM8_g
+ N_BLN<12>_XI62/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI3/MM5 N_XI62/XI3/NET34_XI62/XI3/MM5_d N_XI62/XI3/NET33_XI62/XI3/MM5_g
+ N_VDD_XI62/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI3/MM4 N_XI62/XI3/NET33_XI62/XI3/MM4_d N_XI62/XI3/NET34_XI62/XI3/MM4_g
+ N_VDD_XI62/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI3/MM10 N_XI62/XI3/NET35_XI62/XI3/MM10_d N_XI62/XI3/NET36_XI62/XI3/MM10_g
+ N_VDD_XI62/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI3/MM11 N_XI62/XI3/NET36_XI62/XI3/MM11_d N_XI62/XI3/NET35_XI62/XI3/MM11_g
+ N_VDD_XI62/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI4/MM2 N_XI62/XI4/NET34_XI62/XI4/MM2_d N_XI62/XI4/NET33_XI62/XI4/MM2_g
+ N_VSS_XI62/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI4/MM3 N_XI62/XI4/NET33_XI62/XI4/MM3_d N_WL<120>_XI62/XI4/MM3_g
+ N_BLN<11>_XI62/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI4/MM0 N_XI62/XI4/NET34_XI62/XI4/MM0_d N_WL<120>_XI62/XI4/MM0_g
+ N_BL<11>_XI62/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI4/MM1 N_XI62/XI4/NET33_XI62/XI4/MM1_d N_XI62/XI4/NET34_XI62/XI4/MM1_g
+ N_VSS_XI62/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI4/MM9 N_XI62/XI4/NET36_XI62/XI4/MM9_d N_WL<121>_XI62/XI4/MM9_g
+ N_BL<11>_XI62/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI4/MM6 N_XI62/XI4/NET35_XI62/XI4/MM6_d N_XI62/XI4/NET36_XI62/XI4/MM6_g
+ N_VSS_XI62/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI4/MM7 N_XI62/XI4/NET36_XI62/XI4/MM7_d N_XI62/XI4/NET35_XI62/XI4/MM7_g
+ N_VSS_XI62/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI4/MM8 N_XI62/XI4/NET35_XI62/XI4/MM8_d N_WL<121>_XI62/XI4/MM8_g
+ N_BLN<11>_XI62/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI4/MM5 N_XI62/XI4/NET34_XI62/XI4/MM5_d N_XI62/XI4/NET33_XI62/XI4/MM5_g
+ N_VDD_XI62/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI4/MM4 N_XI62/XI4/NET33_XI62/XI4/MM4_d N_XI62/XI4/NET34_XI62/XI4/MM4_g
+ N_VDD_XI62/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI4/MM10 N_XI62/XI4/NET35_XI62/XI4/MM10_d N_XI62/XI4/NET36_XI62/XI4/MM10_g
+ N_VDD_XI62/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI4/MM11 N_XI62/XI4/NET36_XI62/XI4/MM11_d N_XI62/XI4/NET35_XI62/XI4/MM11_g
+ N_VDD_XI62/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI5/MM2 N_XI62/XI5/NET34_XI62/XI5/MM2_d N_XI62/XI5/NET33_XI62/XI5/MM2_g
+ N_VSS_XI62/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI5/MM3 N_XI62/XI5/NET33_XI62/XI5/MM3_d N_WL<120>_XI62/XI5/MM3_g
+ N_BLN<10>_XI62/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI5/MM0 N_XI62/XI5/NET34_XI62/XI5/MM0_d N_WL<120>_XI62/XI5/MM0_g
+ N_BL<10>_XI62/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI5/MM1 N_XI62/XI5/NET33_XI62/XI5/MM1_d N_XI62/XI5/NET34_XI62/XI5/MM1_g
+ N_VSS_XI62/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI5/MM9 N_XI62/XI5/NET36_XI62/XI5/MM9_d N_WL<121>_XI62/XI5/MM9_g
+ N_BL<10>_XI62/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI5/MM6 N_XI62/XI5/NET35_XI62/XI5/MM6_d N_XI62/XI5/NET36_XI62/XI5/MM6_g
+ N_VSS_XI62/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI5/MM7 N_XI62/XI5/NET36_XI62/XI5/MM7_d N_XI62/XI5/NET35_XI62/XI5/MM7_g
+ N_VSS_XI62/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI5/MM8 N_XI62/XI5/NET35_XI62/XI5/MM8_d N_WL<121>_XI62/XI5/MM8_g
+ N_BLN<10>_XI62/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI5/MM5 N_XI62/XI5/NET34_XI62/XI5/MM5_d N_XI62/XI5/NET33_XI62/XI5/MM5_g
+ N_VDD_XI62/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI5/MM4 N_XI62/XI5/NET33_XI62/XI5/MM4_d N_XI62/XI5/NET34_XI62/XI5/MM4_g
+ N_VDD_XI62/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI5/MM10 N_XI62/XI5/NET35_XI62/XI5/MM10_d N_XI62/XI5/NET36_XI62/XI5/MM10_g
+ N_VDD_XI62/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI5/MM11 N_XI62/XI5/NET36_XI62/XI5/MM11_d N_XI62/XI5/NET35_XI62/XI5/MM11_g
+ N_VDD_XI62/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI6/MM2 N_XI62/XI6/NET34_XI62/XI6/MM2_d N_XI62/XI6/NET33_XI62/XI6/MM2_g
+ N_VSS_XI62/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM3 N_XI62/XI6/NET33_XI62/XI6/MM3_d N_WL<120>_XI62/XI6/MM3_g
+ N_BLN<9>_XI62/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM0 N_XI62/XI6/NET34_XI62/XI6/MM0_d N_WL<120>_XI62/XI6/MM0_g
+ N_BL<9>_XI62/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM1 N_XI62/XI6/NET33_XI62/XI6/MM1_d N_XI62/XI6/NET34_XI62/XI6/MM1_g
+ N_VSS_XI62/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM9 N_XI62/XI6/NET36_XI62/XI6/MM9_d N_WL<121>_XI62/XI6/MM9_g
+ N_BL<9>_XI62/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM6 N_XI62/XI6/NET35_XI62/XI6/MM6_d N_XI62/XI6/NET36_XI62/XI6/MM6_g
+ N_VSS_XI62/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM7 N_XI62/XI6/NET36_XI62/XI6/MM7_d N_XI62/XI6/NET35_XI62/XI6/MM7_g
+ N_VSS_XI62/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM8 N_XI62/XI6/NET35_XI62/XI6/MM8_d N_WL<121>_XI62/XI6/MM8_g
+ N_BLN<9>_XI62/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI6/MM5 N_XI62/XI6/NET34_XI62/XI6/MM5_d N_XI62/XI6/NET33_XI62/XI6/MM5_g
+ N_VDD_XI62/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI6/MM4 N_XI62/XI6/NET33_XI62/XI6/MM4_d N_XI62/XI6/NET34_XI62/XI6/MM4_g
+ N_VDD_XI62/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI6/MM10 N_XI62/XI6/NET35_XI62/XI6/MM10_d N_XI62/XI6/NET36_XI62/XI6/MM10_g
+ N_VDD_XI62/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI6/MM11 N_XI62/XI6/NET36_XI62/XI6/MM11_d N_XI62/XI6/NET35_XI62/XI6/MM11_g
+ N_VDD_XI62/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI7/MM2 N_XI62/XI7/NET34_XI62/XI7/MM2_d N_XI62/XI7/NET33_XI62/XI7/MM2_g
+ N_VSS_XI62/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM3 N_XI62/XI7/NET33_XI62/XI7/MM3_d N_WL<120>_XI62/XI7/MM3_g
+ N_BLN<8>_XI62/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM0 N_XI62/XI7/NET34_XI62/XI7/MM0_d N_WL<120>_XI62/XI7/MM0_g
+ N_BL<8>_XI62/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM1 N_XI62/XI7/NET33_XI62/XI7/MM1_d N_XI62/XI7/NET34_XI62/XI7/MM1_g
+ N_VSS_XI62/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM9 N_XI62/XI7/NET36_XI62/XI7/MM9_d N_WL<121>_XI62/XI7/MM9_g
+ N_BL<8>_XI62/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM6 N_XI62/XI7/NET35_XI62/XI7/MM6_d N_XI62/XI7/NET36_XI62/XI7/MM6_g
+ N_VSS_XI62/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM7 N_XI62/XI7/NET36_XI62/XI7/MM7_d N_XI62/XI7/NET35_XI62/XI7/MM7_g
+ N_VSS_XI62/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM8 N_XI62/XI7/NET35_XI62/XI7/MM8_d N_WL<121>_XI62/XI7/MM8_g
+ N_BLN<8>_XI62/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI7/MM5 N_XI62/XI7/NET34_XI62/XI7/MM5_d N_XI62/XI7/NET33_XI62/XI7/MM5_g
+ N_VDD_XI62/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI7/MM4 N_XI62/XI7/NET33_XI62/XI7/MM4_d N_XI62/XI7/NET34_XI62/XI7/MM4_g
+ N_VDD_XI62/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI7/MM10 N_XI62/XI7/NET35_XI62/XI7/MM10_d N_XI62/XI7/NET36_XI62/XI7/MM10_g
+ N_VDD_XI62/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI7/MM11 N_XI62/XI7/NET36_XI62/XI7/MM11_d N_XI62/XI7/NET35_XI62/XI7/MM11_g
+ N_VDD_XI62/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI8/MM2 N_XI62/XI8/NET34_XI62/XI8/MM2_d N_XI62/XI8/NET33_XI62/XI8/MM2_g
+ N_VSS_XI62/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM3 N_XI62/XI8/NET33_XI62/XI8/MM3_d N_WL<120>_XI62/XI8/MM3_g
+ N_BLN<7>_XI62/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM0 N_XI62/XI8/NET34_XI62/XI8/MM0_d N_WL<120>_XI62/XI8/MM0_g
+ N_BL<7>_XI62/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM1 N_XI62/XI8/NET33_XI62/XI8/MM1_d N_XI62/XI8/NET34_XI62/XI8/MM1_g
+ N_VSS_XI62/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM9 N_XI62/XI8/NET36_XI62/XI8/MM9_d N_WL<121>_XI62/XI8/MM9_g
+ N_BL<7>_XI62/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM6 N_XI62/XI8/NET35_XI62/XI8/MM6_d N_XI62/XI8/NET36_XI62/XI8/MM6_g
+ N_VSS_XI62/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM7 N_XI62/XI8/NET36_XI62/XI8/MM7_d N_XI62/XI8/NET35_XI62/XI8/MM7_g
+ N_VSS_XI62/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM8 N_XI62/XI8/NET35_XI62/XI8/MM8_d N_WL<121>_XI62/XI8/MM8_g
+ N_BLN<7>_XI62/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI8/MM5 N_XI62/XI8/NET34_XI62/XI8/MM5_d N_XI62/XI8/NET33_XI62/XI8/MM5_g
+ N_VDD_XI62/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI8/MM4 N_XI62/XI8/NET33_XI62/XI8/MM4_d N_XI62/XI8/NET34_XI62/XI8/MM4_g
+ N_VDD_XI62/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI8/MM10 N_XI62/XI8/NET35_XI62/XI8/MM10_d N_XI62/XI8/NET36_XI62/XI8/MM10_g
+ N_VDD_XI62/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI8/MM11 N_XI62/XI8/NET36_XI62/XI8/MM11_d N_XI62/XI8/NET35_XI62/XI8/MM11_g
+ N_VDD_XI62/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI9/MM2 N_XI62/XI9/NET34_XI62/XI9/MM2_d N_XI62/XI9/NET33_XI62/XI9/MM2_g
+ N_VSS_XI62/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM3 N_XI62/XI9/NET33_XI62/XI9/MM3_d N_WL<120>_XI62/XI9/MM3_g
+ N_BLN<6>_XI62/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM0 N_XI62/XI9/NET34_XI62/XI9/MM0_d N_WL<120>_XI62/XI9/MM0_g
+ N_BL<6>_XI62/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM1 N_XI62/XI9/NET33_XI62/XI9/MM1_d N_XI62/XI9/NET34_XI62/XI9/MM1_g
+ N_VSS_XI62/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM9 N_XI62/XI9/NET36_XI62/XI9/MM9_d N_WL<121>_XI62/XI9/MM9_g
+ N_BL<6>_XI62/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM6 N_XI62/XI9/NET35_XI62/XI9/MM6_d N_XI62/XI9/NET36_XI62/XI9/MM6_g
+ N_VSS_XI62/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM7 N_XI62/XI9/NET36_XI62/XI9/MM7_d N_XI62/XI9/NET35_XI62/XI9/MM7_g
+ N_VSS_XI62/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM8 N_XI62/XI9/NET35_XI62/XI9/MM8_d N_WL<121>_XI62/XI9/MM8_g
+ N_BLN<6>_XI62/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI9/MM5 N_XI62/XI9/NET34_XI62/XI9/MM5_d N_XI62/XI9/NET33_XI62/XI9/MM5_g
+ N_VDD_XI62/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI9/MM4 N_XI62/XI9/NET33_XI62/XI9/MM4_d N_XI62/XI9/NET34_XI62/XI9/MM4_g
+ N_VDD_XI62/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI9/MM10 N_XI62/XI9/NET35_XI62/XI9/MM10_d N_XI62/XI9/NET36_XI62/XI9/MM10_g
+ N_VDD_XI62/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI9/MM11 N_XI62/XI9/NET36_XI62/XI9/MM11_d N_XI62/XI9/NET35_XI62/XI9/MM11_g
+ N_VDD_XI62/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI10/MM2 N_XI62/XI10/NET34_XI62/XI10/MM2_d
+ N_XI62/XI10/NET33_XI62/XI10/MM2_g N_VSS_XI62/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI10/MM3 N_XI62/XI10/NET33_XI62/XI10/MM3_d N_WL<120>_XI62/XI10/MM3_g
+ N_BLN<5>_XI62/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI10/MM0 N_XI62/XI10/NET34_XI62/XI10/MM0_d N_WL<120>_XI62/XI10/MM0_g
+ N_BL<5>_XI62/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI10/MM1 N_XI62/XI10/NET33_XI62/XI10/MM1_d
+ N_XI62/XI10/NET34_XI62/XI10/MM1_g N_VSS_XI62/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI10/MM9 N_XI62/XI10/NET36_XI62/XI10/MM9_d N_WL<121>_XI62/XI10/MM9_g
+ N_BL<5>_XI62/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI10/MM6 N_XI62/XI10/NET35_XI62/XI10/MM6_d
+ N_XI62/XI10/NET36_XI62/XI10/MM6_g N_VSS_XI62/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI10/MM7 N_XI62/XI10/NET36_XI62/XI10/MM7_d
+ N_XI62/XI10/NET35_XI62/XI10/MM7_g N_VSS_XI62/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI10/MM8 N_XI62/XI10/NET35_XI62/XI10/MM8_d N_WL<121>_XI62/XI10/MM8_g
+ N_BLN<5>_XI62/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI10/MM5 N_XI62/XI10/NET34_XI62/XI10/MM5_d
+ N_XI62/XI10/NET33_XI62/XI10/MM5_g N_VDD_XI62/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI10/MM4 N_XI62/XI10/NET33_XI62/XI10/MM4_d
+ N_XI62/XI10/NET34_XI62/XI10/MM4_g N_VDD_XI62/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI10/MM10 N_XI62/XI10/NET35_XI62/XI10/MM10_d
+ N_XI62/XI10/NET36_XI62/XI10/MM10_g N_VDD_XI62/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI10/MM11 N_XI62/XI10/NET36_XI62/XI10/MM11_d
+ N_XI62/XI10/NET35_XI62/XI10/MM11_g N_VDD_XI62/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI11/MM2 N_XI62/XI11/NET34_XI62/XI11/MM2_d
+ N_XI62/XI11/NET33_XI62/XI11/MM2_g N_VSS_XI62/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI11/MM3 N_XI62/XI11/NET33_XI62/XI11/MM3_d N_WL<120>_XI62/XI11/MM3_g
+ N_BLN<4>_XI62/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI11/MM0 N_XI62/XI11/NET34_XI62/XI11/MM0_d N_WL<120>_XI62/XI11/MM0_g
+ N_BL<4>_XI62/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI11/MM1 N_XI62/XI11/NET33_XI62/XI11/MM1_d
+ N_XI62/XI11/NET34_XI62/XI11/MM1_g N_VSS_XI62/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI11/MM9 N_XI62/XI11/NET36_XI62/XI11/MM9_d N_WL<121>_XI62/XI11/MM9_g
+ N_BL<4>_XI62/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI11/MM6 N_XI62/XI11/NET35_XI62/XI11/MM6_d
+ N_XI62/XI11/NET36_XI62/XI11/MM6_g N_VSS_XI62/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI11/MM7 N_XI62/XI11/NET36_XI62/XI11/MM7_d
+ N_XI62/XI11/NET35_XI62/XI11/MM7_g N_VSS_XI62/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI11/MM8 N_XI62/XI11/NET35_XI62/XI11/MM8_d N_WL<121>_XI62/XI11/MM8_g
+ N_BLN<4>_XI62/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI11/MM5 N_XI62/XI11/NET34_XI62/XI11/MM5_d
+ N_XI62/XI11/NET33_XI62/XI11/MM5_g N_VDD_XI62/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI11/MM4 N_XI62/XI11/NET33_XI62/XI11/MM4_d
+ N_XI62/XI11/NET34_XI62/XI11/MM4_g N_VDD_XI62/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI11/MM10 N_XI62/XI11/NET35_XI62/XI11/MM10_d
+ N_XI62/XI11/NET36_XI62/XI11/MM10_g N_VDD_XI62/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI11/MM11 N_XI62/XI11/NET36_XI62/XI11/MM11_d
+ N_XI62/XI11/NET35_XI62/XI11/MM11_g N_VDD_XI62/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI12/MM2 N_XI62/XI12/NET34_XI62/XI12/MM2_d
+ N_XI62/XI12/NET33_XI62/XI12/MM2_g N_VSS_XI62/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI12/MM3 N_XI62/XI12/NET33_XI62/XI12/MM3_d N_WL<120>_XI62/XI12/MM3_g
+ N_BLN<3>_XI62/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI12/MM0 N_XI62/XI12/NET34_XI62/XI12/MM0_d N_WL<120>_XI62/XI12/MM0_g
+ N_BL<3>_XI62/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI12/MM1 N_XI62/XI12/NET33_XI62/XI12/MM1_d
+ N_XI62/XI12/NET34_XI62/XI12/MM1_g N_VSS_XI62/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI12/MM9 N_XI62/XI12/NET36_XI62/XI12/MM9_d N_WL<121>_XI62/XI12/MM9_g
+ N_BL<3>_XI62/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI12/MM6 N_XI62/XI12/NET35_XI62/XI12/MM6_d
+ N_XI62/XI12/NET36_XI62/XI12/MM6_g N_VSS_XI62/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI12/MM7 N_XI62/XI12/NET36_XI62/XI12/MM7_d
+ N_XI62/XI12/NET35_XI62/XI12/MM7_g N_VSS_XI62/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI12/MM8 N_XI62/XI12/NET35_XI62/XI12/MM8_d N_WL<121>_XI62/XI12/MM8_g
+ N_BLN<3>_XI62/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI12/MM5 N_XI62/XI12/NET34_XI62/XI12/MM5_d
+ N_XI62/XI12/NET33_XI62/XI12/MM5_g N_VDD_XI62/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI12/MM4 N_XI62/XI12/NET33_XI62/XI12/MM4_d
+ N_XI62/XI12/NET34_XI62/XI12/MM4_g N_VDD_XI62/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI12/MM10 N_XI62/XI12/NET35_XI62/XI12/MM10_d
+ N_XI62/XI12/NET36_XI62/XI12/MM10_g N_VDD_XI62/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI12/MM11 N_XI62/XI12/NET36_XI62/XI12/MM11_d
+ N_XI62/XI12/NET35_XI62/XI12/MM11_g N_VDD_XI62/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI13/MM2 N_XI62/XI13/NET34_XI62/XI13/MM2_d
+ N_XI62/XI13/NET33_XI62/XI13/MM2_g N_VSS_XI62/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI13/MM3 N_XI62/XI13/NET33_XI62/XI13/MM3_d N_WL<120>_XI62/XI13/MM3_g
+ N_BLN<2>_XI62/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI13/MM0 N_XI62/XI13/NET34_XI62/XI13/MM0_d N_WL<120>_XI62/XI13/MM0_g
+ N_BL<2>_XI62/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI13/MM1 N_XI62/XI13/NET33_XI62/XI13/MM1_d
+ N_XI62/XI13/NET34_XI62/XI13/MM1_g N_VSS_XI62/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI13/MM9 N_XI62/XI13/NET36_XI62/XI13/MM9_d N_WL<121>_XI62/XI13/MM9_g
+ N_BL<2>_XI62/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI13/MM6 N_XI62/XI13/NET35_XI62/XI13/MM6_d
+ N_XI62/XI13/NET36_XI62/XI13/MM6_g N_VSS_XI62/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI13/MM7 N_XI62/XI13/NET36_XI62/XI13/MM7_d
+ N_XI62/XI13/NET35_XI62/XI13/MM7_g N_VSS_XI62/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI13/MM8 N_XI62/XI13/NET35_XI62/XI13/MM8_d N_WL<121>_XI62/XI13/MM8_g
+ N_BLN<2>_XI62/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI13/MM5 N_XI62/XI13/NET34_XI62/XI13/MM5_d
+ N_XI62/XI13/NET33_XI62/XI13/MM5_g N_VDD_XI62/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI13/MM4 N_XI62/XI13/NET33_XI62/XI13/MM4_d
+ N_XI62/XI13/NET34_XI62/XI13/MM4_g N_VDD_XI62/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI13/MM10 N_XI62/XI13/NET35_XI62/XI13/MM10_d
+ N_XI62/XI13/NET36_XI62/XI13/MM10_g N_VDD_XI62/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI13/MM11 N_XI62/XI13/NET36_XI62/XI13/MM11_d
+ N_XI62/XI13/NET35_XI62/XI13/MM11_g N_VDD_XI62/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI14/MM2 N_XI62/XI14/NET34_XI62/XI14/MM2_d
+ N_XI62/XI14/NET33_XI62/XI14/MM2_g N_VSS_XI62/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI14/MM3 N_XI62/XI14/NET33_XI62/XI14/MM3_d N_WL<120>_XI62/XI14/MM3_g
+ N_BLN<1>_XI62/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI14/MM0 N_XI62/XI14/NET34_XI62/XI14/MM0_d N_WL<120>_XI62/XI14/MM0_g
+ N_BL<1>_XI62/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI14/MM1 N_XI62/XI14/NET33_XI62/XI14/MM1_d
+ N_XI62/XI14/NET34_XI62/XI14/MM1_g N_VSS_XI62/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI14/MM9 N_XI62/XI14/NET36_XI62/XI14/MM9_d N_WL<121>_XI62/XI14/MM9_g
+ N_BL<1>_XI62/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI14/MM6 N_XI62/XI14/NET35_XI62/XI14/MM6_d
+ N_XI62/XI14/NET36_XI62/XI14/MM6_g N_VSS_XI62/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI14/MM7 N_XI62/XI14/NET36_XI62/XI14/MM7_d
+ N_XI62/XI14/NET35_XI62/XI14/MM7_g N_VSS_XI62/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI14/MM8 N_XI62/XI14/NET35_XI62/XI14/MM8_d N_WL<121>_XI62/XI14/MM8_g
+ N_BLN<1>_XI62/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI14/MM5 N_XI62/XI14/NET34_XI62/XI14/MM5_d
+ N_XI62/XI14/NET33_XI62/XI14/MM5_g N_VDD_XI62/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI14/MM4 N_XI62/XI14/NET33_XI62/XI14/MM4_d
+ N_XI62/XI14/NET34_XI62/XI14/MM4_g N_VDD_XI62/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI14/MM10 N_XI62/XI14/NET35_XI62/XI14/MM10_d
+ N_XI62/XI14/NET36_XI62/XI14/MM10_g N_VDD_XI62/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI14/MM11 N_XI62/XI14/NET36_XI62/XI14/MM11_d
+ N_XI62/XI14/NET35_XI62/XI14/MM11_g N_VDD_XI62/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI15/MM2 N_XI62/XI15/NET34_XI62/XI15/MM2_d
+ N_XI62/XI15/NET33_XI62/XI15/MM2_g N_VSS_XI62/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI15/MM3 N_XI62/XI15/NET33_XI62/XI15/MM3_d N_WL<120>_XI62/XI15/MM3_g
+ N_BLN<0>_XI62/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI15/MM0 N_XI62/XI15/NET34_XI62/XI15/MM0_d N_WL<120>_XI62/XI15/MM0_g
+ N_BL<0>_XI62/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI15/MM1 N_XI62/XI15/NET33_XI62/XI15/MM1_d
+ N_XI62/XI15/NET34_XI62/XI15/MM1_g N_VSS_XI62/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI15/MM9 N_XI62/XI15/NET36_XI62/XI15/MM9_d N_WL<121>_XI62/XI15/MM9_g
+ N_BL<0>_XI62/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI15/MM6 N_XI62/XI15/NET35_XI62/XI15/MM6_d
+ N_XI62/XI15/NET36_XI62/XI15/MM6_g N_VSS_XI62/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI15/MM7 N_XI62/XI15/NET36_XI62/XI15/MM7_d
+ N_XI62/XI15/NET35_XI62/XI15/MM7_g N_VSS_XI62/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI62/XI15/MM8 N_XI62/XI15/NET35_XI62/XI15/MM8_d N_WL<121>_XI62/XI15/MM8_g
+ N_BLN<0>_XI62/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI62/XI15/MM5 N_XI62/XI15/NET34_XI62/XI15/MM5_d
+ N_XI62/XI15/NET33_XI62/XI15/MM5_g N_VDD_XI62/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI15/MM4 N_XI62/XI15/NET33_XI62/XI15/MM4_d
+ N_XI62/XI15/NET34_XI62/XI15/MM4_g N_VDD_XI62/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI15/MM10 N_XI62/XI15/NET35_XI62/XI15/MM10_d
+ N_XI62/XI15/NET36_XI62/XI15/MM10_g N_VDD_XI62/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI62/XI15/MM11 N_XI62/XI15/NET36_XI62/XI15/MM11_d
+ N_XI62/XI15/NET35_XI62/XI15/MM11_g N_VDD_XI62/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI0/MM2 N_XI63/XI0/NET34_XI63/XI0/MM2_d N_XI63/XI0/NET33_XI63/XI0/MM2_g
+ N_VSS_XI63/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI0/MM3 N_XI63/XI0/NET33_XI63/XI0/MM3_d N_WL<122>_XI63/XI0/MM3_g
+ N_BLN<15>_XI63/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI0/MM0 N_XI63/XI0/NET34_XI63/XI0/MM0_d N_WL<122>_XI63/XI0/MM0_g
+ N_BL<15>_XI63/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI0/MM1 N_XI63/XI0/NET33_XI63/XI0/MM1_d N_XI63/XI0/NET34_XI63/XI0/MM1_g
+ N_VSS_XI63/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI0/MM9 N_XI63/XI0/NET36_XI63/XI0/MM9_d N_WL<123>_XI63/XI0/MM9_g
+ N_BL<15>_XI63/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI0/MM6 N_XI63/XI0/NET35_XI63/XI0/MM6_d N_XI63/XI0/NET36_XI63/XI0/MM6_g
+ N_VSS_XI63/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI0/MM7 N_XI63/XI0/NET36_XI63/XI0/MM7_d N_XI63/XI0/NET35_XI63/XI0/MM7_g
+ N_VSS_XI63/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI0/MM8 N_XI63/XI0/NET35_XI63/XI0/MM8_d N_WL<123>_XI63/XI0/MM8_g
+ N_BLN<15>_XI63/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI0/MM5 N_XI63/XI0/NET34_XI63/XI0/MM5_d N_XI63/XI0/NET33_XI63/XI0/MM5_g
+ N_VDD_XI63/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI0/MM4 N_XI63/XI0/NET33_XI63/XI0/MM4_d N_XI63/XI0/NET34_XI63/XI0/MM4_g
+ N_VDD_XI63/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI0/MM10 N_XI63/XI0/NET35_XI63/XI0/MM10_d N_XI63/XI0/NET36_XI63/XI0/MM10_g
+ N_VDD_XI63/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI0/MM11 N_XI63/XI0/NET36_XI63/XI0/MM11_d N_XI63/XI0/NET35_XI63/XI0/MM11_g
+ N_VDD_XI63/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI1/MM2 N_XI63/XI1/NET34_XI63/XI1/MM2_d N_XI63/XI1/NET33_XI63/XI1/MM2_g
+ N_VSS_XI63/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI1/MM3 N_XI63/XI1/NET33_XI63/XI1/MM3_d N_WL<122>_XI63/XI1/MM3_g
+ N_BLN<14>_XI63/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI1/MM0 N_XI63/XI1/NET34_XI63/XI1/MM0_d N_WL<122>_XI63/XI1/MM0_g
+ N_BL<14>_XI63/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI1/MM1 N_XI63/XI1/NET33_XI63/XI1/MM1_d N_XI63/XI1/NET34_XI63/XI1/MM1_g
+ N_VSS_XI63/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI1/MM9 N_XI63/XI1/NET36_XI63/XI1/MM9_d N_WL<123>_XI63/XI1/MM9_g
+ N_BL<14>_XI63/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI1/MM6 N_XI63/XI1/NET35_XI63/XI1/MM6_d N_XI63/XI1/NET36_XI63/XI1/MM6_g
+ N_VSS_XI63/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI1/MM7 N_XI63/XI1/NET36_XI63/XI1/MM7_d N_XI63/XI1/NET35_XI63/XI1/MM7_g
+ N_VSS_XI63/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI1/MM8 N_XI63/XI1/NET35_XI63/XI1/MM8_d N_WL<123>_XI63/XI1/MM8_g
+ N_BLN<14>_XI63/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI1/MM5 N_XI63/XI1/NET34_XI63/XI1/MM5_d N_XI63/XI1/NET33_XI63/XI1/MM5_g
+ N_VDD_XI63/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI1/MM4 N_XI63/XI1/NET33_XI63/XI1/MM4_d N_XI63/XI1/NET34_XI63/XI1/MM4_g
+ N_VDD_XI63/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI1/MM10 N_XI63/XI1/NET35_XI63/XI1/MM10_d N_XI63/XI1/NET36_XI63/XI1/MM10_g
+ N_VDD_XI63/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI1/MM11 N_XI63/XI1/NET36_XI63/XI1/MM11_d N_XI63/XI1/NET35_XI63/XI1/MM11_g
+ N_VDD_XI63/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI2/MM2 N_XI63/XI2/NET34_XI63/XI2/MM2_d N_XI63/XI2/NET33_XI63/XI2/MM2_g
+ N_VSS_XI63/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI2/MM3 N_XI63/XI2/NET33_XI63/XI2/MM3_d N_WL<122>_XI63/XI2/MM3_g
+ N_BLN<13>_XI63/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI2/MM0 N_XI63/XI2/NET34_XI63/XI2/MM0_d N_WL<122>_XI63/XI2/MM0_g
+ N_BL<13>_XI63/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI2/MM1 N_XI63/XI2/NET33_XI63/XI2/MM1_d N_XI63/XI2/NET34_XI63/XI2/MM1_g
+ N_VSS_XI63/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI2/MM9 N_XI63/XI2/NET36_XI63/XI2/MM9_d N_WL<123>_XI63/XI2/MM9_g
+ N_BL<13>_XI63/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI2/MM6 N_XI63/XI2/NET35_XI63/XI2/MM6_d N_XI63/XI2/NET36_XI63/XI2/MM6_g
+ N_VSS_XI63/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI2/MM7 N_XI63/XI2/NET36_XI63/XI2/MM7_d N_XI63/XI2/NET35_XI63/XI2/MM7_g
+ N_VSS_XI63/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI2/MM8 N_XI63/XI2/NET35_XI63/XI2/MM8_d N_WL<123>_XI63/XI2/MM8_g
+ N_BLN<13>_XI63/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI2/MM5 N_XI63/XI2/NET34_XI63/XI2/MM5_d N_XI63/XI2/NET33_XI63/XI2/MM5_g
+ N_VDD_XI63/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI2/MM4 N_XI63/XI2/NET33_XI63/XI2/MM4_d N_XI63/XI2/NET34_XI63/XI2/MM4_g
+ N_VDD_XI63/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI2/MM10 N_XI63/XI2/NET35_XI63/XI2/MM10_d N_XI63/XI2/NET36_XI63/XI2/MM10_g
+ N_VDD_XI63/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI2/MM11 N_XI63/XI2/NET36_XI63/XI2/MM11_d N_XI63/XI2/NET35_XI63/XI2/MM11_g
+ N_VDD_XI63/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI3/MM2 N_XI63/XI3/NET34_XI63/XI3/MM2_d N_XI63/XI3/NET33_XI63/XI3/MM2_g
+ N_VSS_XI63/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI3/MM3 N_XI63/XI3/NET33_XI63/XI3/MM3_d N_WL<122>_XI63/XI3/MM3_g
+ N_BLN<12>_XI63/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI3/MM0 N_XI63/XI3/NET34_XI63/XI3/MM0_d N_WL<122>_XI63/XI3/MM0_g
+ N_BL<12>_XI63/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI3/MM1 N_XI63/XI3/NET33_XI63/XI3/MM1_d N_XI63/XI3/NET34_XI63/XI3/MM1_g
+ N_VSS_XI63/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI3/MM9 N_XI63/XI3/NET36_XI63/XI3/MM9_d N_WL<123>_XI63/XI3/MM9_g
+ N_BL<12>_XI63/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI3/MM6 N_XI63/XI3/NET35_XI63/XI3/MM6_d N_XI63/XI3/NET36_XI63/XI3/MM6_g
+ N_VSS_XI63/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI3/MM7 N_XI63/XI3/NET36_XI63/XI3/MM7_d N_XI63/XI3/NET35_XI63/XI3/MM7_g
+ N_VSS_XI63/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI3/MM8 N_XI63/XI3/NET35_XI63/XI3/MM8_d N_WL<123>_XI63/XI3/MM8_g
+ N_BLN<12>_XI63/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI3/MM5 N_XI63/XI3/NET34_XI63/XI3/MM5_d N_XI63/XI3/NET33_XI63/XI3/MM5_g
+ N_VDD_XI63/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI3/MM4 N_XI63/XI3/NET33_XI63/XI3/MM4_d N_XI63/XI3/NET34_XI63/XI3/MM4_g
+ N_VDD_XI63/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI3/MM10 N_XI63/XI3/NET35_XI63/XI3/MM10_d N_XI63/XI3/NET36_XI63/XI3/MM10_g
+ N_VDD_XI63/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI3/MM11 N_XI63/XI3/NET36_XI63/XI3/MM11_d N_XI63/XI3/NET35_XI63/XI3/MM11_g
+ N_VDD_XI63/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI4/MM2 N_XI63/XI4/NET34_XI63/XI4/MM2_d N_XI63/XI4/NET33_XI63/XI4/MM2_g
+ N_VSS_XI63/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI4/MM3 N_XI63/XI4/NET33_XI63/XI4/MM3_d N_WL<122>_XI63/XI4/MM3_g
+ N_BLN<11>_XI63/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI4/MM0 N_XI63/XI4/NET34_XI63/XI4/MM0_d N_WL<122>_XI63/XI4/MM0_g
+ N_BL<11>_XI63/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI4/MM1 N_XI63/XI4/NET33_XI63/XI4/MM1_d N_XI63/XI4/NET34_XI63/XI4/MM1_g
+ N_VSS_XI63/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI4/MM9 N_XI63/XI4/NET36_XI63/XI4/MM9_d N_WL<123>_XI63/XI4/MM9_g
+ N_BL<11>_XI63/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI4/MM6 N_XI63/XI4/NET35_XI63/XI4/MM6_d N_XI63/XI4/NET36_XI63/XI4/MM6_g
+ N_VSS_XI63/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI4/MM7 N_XI63/XI4/NET36_XI63/XI4/MM7_d N_XI63/XI4/NET35_XI63/XI4/MM7_g
+ N_VSS_XI63/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI4/MM8 N_XI63/XI4/NET35_XI63/XI4/MM8_d N_WL<123>_XI63/XI4/MM8_g
+ N_BLN<11>_XI63/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI4/MM5 N_XI63/XI4/NET34_XI63/XI4/MM5_d N_XI63/XI4/NET33_XI63/XI4/MM5_g
+ N_VDD_XI63/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI4/MM4 N_XI63/XI4/NET33_XI63/XI4/MM4_d N_XI63/XI4/NET34_XI63/XI4/MM4_g
+ N_VDD_XI63/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI4/MM10 N_XI63/XI4/NET35_XI63/XI4/MM10_d N_XI63/XI4/NET36_XI63/XI4/MM10_g
+ N_VDD_XI63/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI4/MM11 N_XI63/XI4/NET36_XI63/XI4/MM11_d N_XI63/XI4/NET35_XI63/XI4/MM11_g
+ N_VDD_XI63/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI5/MM2 N_XI63/XI5/NET34_XI63/XI5/MM2_d N_XI63/XI5/NET33_XI63/XI5/MM2_g
+ N_VSS_XI63/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI5/MM3 N_XI63/XI5/NET33_XI63/XI5/MM3_d N_WL<122>_XI63/XI5/MM3_g
+ N_BLN<10>_XI63/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI5/MM0 N_XI63/XI5/NET34_XI63/XI5/MM0_d N_WL<122>_XI63/XI5/MM0_g
+ N_BL<10>_XI63/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI5/MM1 N_XI63/XI5/NET33_XI63/XI5/MM1_d N_XI63/XI5/NET34_XI63/XI5/MM1_g
+ N_VSS_XI63/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI5/MM9 N_XI63/XI5/NET36_XI63/XI5/MM9_d N_WL<123>_XI63/XI5/MM9_g
+ N_BL<10>_XI63/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI5/MM6 N_XI63/XI5/NET35_XI63/XI5/MM6_d N_XI63/XI5/NET36_XI63/XI5/MM6_g
+ N_VSS_XI63/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI5/MM7 N_XI63/XI5/NET36_XI63/XI5/MM7_d N_XI63/XI5/NET35_XI63/XI5/MM7_g
+ N_VSS_XI63/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI5/MM8 N_XI63/XI5/NET35_XI63/XI5/MM8_d N_WL<123>_XI63/XI5/MM8_g
+ N_BLN<10>_XI63/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI5/MM5 N_XI63/XI5/NET34_XI63/XI5/MM5_d N_XI63/XI5/NET33_XI63/XI5/MM5_g
+ N_VDD_XI63/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI5/MM4 N_XI63/XI5/NET33_XI63/XI5/MM4_d N_XI63/XI5/NET34_XI63/XI5/MM4_g
+ N_VDD_XI63/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI5/MM10 N_XI63/XI5/NET35_XI63/XI5/MM10_d N_XI63/XI5/NET36_XI63/XI5/MM10_g
+ N_VDD_XI63/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI5/MM11 N_XI63/XI5/NET36_XI63/XI5/MM11_d N_XI63/XI5/NET35_XI63/XI5/MM11_g
+ N_VDD_XI63/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI6/MM2 N_XI63/XI6/NET34_XI63/XI6/MM2_d N_XI63/XI6/NET33_XI63/XI6/MM2_g
+ N_VSS_XI63/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM3 N_XI63/XI6/NET33_XI63/XI6/MM3_d N_WL<122>_XI63/XI6/MM3_g
+ N_BLN<9>_XI63/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM0 N_XI63/XI6/NET34_XI63/XI6/MM0_d N_WL<122>_XI63/XI6/MM0_g
+ N_BL<9>_XI63/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM1 N_XI63/XI6/NET33_XI63/XI6/MM1_d N_XI63/XI6/NET34_XI63/XI6/MM1_g
+ N_VSS_XI63/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM9 N_XI63/XI6/NET36_XI63/XI6/MM9_d N_WL<123>_XI63/XI6/MM9_g
+ N_BL<9>_XI63/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM6 N_XI63/XI6/NET35_XI63/XI6/MM6_d N_XI63/XI6/NET36_XI63/XI6/MM6_g
+ N_VSS_XI63/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM7 N_XI63/XI6/NET36_XI63/XI6/MM7_d N_XI63/XI6/NET35_XI63/XI6/MM7_g
+ N_VSS_XI63/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM8 N_XI63/XI6/NET35_XI63/XI6/MM8_d N_WL<123>_XI63/XI6/MM8_g
+ N_BLN<9>_XI63/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI6/MM5 N_XI63/XI6/NET34_XI63/XI6/MM5_d N_XI63/XI6/NET33_XI63/XI6/MM5_g
+ N_VDD_XI63/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI6/MM4 N_XI63/XI6/NET33_XI63/XI6/MM4_d N_XI63/XI6/NET34_XI63/XI6/MM4_g
+ N_VDD_XI63/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI6/MM10 N_XI63/XI6/NET35_XI63/XI6/MM10_d N_XI63/XI6/NET36_XI63/XI6/MM10_g
+ N_VDD_XI63/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI6/MM11 N_XI63/XI6/NET36_XI63/XI6/MM11_d N_XI63/XI6/NET35_XI63/XI6/MM11_g
+ N_VDD_XI63/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI7/MM2 N_XI63/XI7/NET34_XI63/XI7/MM2_d N_XI63/XI7/NET33_XI63/XI7/MM2_g
+ N_VSS_XI63/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM3 N_XI63/XI7/NET33_XI63/XI7/MM3_d N_WL<122>_XI63/XI7/MM3_g
+ N_BLN<8>_XI63/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM0 N_XI63/XI7/NET34_XI63/XI7/MM0_d N_WL<122>_XI63/XI7/MM0_g
+ N_BL<8>_XI63/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM1 N_XI63/XI7/NET33_XI63/XI7/MM1_d N_XI63/XI7/NET34_XI63/XI7/MM1_g
+ N_VSS_XI63/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM9 N_XI63/XI7/NET36_XI63/XI7/MM9_d N_WL<123>_XI63/XI7/MM9_g
+ N_BL<8>_XI63/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM6 N_XI63/XI7/NET35_XI63/XI7/MM6_d N_XI63/XI7/NET36_XI63/XI7/MM6_g
+ N_VSS_XI63/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM7 N_XI63/XI7/NET36_XI63/XI7/MM7_d N_XI63/XI7/NET35_XI63/XI7/MM7_g
+ N_VSS_XI63/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM8 N_XI63/XI7/NET35_XI63/XI7/MM8_d N_WL<123>_XI63/XI7/MM8_g
+ N_BLN<8>_XI63/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI7/MM5 N_XI63/XI7/NET34_XI63/XI7/MM5_d N_XI63/XI7/NET33_XI63/XI7/MM5_g
+ N_VDD_XI63/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI7/MM4 N_XI63/XI7/NET33_XI63/XI7/MM4_d N_XI63/XI7/NET34_XI63/XI7/MM4_g
+ N_VDD_XI63/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI7/MM10 N_XI63/XI7/NET35_XI63/XI7/MM10_d N_XI63/XI7/NET36_XI63/XI7/MM10_g
+ N_VDD_XI63/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI7/MM11 N_XI63/XI7/NET36_XI63/XI7/MM11_d N_XI63/XI7/NET35_XI63/XI7/MM11_g
+ N_VDD_XI63/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI8/MM2 N_XI63/XI8/NET34_XI63/XI8/MM2_d N_XI63/XI8/NET33_XI63/XI8/MM2_g
+ N_VSS_XI63/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM3 N_XI63/XI8/NET33_XI63/XI8/MM3_d N_WL<122>_XI63/XI8/MM3_g
+ N_BLN<7>_XI63/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM0 N_XI63/XI8/NET34_XI63/XI8/MM0_d N_WL<122>_XI63/XI8/MM0_g
+ N_BL<7>_XI63/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM1 N_XI63/XI8/NET33_XI63/XI8/MM1_d N_XI63/XI8/NET34_XI63/XI8/MM1_g
+ N_VSS_XI63/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM9 N_XI63/XI8/NET36_XI63/XI8/MM9_d N_WL<123>_XI63/XI8/MM9_g
+ N_BL<7>_XI63/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM6 N_XI63/XI8/NET35_XI63/XI8/MM6_d N_XI63/XI8/NET36_XI63/XI8/MM6_g
+ N_VSS_XI63/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM7 N_XI63/XI8/NET36_XI63/XI8/MM7_d N_XI63/XI8/NET35_XI63/XI8/MM7_g
+ N_VSS_XI63/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM8 N_XI63/XI8/NET35_XI63/XI8/MM8_d N_WL<123>_XI63/XI8/MM8_g
+ N_BLN<7>_XI63/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI8/MM5 N_XI63/XI8/NET34_XI63/XI8/MM5_d N_XI63/XI8/NET33_XI63/XI8/MM5_g
+ N_VDD_XI63/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI8/MM4 N_XI63/XI8/NET33_XI63/XI8/MM4_d N_XI63/XI8/NET34_XI63/XI8/MM4_g
+ N_VDD_XI63/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI8/MM10 N_XI63/XI8/NET35_XI63/XI8/MM10_d N_XI63/XI8/NET36_XI63/XI8/MM10_g
+ N_VDD_XI63/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI8/MM11 N_XI63/XI8/NET36_XI63/XI8/MM11_d N_XI63/XI8/NET35_XI63/XI8/MM11_g
+ N_VDD_XI63/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI9/MM2 N_XI63/XI9/NET34_XI63/XI9/MM2_d N_XI63/XI9/NET33_XI63/XI9/MM2_g
+ N_VSS_XI63/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM3 N_XI63/XI9/NET33_XI63/XI9/MM3_d N_WL<122>_XI63/XI9/MM3_g
+ N_BLN<6>_XI63/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM0 N_XI63/XI9/NET34_XI63/XI9/MM0_d N_WL<122>_XI63/XI9/MM0_g
+ N_BL<6>_XI63/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM1 N_XI63/XI9/NET33_XI63/XI9/MM1_d N_XI63/XI9/NET34_XI63/XI9/MM1_g
+ N_VSS_XI63/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM9 N_XI63/XI9/NET36_XI63/XI9/MM9_d N_WL<123>_XI63/XI9/MM9_g
+ N_BL<6>_XI63/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM6 N_XI63/XI9/NET35_XI63/XI9/MM6_d N_XI63/XI9/NET36_XI63/XI9/MM6_g
+ N_VSS_XI63/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM7 N_XI63/XI9/NET36_XI63/XI9/MM7_d N_XI63/XI9/NET35_XI63/XI9/MM7_g
+ N_VSS_XI63/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM8 N_XI63/XI9/NET35_XI63/XI9/MM8_d N_WL<123>_XI63/XI9/MM8_g
+ N_BLN<6>_XI63/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI9/MM5 N_XI63/XI9/NET34_XI63/XI9/MM5_d N_XI63/XI9/NET33_XI63/XI9/MM5_g
+ N_VDD_XI63/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI9/MM4 N_XI63/XI9/NET33_XI63/XI9/MM4_d N_XI63/XI9/NET34_XI63/XI9/MM4_g
+ N_VDD_XI63/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI9/MM10 N_XI63/XI9/NET35_XI63/XI9/MM10_d N_XI63/XI9/NET36_XI63/XI9/MM10_g
+ N_VDD_XI63/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI9/MM11 N_XI63/XI9/NET36_XI63/XI9/MM11_d N_XI63/XI9/NET35_XI63/XI9/MM11_g
+ N_VDD_XI63/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI10/MM2 N_XI63/XI10/NET34_XI63/XI10/MM2_d
+ N_XI63/XI10/NET33_XI63/XI10/MM2_g N_VSS_XI63/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI10/MM3 N_XI63/XI10/NET33_XI63/XI10/MM3_d N_WL<122>_XI63/XI10/MM3_g
+ N_BLN<5>_XI63/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI10/MM0 N_XI63/XI10/NET34_XI63/XI10/MM0_d N_WL<122>_XI63/XI10/MM0_g
+ N_BL<5>_XI63/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI10/MM1 N_XI63/XI10/NET33_XI63/XI10/MM1_d
+ N_XI63/XI10/NET34_XI63/XI10/MM1_g N_VSS_XI63/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI10/MM9 N_XI63/XI10/NET36_XI63/XI10/MM9_d N_WL<123>_XI63/XI10/MM9_g
+ N_BL<5>_XI63/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI10/MM6 N_XI63/XI10/NET35_XI63/XI10/MM6_d
+ N_XI63/XI10/NET36_XI63/XI10/MM6_g N_VSS_XI63/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI10/MM7 N_XI63/XI10/NET36_XI63/XI10/MM7_d
+ N_XI63/XI10/NET35_XI63/XI10/MM7_g N_VSS_XI63/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI10/MM8 N_XI63/XI10/NET35_XI63/XI10/MM8_d N_WL<123>_XI63/XI10/MM8_g
+ N_BLN<5>_XI63/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI10/MM5 N_XI63/XI10/NET34_XI63/XI10/MM5_d
+ N_XI63/XI10/NET33_XI63/XI10/MM5_g N_VDD_XI63/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI10/MM4 N_XI63/XI10/NET33_XI63/XI10/MM4_d
+ N_XI63/XI10/NET34_XI63/XI10/MM4_g N_VDD_XI63/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI10/MM10 N_XI63/XI10/NET35_XI63/XI10/MM10_d
+ N_XI63/XI10/NET36_XI63/XI10/MM10_g N_VDD_XI63/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI10/MM11 N_XI63/XI10/NET36_XI63/XI10/MM11_d
+ N_XI63/XI10/NET35_XI63/XI10/MM11_g N_VDD_XI63/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI11/MM2 N_XI63/XI11/NET34_XI63/XI11/MM2_d
+ N_XI63/XI11/NET33_XI63/XI11/MM2_g N_VSS_XI63/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI11/MM3 N_XI63/XI11/NET33_XI63/XI11/MM3_d N_WL<122>_XI63/XI11/MM3_g
+ N_BLN<4>_XI63/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI11/MM0 N_XI63/XI11/NET34_XI63/XI11/MM0_d N_WL<122>_XI63/XI11/MM0_g
+ N_BL<4>_XI63/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI11/MM1 N_XI63/XI11/NET33_XI63/XI11/MM1_d
+ N_XI63/XI11/NET34_XI63/XI11/MM1_g N_VSS_XI63/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI11/MM9 N_XI63/XI11/NET36_XI63/XI11/MM9_d N_WL<123>_XI63/XI11/MM9_g
+ N_BL<4>_XI63/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI11/MM6 N_XI63/XI11/NET35_XI63/XI11/MM6_d
+ N_XI63/XI11/NET36_XI63/XI11/MM6_g N_VSS_XI63/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI11/MM7 N_XI63/XI11/NET36_XI63/XI11/MM7_d
+ N_XI63/XI11/NET35_XI63/XI11/MM7_g N_VSS_XI63/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI11/MM8 N_XI63/XI11/NET35_XI63/XI11/MM8_d N_WL<123>_XI63/XI11/MM8_g
+ N_BLN<4>_XI63/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI11/MM5 N_XI63/XI11/NET34_XI63/XI11/MM5_d
+ N_XI63/XI11/NET33_XI63/XI11/MM5_g N_VDD_XI63/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI11/MM4 N_XI63/XI11/NET33_XI63/XI11/MM4_d
+ N_XI63/XI11/NET34_XI63/XI11/MM4_g N_VDD_XI63/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI11/MM10 N_XI63/XI11/NET35_XI63/XI11/MM10_d
+ N_XI63/XI11/NET36_XI63/XI11/MM10_g N_VDD_XI63/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI11/MM11 N_XI63/XI11/NET36_XI63/XI11/MM11_d
+ N_XI63/XI11/NET35_XI63/XI11/MM11_g N_VDD_XI63/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI12/MM2 N_XI63/XI12/NET34_XI63/XI12/MM2_d
+ N_XI63/XI12/NET33_XI63/XI12/MM2_g N_VSS_XI63/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI12/MM3 N_XI63/XI12/NET33_XI63/XI12/MM3_d N_WL<122>_XI63/XI12/MM3_g
+ N_BLN<3>_XI63/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI12/MM0 N_XI63/XI12/NET34_XI63/XI12/MM0_d N_WL<122>_XI63/XI12/MM0_g
+ N_BL<3>_XI63/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI12/MM1 N_XI63/XI12/NET33_XI63/XI12/MM1_d
+ N_XI63/XI12/NET34_XI63/XI12/MM1_g N_VSS_XI63/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI12/MM9 N_XI63/XI12/NET36_XI63/XI12/MM9_d N_WL<123>_XI63/XI12/MM9_g
+ N_BL<3>_XI63/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI12/MM6 N_XI63/XI12/NET35_XI63/XI12/MM6_d
+ N_XI63/XI12/NET36_XI63/XI12/MM6_g N_VSS_XI63/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI12/MM7 N_XI63/XI12/NET36_XI63/XI12/MM7_d
+ N_XI63/XI12/NET35_XI63/XI12/MM7_g N_VSS_XI63/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI12/MM8 N_XI63/XI12/NET35_XI63/XI12/MM8_d N_WL<123>_XI63/XI12/MM8_g
+ N_BLN<3>_XI63/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI12/MM5 N_XI63/XI12/NET34_XI63/XI12/MM5_d
+ N_XI63/XI12/NET33_XI63/XI12/MM5_g N_VDD_XI63/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI12/MM4 N_XI63/XI12/NET33_XI63/XI12/MM4_d
+ N_XI63/XI12/NET34_XI63/XI12/MM4_g N_VDD_XI63/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI12/MM10 N_XI63/XI12/NET35_XI63/XI12/MM10_d
+ N_XI63/XI12/NET36_XI63/XI12/MM10_g N_VDD_XI63/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI12/MM11 N_XI63/XI12/NET36_XI63/XI12/MM11_d
+ N_XI63/XI12/NET35_XI63/XI12/MM11_g N_VDD_XI63/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI13/MM2 N_XI63/XI13/NET34_XI63/XI13/MM2_d
+ N_XI63/XI13/NET33_XI63/XI13/MM2_g N_VSS_XI63/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI13/MM3 N_XI63/XI13/NET33_XI63/XI13/MM3_d N_WL<122>_XI63/XI13/MM3_g
+ N_BLN<2>_XI63/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI13/MM0 N_XI63/XI13/NET34_XI63/XI13/MM0_d N_WL<122>_XI63/XI13/MM0_g
+ N_BL<2>_XI63/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI13/MM1 N_XI63/XI13/NET33_XI63/XI13/MM1_d
+ N_XI63/XI13/NET34_XI63/XI13/MM1_g N_VSS_XI63/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI13/MM9 N_XI63/XI13/NET36_XI63/XI13/MM9_d N_WL<123>_XI63/XI13/MM9_g
+ N_BL<2>_XI63/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI13/MM6 N_XI63/XI13/NET35_XI63/XI13/MM6_d
+ N_XI63/XI13/NET36_XI63/XI13/MM6_g N_VSS_XI63/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI13/MM7 N_XI63/XI13/NET36_XI63/XI13/MM7_d
+ N_XI63/XI13/NET35_XI63/XI13/MM7_g N_VSS_XI63/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI13/MM8 N_XI63/XI13/NET35_XI63/XI13/MM8_d N_WL<123>_XI63/XI13/MM8_g
+ N_BLN<2>_XI63/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI13/MM5 N_XI63/XI13/NET34_XI63/XI13/MM5_d
+ N_XI63/XI13/NET33_XI63/XI13/MM5_g N_VDD_XI63/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI13/MM4 N_XI63/XI13/NET33_XI63/XI13/MM4_d
+ N_XI63/XI13/NET34_XI63/XI13/MM4_g N_VDD_XI63/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI13/MM10 N_XI63/XI13/NET35_XI63/XI13/MM10_d
+ N_XI63/XI13/NET36_XI63/XI13/MM10_g N_VDD_XI63/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI13/MM11 N_XI63/XI13/NET36_XI63/XI13/MM11_d
+ N_XI63/XI13/NET35_XI63/XI13/MM11_g N_VDD_XI63/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI14/MM2 N_XI63/XI14/NET34_XI63/XI14/MM2_d
+ N_XI63/XI14/NET33_XI63/XI14/MM2_g N_VSS_XI63/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI14/MM3 N_XI63/XI14/NET33_XI63/XI14/MM3_d N_WL<122>_XI63/XI14/MM3_g
+ N_BLN<1>_XI63/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI14/MM0 N_XI63/XI14/NET34_XI63/XI14/MM0_d N_WL<122>_XI63/XI14/MM0_g
+ N_BL<1>_XI63/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI14/MM1 N_XI63/XI14/NET33_XI63/XI14/MM1_d
+ N_XI63/XI14/NET34_XI63/XI14/MM1_g N_VSS_XI63/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI14/MM9 N_XI63/XI14/NET36_XI63/XI14/MM9_d N_WL<123>_XI63/XI14/MM9_g
+ N_BL<1>_XI63/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI14/MM6 N_XI63/XI14/NET35_XI63/XI14/MM6_d
+ N_XI63/XI14/NET36_XI63/XI14/MM6_g N_VSS_XI63/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI14/MM7 N_XI63/XI14/NET36_XI63/XI14/MM7_d
+ N_XI63/XI14/NET35_XI63/XI14/MM7_g N_VSS_XI63/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI14/MM8 N_XI63/XI14/NET35_XI63/XI14/MM8_d N_WL<123>_XI63/XI14/MM8_g
+ N_BLN<1>_XI63/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI14/MM5 N_XI63/XI14/NET34_XI63/XI14/MM5_d
+ N_XI63/XI14/NET33_XI63/XI14/MM5_g N_VDD_XI63/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI14/MM4 N_XI63/XI14/NET33_XI63/XI14/MM4_d
+ N_XI63/XI14/NET34_XI63/XI14/MM4_g N_VDD_XI63/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI14/MM10 N_XI63/XI14/NET35_XI63/XI14/MM10_d
+ N_XI63/XI14/NET36_XI63/XI14/MM10_g N_VDD_XI63/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI14/MM11 N_XI63/XI14/NET36_XI63/XI14/MM11_d
+ N_XI63/XI14/NET35_XI63/XI14/MM11_g N_VDD_XI63/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI15/MM2 N_XI63/XI15/NET34_XI63/XI15/MM2_d
+ N_XI63/XI15/NET33_XI63/XI15/MM2_g N_VSS_XI63/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI15/MM3 N_XI63/XI15/NET33_XI63/XI15/MM3_d N_WL<122>_XI63/XI15/MM3_g
+ N_BLN<0>_XI63/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI15/MM0 N_XI63/XI15/NET34_XI63/XI15/MM0_d N_WL<122>_XI63/XI15/MM0_g
+ N_BL<0>_XI63/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI15/MM1 N_XI63/XI15/NET33_XI63/XI15/MM1_d
+ N_XI63/XI15/NET34_XI63/XI15/MM1_g N_VSS_XI63/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI15/MM9 N_XI63/XI15/NET36_XI63/XI15/MM9_d N_WL<123>_XI63/XI15/MM9_g
+ N_BL<0>_XI63/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI15/MM6 N_XI63/XI15/NET35_XI63/XI15/MM6_d
+ N_XI63/XI15/NET36_XI63/XI15/MM6_g N_VSS_XI63/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI15/MM7 N_XI63/XI15/NET36_XI63/XI15/MM7_d
+ N_XI63/XI15/NET35_XI63/XI15/MM7_g N_VSS_XI63/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI63/XI15/MM8 N_XI63/XI15/NET35_XI63/XI15/MM8_d N_WL<123>_XI63/XI15/MM8_g
+ N_BLN<0>_XI63/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI63/XI15/MM5 N_XI63/XI15/NET34_XI63/XI15/MM5_d
+ N_XI63/XI15/NET33_XI63/XI15/MM5_g N_VDD_XI63/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI15/MM4 N_XI63/XI15/NET33_XI63/XI15/MM4_d
+ N_XI63/XI15/NET34_XI63/XI15/MM4_g N_VDD_XI63/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI15/MM10 N_XI63/XI15/NET35_XI63/XI15/MM10_d
+ N_XI63/XI15/NET36_XI63/XI15/MM10_g N_VDD_XI63/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI63/XI15/MM11 N_XI63/XI15/NET36_XI63/XI15/MM11_d
+ N_XI63/XI15/NET35_XI63/XI15/MM11_g N_VDD_XI63/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI0/MM2 N_XI64/XI0/NET34_XI64/XI0/MM2_d N_XI64/XI0/NET33_XI64/XI0/MM2_g
+ N_VSS_XI64/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI0/MM3 N_XI64/XI0/NET33_XI64/XI0/MM3_d N_WL<124>_XI64/XI0/MM3_g
+ N_BLN<15>_XI64/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI0/MM0 N_XI64/XI0/NET34_XI64/XI0/MM0_d N_WL<124>_XI64/XI0/MM0_g
+ N_BL<15>_XI64/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI0/MM1 N_XI64/XI0/NET33_XI64/XI0/MM1_d N_XI64/XI0/NET34_XI64/XI0/MM1_g
+ N_VSS_XI64/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI0/MM9 N_XI64/XI0/NET36_XI64/XI0/MM9_d N_WL<125>_XI64/XI0/MM9_g
+ N_BL<15>_XI64/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI0/MM6 N_XI64/XI0/NET35_XI64/XI0/MM6_d N_XI64/XI0/NET36_XI64/XI0/MM6_g
+ N_VSS_XI64/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI0/MM7 N_XI64/XI0/NET36_XI64/XI0/MM7_d N_XI64/XI0/NET35_XI64/XI0/MM7_g
+ N_VSS_XI64/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI0/MM8 N_XI64/XI0/NET35_XI64/XI0/MM8_d N_WL<125>_XI64/XI0/MM8_g
+ N_BLN<15>_XI64/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI0/MM5 N_XI64/XI0/NET34_XI64/XI0/MM5_d N_XI64/XI0/NET33_XI64/XI0/MM5_g
+ N_VDD_XI64/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI0/MM4 N_XI64/XI0/NET33_XI64/XI0/MM4_d N_XI64/XI0/NET34_XI64/XI0/MM4_g
+ N_VDD_XI64/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI0/MM10 N_XI64/XI0/NET35_XI64/XI0/MM10_d N_XI64/XI0/NET36_XI64/XI0/MM10_g
+ N_VDD_XI64/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI0/MM11 N_XI64/XI0/NET36_XI64/XI0/MM11_d N_XI64/XI0/NET35_XI64/XI0/MM11_g
+ N_VDD_XI64/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI1/MM2 N_XI64/XI1/NET34_XI64/XI1/MM2_d N_XI64/XI1/NET33_XI64/XI1/MM2_g
+ N_VSS_XI64/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI1/MM3 N_XI64/XI1/NET33_XI64/XI1/MM3_d N_WL<124>_XI64/XI1/MM3_g
+ N_BLN<14>_XI64/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI1/MM0 N_XI64/XI1/NET34_XI64/XI1/MM0_d N_WL<124>_XI64/XI1/MM0_g
+ N_BL<14>_XI64/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI1/MM1 N_XI64/XI1/NET33_XI64/XI1/MM1_d N_XI64/XI1/NET34_XI64/XI1/MM1_g
+ N_VSS_XI64/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI1/MM9 N_XI64/XI1/NET36_XI64/XI1/MM9_d N_WL<125>_XI64/XI1/MM9_g
+ N_BL<14>_XI64/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI1/MM6 N_XI64/XI1/NET35_XI64/XI1/MM6_d N_XI64/XI1/NET36_XI64/XI1/MM6_g
+ N_VSS_XI64/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI1/MM7 N_XI64/XI1/NET36_XI64/XI1/MM7_d N_XI64/XI1/NET35_XI64/XI1/MM7_g
+ N_VSS_XI64/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI1/MM8 N_XI64/XI1/NET35_XI64/XI1/MM8_d N_WL<125>_XI64/XI1/MM8_g
+ N_BLN<14>_XI64/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI1/MM5 N_XI64/XI1/NET34_XI64/XI1/MM5_d N_XI64/XI1/NET33_XI64/XI1/MM5_g
+ N_VDD_XI64/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI1/MM4 N_XI64/XI1/NET33_XI64/XI1/MM4_d N_XI64/XI1/NET34_XI64/XI1/MM4_g
+ N_VDD_XI64/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI1/MM10 N_XI64/XI1/NET35_XI64/XI1/MM10_d N_XI64/XI1/NET36_XI64/XI1/MM10_g
+ N_VDD_XI64/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI1/MM11 N_XI64/XI1/NET36_XI64/XI1/MM11_d N_XI64/XI1/NET35_XI64/XI1/MM11_g
+ N_VDD_XI64/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI2/MM2 N_XI64/XI2/NET34_XI64/XI2/MM2_d N_XI64/XI2/NET33_XI64/XI2/MM2_g
+ N_VSS_XI64/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI2/MM3 N_XI64/XI2/NET33_XI64/XI2/MM3_d N_WL<124>_XI64/XI2/MM3_g
+ N_BLN<13>_XI64/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI2/MM0 N_XI64/XI2/NET34_XI64/XI2/MM0_d N_WL<124>_XI64/XI2/MM0_g
+ N_BL<13>_XI64/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI2/MM1 N_XI64/XI2/NET33_XI64/XI2/MM1_d N_XI64/XI2/NET34_XI64/XI2/MM1_g
+ N_VSS_XI64/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI2/MM9 N_XI64/XI2/NET36_XI64/XI2/MM9_d N_WL<125>_XI64/XI2/MM9_g
+ N_BL<13>_XI64/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI2/MM6 N_XI64/XI2/NET35_XI64/XI2/MM6_d N_XI64/XI2/NET36_XI64/XI2/MM6_g
+ N_VSS_XI64/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI2/MM7 N_XI64/XI2/NET36_XI64/XI2/MM7_d N_XI64/XI2/NET35_XI64/XI2/MM7_g
+ N_VSS_XI64/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI2/MM8 N_XI64/XI2/NET35_XI64/XI2/MM8_d N_WL<125>_XI64/XI2/MM8_g
+ N_BLN<13>_XI64/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI2/MM5 N_XI64/XI2/NET34_XI64/XI2/MM5_d N_XI64/XI2/NET33_XI64/XI2/MM5_g
+ N_VDD_XI64/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI2/MM4 N_XI64/XI2/NET33_XI64/XI2/MM4_d N_XI64/XI2/NET34_XI64/XI2/MM4_g
+ N_VDD_XI64/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI2/MM10 N_XI64/XI2/NET35_XI64/XI2/MM10_d N_XI64/XI2/NET36_XI64/XI2/MM10_g
+ N_VDD_XI64/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI2/MM11 N_XI64/XI2/NET36_XI64/XI2/MM11_d N_XI64/XI2/NET35_XI64/XI2/MM11_g
+ N_VDD_XI64/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI3/MM2 N_XI64/XI3/NET34_XI64/XI3/MM2_d N_XI64/XI3/NET33_XI64/XI3/MM2_g
+ N_VSS_XI64/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI3/MM3 N_XI64/XI3/NET33_XI64/XI3/MM3_d N_WL<124>_XI64/XI3/MM3_g
+ N_BLN<12>_XI64/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI3/MM0 N_XI64/XI3/NET34_XI64/XI3/MM0_d N_WL<124>_XI64/XI3/MM0_g
+ N_BL<12>_XI64/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI3/MM1 N_XI64/XI3/NET33_XI64/XI3/MM1_d N_XI64/XI3/NET34_XI64/XI3/MM1_g
+ N_VSS_XI64/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI3/MM9 N_XI64/XI3/NET36_XI64/XI3/MM9_d N_WL<125>_XI64/XI3/MM9_g
+ N_BL<12>_XI64/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI3/MM6 N_XI64/XI3/NET35_XI64/XI3/MM6_d N_XI64/XI3/NET36_XI64/XI3/MM6_g
+ N_VSS_XI64/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI3/MM7 N_XI64/XI3/NET36_XI64/XI3/MM7_d N_XI64/XI3/NET35_XI64/XI3/MM7_g
+ N_VSS_XI64/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI3/MM8 N_XI64/XI3/NET35_XI64/XI3/MM8_d N_WL<125>_XI64/XI3/MM8_g
+ N_BLN<12>_XI64/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI3/MM5 N_XI64/XI3/NET34_XI64/XI3/MM5_d N_XI64/XI3/NET33_XI64/XI3/MM5_g
+ N_VDD_XI64/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI3/MM4 N_XI64/XI3/NET33_XI64/XI3/MM4_d N_XI64/XI3/NET34_XI64/XI3/MM4_g
+ N_VDD_XI64/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI3/MM10 N_XI64/XI3/NET35_XI64/XI3/MM10_d N_XI64/XI3/NET36_XI64/XI3/MM10_g
+ N_VDD_XI64/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI3/MM11 N_XI64/XI3/NET36_XI64/XI3/MM11_d N_XI64/XI3/NET35_XI64/XI3/MM11_g
+ N_VDD_XI64/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI4/MM2 N_XI64/XI4/NET34_XI64/XI4/MM2_d N_XI64/XI4/NET33_XI64/XI4/MM2_g
+ N_VSS_XI64/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI4/MM3 N_XI64/XI4/NET33_XI64/XI4/MM3_d N_WL<124>_XI64/XI4/MM3_g
+ N_BLN<11>_XI64/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI4/MM0 N_XI64/XI4/NET34_XI64/XI4/MM0_d N_WL<124>_XI64/XI4/MM0_g
+ N_BL<11>_XI64/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI4/MM1 N_XI64/XI4/NET33_XI64/XI4/MM1_d N_XI64/XI4/NET34_XI64/XI4/MM1_g
+ N_VSS_XI64/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI4/MM9 N_XI64/XI4/NET36_XI64/XI4/MM9_d N_WL<125>_XI64/XI4/MM9_g
+ N_BL<11>_XI64/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI4/MM6 N_XI64/XI4/NET35_XI64/XI4/MM6_d N_XI64/XI4/NET36_XI64/XI4/MM6_g
+ N_VSS_XI64/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI4/MM7 N_XI64/XI4/NET36_XI64/XI4/MM7_d N_XI64/XI4/NET35_XI64/XI4/MM7_g
+ N_VSS_XI64/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI4/MM8 N_XI64/XI4/NET35_XI64/XI4/MM8_d N_WL<125>_XI64/XI4/MM8_g
+ N_BLN<11>_XI64/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI4/MM5 N_XI64/XI4/NET34_XI64/XI4/MM5_d N_XI64/XI4/NET33_XI64/XI4/MM5_g
+ N_VDD_XI64/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI4/MM4 N_XI64/XI4/NET33_XI64/XI4/MM4_d N_XI64/XI4/NET34_XI64/XI4/MM4_g
+ N_VDD_XI64/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI4/MM10 N_XI64/XI4/NET35_XI64/XI4/MM10_d N_XI64/XI4/NET36_XI64/XI4/MM10_g
+ N_VDD_XI64/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI4/MM11 N_XI64/XI4/NET36_XI64/XI4/MM11_d N_XI64/XI4/NET35_XI64/XI4/MM11_g
+ N_VDD_XI64/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI5/MM2 N_XI64/XI5/NET34_XI64/XI5/MM2_d N_XI64/XI5/NET33_XI64/XI5/MM2_g
+ N_VSS_XI64/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI5/MM3 N_XI64/XI5/NET33_XI64/XI5/MM3_d N_WL<124>_XI64/XI5/MM3_g
+ N_BLN<10>_XI64/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI5/MM0 N_XI64/XI5/NET34_XI64/XI5/MM0_d N_WL<124>_XI64/XI5/MM0_g
+ N_BL<10>_XI64/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI5/MM1 N_XI64/XI5/NET33_XI64/XI5/MM1_d N_XI64/XI5/NET34_XI64/XI5/MM1_g
+ N_VSS_XI64/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI5/MM9 N_XI64/XI5/NET36_XI64/XI5/MM9_d N_WL<125>_XI64/XI5/MM9_g
+ N_BL<10>_XI64/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI5/MM6 N_XI64/XI5/NET35_XI64/XI5/MM6_d N_XI64/XI5/NET36_XI64/XI5/MM6_g
+ N_VSS_XI64/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI5/MM7 N_XI64/XI5/NET36_XI64/XI5/MM7_d N_XI64/XI5/NET35_XI64/XI5/MM7_g
+ N_VSS_XI64/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI5/MM8 N_XI64/XI5/NET35_XI64/XI5/MM8_d N_WL<125>_XI64/XI5/MM8_g
+ N_BLN<10>_XI64/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI5/MM5 N_XI64/XI5/NET34_XI64/XI5/MM5_d N_XI64/XI5/NET33_XI64/XI5/MM5_g
+ N_VDD_XI64/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI5/MM4 N_XI64/XI5/NET33_XI64/XI5/MM4_d N_XI64/XI5/NET34_XI64/XI5/MM4_g
+ N_VDD_XI64/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI5/MM10 N_XI64/XI5/NET35_XI64/XI5/MM10_d N_XI64/XI5/NET36_XI64/XI5/MM10_g
+ N_VDD_XI64/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI5/MM11 N_XI64/XI5/NET36_XI64/XI5/MM11_d N_XI64/XI5/NET35_XI64/XI5/MM11_g
+ N_VDD_XI64/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI6/MM2 N_XI64/XI6/NET34_XI64/XI6/MM2_d N_XI64/XI6/NET33_XI64/XI6/MM2_g
+ N_VSS_XI64/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM3 N_XI64/XI6/NET33_XI64/XI6/MM3_d N_WL<124>_XI64/XI6/MM3_g
+ N_BLN<9>_XI64/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM0 N_XI64/XI6/NET34_XI64/XI6/MM0_d N_WL<124>_XI64/XI6/MM0_g
+ N_BL<9>_XI64/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM1 N_XI64/XI6/NET33_XI64/XI6/MM1_d N_XI64/XI6/NET34_XI64/XI6/MM1_g
+ N_VSS_XI64/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM9 N_XI64/XI6/NET36_XI64/XI6/MM9_d N_WL<125>_XI64/XI6/MM9_g
+ N_BL<9>_XI64/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM6 N_XI64/XI6/NET35_XI64/XI6/MM6_d N_XI64/XI6/NET36_XI64/XI6/MM6_g
+ N_VSS_XI64/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM7 N_XI64/XI6/NET36_XI64/XI6/MM7_d N_XI64/XI6/NET35_XI64/XI6/MM7_g
+ N_VSS_XI64/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM8 N_XI64/XI6/NET35_XI64/XI6/MM8_d N_WL<125>_XI64/XI6/MM8_g
+ N_BLN<9>_XI64/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI6/MM5 N_XI64/XI6/NET34_XI64/XI6/MM5_d N_XI64/XI6/NET33_XI64/XI6/MM5_g
+ N_VDD_XI64/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI6/MM4 N_XI64/XI6/NET33_XI64/XI6/MM4_d N_XI64/XI6/NET34_XI64/XI6/MM4_g
+ N_VDD_XI64/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI6/MM10 N_XI64/XI6/NET35_XI64/XI6/MM10_d N_XI64/XI6/NET36_XI64/XI6/MM10_g
+ N_VDD_XI64/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI6/MM11 N_XI64/XI6/NET36_XI64/XI6/MM11_d N_XI64/XI6/NET35_XI64/XI6/MM11_g
+ N_VDD_XI64/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI7/MM2 N_XI64/XI7/NET34_XI64/XI7/MM2_d N_XI64/XI7/NET33_XI64/XI7/MM2_g
+ N_VSS_XI64/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM3 N_XI64/XI7/NET33_XI64/XI7/MM3_d N_WL<124>_XI64/XI7/MM3_g
+ N_BLN<8>_XI64/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM0 N_XI64/XI7/NET34_XI64/XI7/MM0_d N_WL<124>_XI64/XI7/MM0_g
+ N_BL<8>_XI64/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM1 N_XI64/XI7/NET33_XI64/XI7/MM1_d N_XI64/XI7/NET34_XI64/XI7/MM1_g
+ N_VSS_XI64/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM9 N_XI64/XI7/NET36_XI64/XI7/MM9_d N_WL<125>_XI64/XI7/MM9_g
+ N_BL<8>_XI64/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM6 N_XI64/XI7/NET35_XI64/XI7/MM6_d N_XI64/XI7/NET36_XI64/XI7/MM6_g
+ N_VSS_XI64/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM7 N_XI64/XI7/NET36_XI64/XI7/MM7_d N_XI64/XI7/NET35_XI64/XI7/MM7_g
+ N_VSS_XI64/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM8 N_XI64/XI7/NET35_XI64/XI7/MM8_d N_WL<125>_XI64/XI7/MM8_g
+ N_BLN<8>_XI64/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI7/MM5 N_XI64/XI7/NET34_XI64/XI7/MM5_d N_XI64/XI7/NET33_XI64/XI7/MM5_g
+ N_VDD_XI64/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI7/MM4 N_XI64/XI7/NET33_XI64/XI7/MM4_d N_XI64/XI7/NET34_XI64/XI7/MM4_g
+ N_VDD_XI64/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI7/MM10 N_XI64/XI7/NET35_XI64/XI7/MM10_d N_XI64/XI7/NET36_XI64/XI7/MM10_g
+ N_VDD_XI64/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI7/MM11 N_XI64/XI7/NET36_XI64/XI7/MM11_d N_XI64/XI7/NET35_XI64/XI7/MM11_g
+ N_VDD_XI64/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI8/MM2 N_XI64/XI8/NET34_XI64/XI8/MM2_d N_XI64/XI8/NET33_XI64/XI8/MM2_g
+ N_VSS_XI64/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM3 N_XI64/XI8/NET33_XI64/XI8/MM3_d N_WL<124>_XI64/XI8/MM3_g
+ N_BLN<7>_XI64/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM0 N_XI64/XI8/NET34_XI64/XI8/MM0_d N_WL<124>_XI64/XI8/MM0_g
+ N_BL<7>_XI64/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM1 N_XI64/XI8/NET33_XI64/XI8/MM1_d N_XI64/XI8/NET34_XI64/XI8/MM1_g
+ N_VSS_XI64/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM9 N_XI64/XI8/NET36_XI64/XI8/MM9_d N_WL<125>_XI64/XI8/MM9_g
+ N_BL<7>_XI64/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM6 N_XI64/XI8/NET35_XI64/XI8/MM6_d N_XI64/XI8/NET36_XI64/XI8/MM6_g
+ N_VSS_XI64/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM7 N_XI64/XI8/NET36_XI64/XI8/MM7_d N_XI64/XI8/NET35_XI64/XI8/MM7_g
+ N_VSS_XI64/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM8 N_XI64/XI8/NET35_XI64/XI8/MM8_d N_WL<125>_XI64/XI8/MM8_g
+ N_BLN<7>_XI64/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI8/MM5 N_XI64/XI8/NET34_XI64/XI8/MM5_d N_XI64/XI8/NET33_XI64/XI8/MM5_g
+ N_VDD_XI64/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI8/MM4 N_XI64/XI8/NET33_XI64/XI8/MM4_d N_XI64/XI8/NET34_XI64/XI8/MM4_g
+ N_VDD_XI64/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI8/MM10 N_XI64/XI8/NET35_XI64/XI8/MM10_d N_XI64/XI8/NET36_XI64/XI8/MM10_g
+ N_VDD_XI64/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI8/MM11 N_XI64/XI8/NET36_XI64/XI8/MM11_d N_XI64/XI8/NET35_XI64/XI8/MM11_g
+ N_VDD_XI64/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI9/MM2 N_XI64/XI9/NET34_XI64/XI9/MM2_d N_XI64/XI9/NET33_XI64/XI9/MM2_g
+ N_VSS_XI64/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM3 N_XI64/XI9/NET33_XI64/XI9/MM3_d N_WL<124>_XI64/XI9/MM3_g
+ N_BLN<6>_XI64/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM0 N_XI64/XI9/NET34_XI64/XI9/MM0_d N_WL<124>_XI64/XI9/MM0_g
+ N_BL<6>_XI64/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM1 N_XI64/XI9/NET33_XI64/XI9/MM1_d N_XI64/XI9/NET34_XI64/XI9/MM1_g
+ N_VSS_XI64/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM9 N_XI64/XI9/NET36_XI64/XI9/MM9_d N_WL<125>_XI64/XI9/MM9_g
+ N_BL<6>_XI64/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM6 N_XI64/XI9/NET35_XI64/XI9/MM6_d N_XI64/XI9/NET36_XI64/XI9/MM6_g
+ N_VSS_XI64/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM7 N_XI64/XI9/NET36_XI64/XI9/MM7_d N_XI64/XI9/NET35_XI64/XI9/MM7_g
+ N_VSS_XI64/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM8 N_XI64/XI9/NET35_XI64/XI9/MM8_d N_WL<125>_XI64/XI9/MM8_g
+ N_BLN<6>_XI64/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI9/MM5 N_XI64/XI9/NET34_XI64/XI9/MM5_d N_XI64/XI9/NET33_XI64/XI9/MM5_g
+ N_VDD_XI64/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI9/MM4 N_XI64/XI9/NET33_XI64/XI9/MM4_d N_XI64/XI9/NET34_XI64/XI9/MM4_g
+ N_VDD_XI64/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI9/MM10 N_XI64/XI9/NET35_XI64/XI9/MM10_d N_XI64/XI9/NET36_XI64/XI9/MM10_g
+ N_VDD_XI64/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI9/MM11 N_XI64/XI9/NET36_XI64/XI9/MM11_d N_XI64/XI9/NET35_XI64/XI9/MM11_g
+ N_VDD_XI64/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI10/MM2 N_XI64/XI10/NET34_XI64/XI10/MM2_d
+ N_XI64/XI10/NET33_XI64/XI10/MM2_g N_VSS_XI64/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI10/MM3 N_XI64/XI10/NET33_XI64/XI10/MM3_d N_WL<124>_XI64/XI10/MM3_g
+ N_BLN<5>_XI64/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI10/MM0 N_XI64/XI10/NET34_XI64/XI10/MM0_d N_WL<124>_XI64/XI10/MM0_g
+ N_BL<5>_XI64/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI10/MM1 N_XI64/XI10/NET33_XI64/XI10/MM1_d
+ N_XI64/XI10/NET34_XI64/XI10/MM1_g N_VSS_XI64/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI10/MM9 N_XI64/XI10/NET36_XI64/XI10/MM9_d N_WL<125>_XI64/XI10/MM9_g
+ N_BL<5>_XI64/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI10/MM6 N_XI64/XI10/NET35_XI64/XI10/MM6_d
+ N_XI64/XI10/NET36_XI64/XI10/MM6_g N_VSS_XI64/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI10/MM7 N_XI64/XI10/NET36_XI64/XI10/MM7_d
+ N_XI64/XI10/NET35_XI64/XI10/MM7_g N_VSS_XI64/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI10/MM8 N_XI64/XI10/NET35_XI64/XI10/MM8_d N_WL<125>_XI64/XI10/MM8_g
+ N_BLN<5>_XI64/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI10/MM5 N_XI64/XI10/NET34_XI64/XI10/MM5_d
+ N_XI64/XI10/NET33_XI64/XI10/MM5_g N_VDD_XI64/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI10/MM4 N_XI64/XI10/NET33_XI64/XI10/MM4_d
+ N_XI64/XI10/NET34_XI64/XI10/MM4_g N_VDD_XI64/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI10/MM10 N_XI64/XI10/NET35_XI64/XI10/MM10_d
+ N_XI64/XI10/NET36_XI64/XI10/MM10_g N_VDD_XI64/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI10/MM11 N_XI64/XI10/NET36_XI64/XI10/MM11_d
+ N_XI64/XI10/NET35_XI64/XI10/MM11_g N_VDD_XI64/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI11/MM2 N_XI64/XI11/NET34_XI64/XI11/MM2_d
+ N_XI64/XI11/NET33_XI64/XI11/MM2_g N_VSS_XI64/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI11/MM3 N_XI64/XI11/NET33_XI64/XI11/MM3_d N_WL<124>_XI64/XI11/MM3_g
+ N_BLN<4>_XI64/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI11/MM0 N_XI64/XI11/NET34_XI64/XI11/MM0_d N_WL<124>_XI64/XI11/MM0_g
+ N_BL<4>_XI64/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI11/MM1 N_XI64/XI11/NET33_XI64/XI11/MM1_d
+ N_XI64/XI11/NET34_XI64/XI11/MM1_g N_VSS_XI64/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI11/MM9 N_XI64/XI11/NET36_XI64/XI11/MM9_d N_WL<125>_XI64/XI11/MM9_g
+ N_BL<4>_XI64/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI11/MM6 N_XI64/XI11/NET35_XI64/XI11/MM6_d
+ N_XI64/XI11/NET36_XI64/XI11/MM6_g N_VSS_XI64/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI11/MM7 N_XI64/XI11/NET36_XI64/XI11/MM7_d
+ N_XI64/XI11/NET35_XI64/XI11/MM7_g N_VSS_XI64/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI11/MM8 N_XI64/XI11/NET35_XI64/XI11/MM8_d N_WL<125>_XI64/XI11/MM8_g
+ N_BLN<4>_XI64/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI11/MM5 N_XI64/XI11/NET34_XI64/XI11/MM5_d
+ N_XI64/XI11/NET33_XI64/XI11/MM5_g N_VDD_XI64/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI11/MM4 N_XI64/XI11/NET33_XI64/XI11/MM4_d
+ N_XI64/XI11/NET34_XI64/XI11/MM4_g N_VDD_XI64/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI11/MM10 N_XI64/XI11/NET35_XI64/XI11/MM10_d
+ N_XI64/XI11/NET36_XI64/XI11/MM10_g N_VDD_XI64/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI11/MM11 N_XI64/XI11/NET36_XI64/XI11/MM11_d
+ N_XI64/XI11/NET35_XI64/XI11/MM11_g N_VDD_XI64/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI12/MM2 N_XI64/XI12/NET34_XI64/XI12/MM2_d
+ N_XI64/XI12/NET33_XI64/XI12/MM2_g N_VSS_XI64/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI12/MM3 N_XI64/XI12/NET33_XI64/XI12/MM3_d N_WL<124>_XI64/XI12/MM3_g
+ N_BLN<3>_XI64/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI12/MM0 N_XI64/XI12/NET34_XI64/XI12/MM0_d N_WL<124>_XI64/XI12/MM0_g
+ N_BL<3>_XI64/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI12/MM1 N_XI64/XI12/NET33_XI64/XI12/MM1_d
+ N_XI64/XI12/NET34_XI64/XI12/MM1_g N_VSS_XI64/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI12/MM9 N_XI64/XI12/NET36_XI64/XI12/MM9_d N_WL<125>_XI64/XI12/MM9_g
+ N_BL<3>_XI64/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI12/MM6 N_XI64/XI12/NET35_XI64/XI12/MM6_d
+ N_XI64/XI12/NET36_XI64/XI12/MM6_g N_VSS_XI64/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI12/MM7 N_XI64/XI12/NET36_XI64/XI12/MM7_d
+ N_XI64/XI12/NET35_XI64/XI12/MM7_g N_VSS_XI64/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI12/MM8 N_XI64/XI12/NET35_XI64/XI12/MM8_d N_WL<125>_XI64/XI12/MM8_g
+ N_BLN<3>_XI64/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI12/MM5 N_XI64/XI12/NET34_XI64/XI12/MM5_d
+ N_XI64/XI12/NET33_XI64/XI12/MM5_g N_VDD_XI64/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI12/MM4 N_XI64/XI12/NET33_XI64/XI12/MM4_d
+ N_XI64/XI12/NET34_XI64/XI12/MM4_g N_VDD_XI64/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI12/MM10 N_XI64/XI12/NET35_XI64/XI12/MM10_d
+ N_XI64/XI12/NET36_XI64/XI12/MM10_g N_VDD_XI64/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI12/MM11 N_XI64/XI12/NET36_XI64/XI12/MM11_d
+ N_XI64/XI12/NET35_XI64/XI12/MM11_g N_VDD_XI64/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI13/MM2 N_XI64/XI13/NET34_XI64/XI13/MM2_d
+ N_XI64/XI13/NET33_XI64/XI13/MM2_g N_VSS_XI64/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI13/MM3 N_XI64/XI13/NET33_XI64/XI13/MM3_d N_WL<124>_XI64/XI13/MM3_g
+ N_BLN<2>_XI64/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI13/MM0 N_XI64/XI13/NET34_XI64/XI13/MM0_d N_WL<124>_XI64/XI13/MM0_g
+ N_BL<2>_XI64/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI13/MM1 N_XI64/XI13/NET33_XI64/XI13/MM1_d
+ N_XI64/XI13/NET34_XI64/XI13/MM1_g N_VSS_XI64/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI13/MM9 N_XI64/XI13/NET36_XI64/XI13/MM9_d N_WL<125>_XI64/XI13/MM9_g
+ N_BL<2>_XI64/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI13/MM6 N_XI64/XI13/NET35_XI64/XI13/MM6_d
+ N_XI64/XI13/NET36_XI64/XI13/MM6_g N_VSS_XI64/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI13/MM7 N_XI64/XI13/NET36_XI64/XI13/MM7_d
+ N_XI64/XI13/NET35_XI64/XI13/MM7_g N_VSS_XI64/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI13/MM8 N_XI64/XI13/NET35_XI64/XI13/MM8_d N_WL<125>_XI64/XI13/MM8_g
+ N_BLN<2>_XI64/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI13/MM5 N_XI64/XI13/NET34_XI64/XI13/MM5_d
+ N_XI64/XI13/NET33_XI64/XI13/MM5_g N_VDD_XI64/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI13/MM4 N_XI64/XI13/NET33_XI64/XI13/MM4_d
+ N_XI64/XI13/NET34_XI64/XI13/MM4_g N_VDD_XI64/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI13/MM10 N_XI64/XI13/NET35_XI64/XI13/MM10_d
+ N_XI64/XI13/NET36_XI64/XI13/MM10_g N_VDD_XI64/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI13/MM11 N_XI64/XI13/NET36_XI64/XI13/MM11_d
+ N_XI64/XI13/NET35_XI64/XI13/MM11_g N_VDD_XI64/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI14/MM2 N_XI64/XI14/NET34_XI64/XI14/MM2_d
+ N_XI64/XI14/NET33_XI64/XI14/MM2_g N_VSS_XI64/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI14/MM3 N_XI64/XI14/NET33_XI64/XI14/MM3_d N_WL<124>_XI64/XI14/MM3_g
+ N_BLN<1>_XI64/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI14/MM0 N_XI64/XI14/NET34_XI64/XI14/MM0_d N_WL<124>_XI64/XI14/MM0_g
+ N_BL<1>_XI64/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI14/MM1 N_XI64/XI14/NET33_XI64/XI14/MM1_d
+ N_XI64/XI14/NET34_XI64/XI14/MM1_g N_VSS_XI64/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI14/MM9 N_XI64/XI14/NET36_XI64/XI14/MM9_d N_WL<125>_XI64/XI14/MM9_g
+ N_BL<1>_XI64/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI14/MM6 N_XI64/XI14/NET35_XI64/XI14/MM6_d
+ N_XI64/XI14/NET36_XI64/XI14/MM6_g N_VSS_XI64/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI14/MM7 N_XI64/XI14/NET36_XI64/XI14/MM7_d
+ N_XI64/XI14/NET35_XI64/XI14/MM7_g N_VSS_XI64/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI14/MM8 N_XI64/XI14/NET35_XI64/XI14/MM8_d N_WL<125>_XI64/XI14/MM8_g
+ N_BLN<1>_XI64/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI14/MM5 N_XI64/XI14/NET34_XI64/XI14/MM5_d
+ N_XI64/XI14/NET33_XI64/XI14/MM5_g N_VDD_XI64/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI14/MM4 N_XI64/XI14/NET33_XI64/XI14/MM4_d
+ N_XI64/XI14/NET34_XI64/XI14/MM4_g N_VDD_XI64/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI14/MM10 N_XI64/XI14/NET35_XI64/XI14/MM10_d
+ N_XI64/XI14/NET36_XI64/XI14/MM10_g N_VDD_XI64/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI14/MM11 N_XI64/XI14/NET36_XI64/XI14/MM11_d
+ N_XI64/XI14/NET35_XI64/XI14/MM11_g N_VDD_XI64/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI15/MM2 N_XI64/XI15/NET34_XI64/XI15/MM2_d
+ N_XI64/XI15/NET33_XI64/XI15/MM2_g N_VSS_XI64/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI15/MM3 N_XI64/XI15/NET33_XI64/XI15/MM3_d N_WL<124>_XI64/XI15/MM3_g
+ N_BLN<0>_XI64/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI15/MM0 N_XI64/XI15/NET34_XI64/XI15/MM0_d N_WL<124>_XI64/XI15/MM0_g
+ N_BL<0>_XI64/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI15/MM1 N_XI64/XI15/NET33_XI64/XI15/MM1_d
+ N_XI64/XI15/NET34_XI64/XI15/MM1_g N_VSS_XI64/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI15/MM9 N_XI64/XI15/NET36_XI64/XI15/MM9_d N_WL<125>_XI64/XI15/MM9_g
+ N_BL<0>_XI64/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI15/MM6 N_XI64/XI15/NET35_XI64/XI15/MM6_d
+ N_XI64/XI15/NET36_XI64/XI15/MM6_g N_VSS_XI64/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI15/MM7 N_XI64/XI15/NET36_XI64/XI15/MM7_d
+ N_XI64/XI15/NET35_XI64/XI15/MM7_g N_VSS_XI64/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI64/XI15/MM8 N_XI64/XI15/NET35_XI64/XI15/MM8_d N_WL<125>_XI64/XI15/MM8_g
+ N_BLN<0>_XI64/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI64/XI15/MM5 N_XI64/XI15/NET34_XI64/XI15/MM5_d
+ N_XI64/XI15/NET33_XI64/XI15/MM5_g N_VDD_XI64/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI15/MM4 N_XI64/XI15/NET33_XI64/XI15/MM4_d
+ N_XI64/XI15/NET34_XI64/XI15/MM4_g N_VDD_XI64/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI15/MM10 N_XI64/XI15/NET35_XI64/XI15/MM10_d
+ N_XI64/XI15/NET36_XI64/XI15/MM10_g N_VDD_XI64/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI64/XI15/MM11 N_XI64/XI15/NET36_XI64/XI15/MM11_d
+ N_XI64/XI15/NET35_XI64/XI15/MM11_g N_VDD_XI64/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI0/MM2 N_XI65/XI0/NET34_XI65/XI0/MM2_d N_XI65/XI0/NET33_XI65/XI0/MM2_g
+ N_VSS_XI65/XI0/MM2_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI0/MM3 N_XI65/XI0/NET33_XI65/XI0/MM3_d N_WL<126>_XI65/XI0/MM3_g
+ N_BLN<15>_XI65/XI0/MM3_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI0/MM0 N_XI65/XI0/NET34_XI65/XI0/MM0_d N_WL<126>_XI65/XI0/MM0_g
+ N_BL<15>_XI65/XI0/MM0_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI0/MM1 N_XI65/XI0/NET33_XI65/XI0/MM1_d N_XI65/XI0/NET34_XI65/XI0/MM1_g
+ N_VSS_XI65/XI0/MM1_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI0/MM9 N_XI65/XI0/NET36_XI65/XI0/MM9_d N_WL<127>_XI65/XI0/MM9_g
+ N_BL<15>_XI65/XI0/MM9_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI0/MM6 N_XI65/XI0/NET35_XI65/XI0/MM6_d N_XI65/XI0/NET36_XI65/XI0/MM6_g
+ N_VSS_XI65/XI0/MM6_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI0/MM7 N_XI65/XI0/NET36_XI65/XI0/MM7_d N_XI65/XI0/NET35_XI65/XI0/MM7_g
+ N_VSS_XI65/XI0/MM7_s N_VSS_XI0/XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI0/MM8 N_XI65/XI0/NET35_XI65/XI0/MM8_d N_WL<127>_XI65/XI0/MM8_g
+ N_BLN<15>_XI65/XI0/MM8_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI0/MM5 N_XI65/XI0/NET34_XI65/XI0/MM5_d N_XI65/XI0/NET33_XI65/XI0/MM5_g
+ N_VDD_XI65/XI0/MM5_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI0/MM4 N_XI65/XI0/NET33_XI65/XI0/MM4_d N_XI65/XI0/NET34_XI65/XI0/MM4_g
+ N_VDD_XI65/XI0/MM4_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI0/MM10 N_XI65/XI0/NET35_XI65/XI0/MM10_d N_XI65/XI0/NET36_XI65/XI0/MM10_g
+ N_VDD_XI65/XI0/MM10_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI0/MM11 N_XI65/XI0/NET36_XI65/XI0/MM11_d N_XI65/XI0/NET35_XI65/XI0/MM11_g
+ N_VDD_XI65/XI0/MM11_s N_VDD_XI0/XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI1/MM2 N_XI65/XI1/NET34_XI65/XI1/MM2_d N_XI65/XI1/NET33_XI65/XI1/MM2_g
+ N_VSS_XI65/XI1/MM2_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI1/MM3 N_XI65/XI1/NET33_XI65/XI1/MM3_d N_WL<126>_XI65/XI1/MM3_g
+ N_BLN<14>_XI65/XI1/MM3_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI1/MM0 N_XI65/XI1/NET34_XI65/XI1/MM0_d N_WL<126>_XI65/XI1/MM0_g
+ N_BL<14>_XI65/XI1/MM0_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI1/MM1 N_XI65/XI1/NET33_XI65/XI1/MM1_d N_XI65/XI1/NET34_XI65/XI1/MM1_g
+ N_VSS_XI65/XI1/MM1_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI1/MM9 N_XI65/XI1/NET36_XI65/XI1/MM9_d N_WL<127>_XI65/XI1/MM9_g
+ N_BL<14>_XI65/XI1/MM9_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI1/MM6 N_XI65/XI1/NET35_XI65/XI1/MM6_d N_XI65/XI1/NET36_XI65/XI1/MM6_g
+ N_VSS_XI65/XI1/MM6_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI1/MM7 N_XI65/XI1/NET36_XI65/XI1/MM7_d N_XI65/XI1/NET35_XI65/XI1/MM7_g
+ N_VSS_XI65/XI1/MM7_s N_VSS_XI0/XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI1/MM8 N_XI65/XI1/NET35_XI65/XI1/MM8_d N_WL<127>_XI65/XI1/MM8_g
+ N_BLN<14>_XI65/XI1/MM8_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI1/MM5 N_XI65/XI1/NET34_XI65/XI1/MM5_d N_XI65/XI1/NET33_XI65/XI1/MM5_g
+ N_VDD_XI65/XI1/MM5_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI1/MM4 N_XI65/XI1/NET33_XI65/XI1/MM4_d N_XI65/XI1/NET34_XI65/XI1/MM4_g
+ N_VDD_XI65/XI1/MM4_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI1/MM10 N_XI65/XI1/NET35_XI65/XI1/MM10_d N_XI65/XI1/NET36_XI65/XI1/MM10_g
+ N_VDD_XI65/XI1/MM10_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI1/MM11 N_XI65/XI1/NET36_XI65/XI1/MM11_d N_XI65/XI1/NET35_XI65/XI1/MM11_g
+ N_VDD_XI65/XI1/MM11_s N_VDD_XI0/XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI2/MM2 N_XI65/XI2/NET34_XI65/XI2/MM2_d N_XI65/XI2/NET33_XI65/XI2/MM2_g
+ N_VSS_XI65/XI2/MM2_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI2/MM3 N_XI65/XI2/NET33_XI65/XI2/MM3_d N_WL<126>_XI65/XI2/MM3_g
+ N_BLN<13>_XI65/XI2/MM3_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI2/MM0 N_XI65/XI2/NET34_XI65/XI2/MM0_d N_WL<126>_XI65/XI2/MM0_g
+ N_BL<13>_XI65/XI2/MM0_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI2/MM1 N_XI65/XI2/NET33_XI65/XI2/MM1_d N_XI65/XI2/NET34_XI65/XI2/MM1_g
+ N_VSS_XI65/XI2/MM1_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI2/MM9 N_XI65/XI2/NET36_XI65/XI2/MM9_d N_WL<127>_XI65/XI2/MM9_g
+ N_BL<13>_XI65/XI2/MM9_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI2/MM6 N_XI65/XI2/NET35_XI65/XI2/MM6_d N_XI65/XI2/NET36_XI65/XI2/MM6_g
+ N_VSS_XI65/XI2/MM6_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI2/MM7 N_XI65/XI2/NET36_XI65/XI2/MM7_d N_XI65/XI2/NET35_XI65/XI2/MM7_g
+ N_VSS_XI65/XI2/MM7_s N_VSS_XI0/XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI2/MM8 N_XI65/XI2/NET35_XI65/XI2/MM8_d N_WL<127>_XI65/XI2/MM8_g
+ N_BLN<13>_XI65/XI2/MM8_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI2/MM5 N_XI65/XI2/NET34_XI65/XI2/MM5_d N_XI65/XI2/NET33_XI65/XI2/MM5_g
+ N_VDD_XI65/XI2/MM5_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI2/MM4 N_XI65/XI2/NET33_XI65/XI2/MM4_d N_XI65/XI2/NET34_XI65/XI2/MM4_g
+ N_VDD_XI65/XI2/MM4_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI2/MM10 N_XI65/XI2/NET35_XI65/XI2/MM10_d N_XI65/XI2/NET36_XI65/XI2/MM10_g
+ N_VDD_XI65/XI2/MM10_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI2/MM11 N_XI65/XI2/NET36_XI65/XI2/MM11_d N_XI65/XI2/NET35_XI65/XI2/MM11_g
+ N_VDD_XI65/XI2/MM11_s N_VDD_XI0/XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI3/MM2 N_XI65/XI3/NET34_XI65/XI3/MM2_d N_XI65/XI3/NET33_XI65/XI3/MM2_g
+ N_VSS_XI65/XI3/MM2_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI3/MM3 N_XI65/XI3/NET33_XI65/XI3/MM3_d N_WL<126>_XI65/XI3/MM3_g
+ N_BLN<12>_XI65/XI3/MM3_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI3/MM0 N_XI65/XI3/NET34_XI65/XI3/MM0_d N_WL<126>_XI65/XI3/MM0_g
+ N_BL<12>_XI65/XI3/MM0_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI3/MM1 N_XI65/XI3/NET33_XI65/XI3/MM1_d N_XI65/XI3/NET34_XI65/XI3/MM1_g
+ N_VSS_XI65/XI3/MM1_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI3/MM9 N_XI65/XI3/NET36_XI65/XI3/MM9_d N_WL<127>_XI65/XI3/MM9_g
+ N_BL<12>_XI65/XI3/MM9_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI3/MM6 N_XI65/XI3/NET35_XI65/XI3/MM6_d N_XI65/XI3/NET36_XI65/XI3/MM6_g
+ N_VSS_XI65/XI3/MM6_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI3/MM7 N_XI65/XI3/NET36_XI65/XI3/MM7_d N_XI65/XI3/NET35_XI65/XI3/MM7_g
+ N_VSS_XI65/XI3/MM7_s N_VSS_XI0/XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI3/MM8 N_XI65/XI3/NET35_XI65/XI3/MM8_d N_WL<127>_XI65/XI3/MM8_g
+ N_BLN<12>_XI65/XI3/MM8_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI3/MM5 N_XI65/XI3/NET34_XI65/XI3/MM5_d N_XI65/XI3/NET33_XI65/XI3/MM5_g
+ N_VDD_XI65/XI3/MM5_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI3/MM4 N_XI65/XI3/NET33_XI65/XI3/MM4_d N_XI65/XI3/NET34_XI65/XI3/MM4_g
+ N_VDD_XI65/XI3/MM4_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI3/MM10 N_XI65/XI3/NET35_XI65/XI3/MM10_d N_XI65/XI3/NET36_XI65/XI3/MM10_g
+ N_VDD_XI65/XI3/MM10_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI3/MM11 N_XI65/XI3/NET36_XI65/XI3/MM11_d N_XI65/XI3/NET35_XI65/XI3/MM11_g
+ N_VDD_XI65/XI3/MM11_s N_VDD_XI0/XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI4/MM2 N_XI65/XI4/NET34_XI65/XI4/MM2_d N_XI65/XI4/NET33_XI65/XI4/MM2_g
+ N_VSS_XI65/XI4/MM2_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI4/MM3 N_XI65/XI4/NET33_XI65/XI4/MM3_d N_WL<126>_XI65/XI4/MM3_g
+ N_BLN<11>_XI65/XI4/MM3_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI4/MM0 N_XI65/XI4/NET34_XI65/XI4/MM0_d N_WL<126>_XI65/XI4/MM0_g
+ N_BL<11>_XI65/XI4/MM0_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI4/MM1 N_XI65/XI4/NET33_XI65/XI4/MM1_d N_XI65/XI4/NET34_XI65/XI4/MM1_g
+ N_VSS_XI65/XI4/MM1_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI4/MM9 N_XI65/XI4/NET36_XI65/XI4/MM9_d N_WL<127>_XI65/XI4/MM9_g
+ N_BL<11>_XI65/XI4/MM9_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI4/MM6 N_XI65/XI4/NET35_XI65/XI4/MM6_d N_XI65/XI4/NET36_XI65/XI4/MM6_g
+ N_VSS_XI65/XI4/MM6_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI4/MM7 N_XI65/XI4/NET36_XI65/XI4/MM7_d N_XI65/XI4/NET35_XI65/XI4/MM7_g
+ N_VSS_XI65/XI4/MM7_s N_VSS_XI0/XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI4/MM8 N_XI65/XI4/NET35_XI65/XI4/MM8_d N_WL<127>_XI65/XI4/MM8_g
+ N_BLN<11>_XI65/XI4/MM8_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI4/MM5 N_XI65/XI4/NET34_XI65/XI4/MM5_d N_XI65/XI4/NET33_XI65/XI4/MM5_g
+ N_VDD_XI65/XI4/MM5_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI4/MM4 N_XI65/XI4/NET33_XI65/XI4/MM4_d N_XI65/XI4/NET34_XI65/XI4/MM4_g
+ N_VDD_XI65/XI4/MM4_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI4/MM10 N_XI65/XI4/NET35_XI65/XI4/MM10_d N_XI65/XI4/NET36_XI65/XI4/MM10_g
+ N_VDD_XI65/XI4/MM10_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI4/MM11 N_XI65/XI4/NET36_XI65/XI4/MM11_d N_XI65/XI4/NET35_XI65/XI4/MM11_g
+ N_VDD_XI65/XI4/MM11_s N_VDD_XI0/XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI5/MM2 N_XI65/XI5/NET34_XI65/XI5/MM2_d N_XI65/XI5/NET33_XI65/XI5/MM2_g
+ N_VSS_XI65/XI5/MM2_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI5/MM3 N_XI65/XI5/NET33_XI65/XI5/MM3_d N_WL<126>_XI65/XI5/MM3_g
+ N_BLN<10>_XI65/XI5/MM3_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI5/MM0 N_XI65/XI5/NET34_XI65/XI5/MM0_d N_WL<126>_XI65/XI5/MM0_g
+ N_BL<10>_XI65/XI5/MM0_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI5/MM1 N_XI65/XI5/NET33_XI65/XI5/MM1_d N_XI65/XI5/NET34_XI65/XI5/MM1_g
+ N_VSS_XI65/XI5/MM1_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI5/MM9 N_XI65/XI5/NET36_XI65/XI5/MM9_d N_WL<127>_XI65/XI5/MM9_g
+ N_BL<10>_XI65/XI5/MM9_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI5/MM6 N_XI65/XI5/NET35_XI65/XI5/MM6_d N_XI65/XI5/NET36_XI65/XI5/MM6_g
+ N_VSS_XI65/XI5/MM6_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI5/MM7 N_XI65/XI5/NET36_XI65/XI5/MM7_d N_XI65/XI5/NET35_XI65/XI5/MM7_g
+ N_VSS_XI65/XI5/MM7_s N_VSS_XI0/XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI5/MM8 N_XI65/XI5/NET35_XI65/XI5/MM8_d N_WL<127>_XI65/XI5/MM8_g
+ N_BLN<10>_XI65/XI5/MM8_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI5/MM5 N_XI65/XI5/NET34_XI65/XI5/MM5_d N_XI65/XI5/NET33_XI65/XI5/MM5_g
+ N_VDD_XI65/XI5/MM5_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI5/MM4 N_XI65/XI5/NET33_XI65/XI5/MM4_d N_XI65/XI5/NET34_XI65/XI5/MM4_g
+ N_VDD_XI65/XI5/MM4_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI5/MM10 N_XI65/XI5/NET35_XI65/XI5/MM10_d N_XI65/XI5/NET36_XI65/XI5/MM10_g
+ N_VDD_XI65/XI5/MM10_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI5/MM11 N_XI65/XI5/NET36_XI65/XI5/MM11_d N_XI65/XI5/NET35_XI65/XI5/MM11_g
+ N_VDD_XI65/XI5/MM11_s N_VDD_XI0/XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI6/MM2 N_XI65/XI6/NET34_XI65/XI6/MM2_d N_XI65/XI6/NET33_XI65/XI6/MM2_g
+ N_VSS_XI65/XI6/MM2_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM3 N_XI65/XI6/NET33_XI65/XI6/MM3_d N_WL<126>_XI65/XI6/MM3_g
+ N_BLN<9>_XI65/XI6/MM3_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM0 N_XI65/XI6/NET34_XI65/XI6/MM0_d N_WL<126>_XI65/XI6/MM0_g
+ N_BL<9>_XI65/XI6/MM0_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM1 N_XI65/XI6/NET33_XI65/XI6/MM1_d N_XI65/XI6/NET34_XI65/XI6/MM1_g
+ N_VSS_XI65/XI6/MM1_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM9 N_XI65/XI6/NET36_XI65/XI6/MM9_d N_WL<127>_XI65/XI6/MM9_g
+ N_BL<9>_XI65/XI6/MM9_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM6 N_XI65/XI6/NET35_XI65/XI6/MM6_d N_XI65/XI6/NET36_XI65/XI6/MM6_g
+ N_VSS_XI65/XI6/MM6_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM7 N_XI65/XI6/NET36_XI65/XI6/MM7_d N_XI65/XI6/NET35_XI65/XI6/MM7_g
+ N_VSS_XI65/XI6/MM7_s N_VSS_XI0/XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM8 N_XI65/XI6/NET35_XI65/XI6/MM8_d N_WL<127>_XI65/XI6/MM8_g
+ N_BLN<9>_XI65/XI6/MM8_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI6/MM5 N_XI65/XI6/NET34_XI65/XI6/MM5_d N_XI65/XI6/NET33_XI65/XI6/MM5_g
+ N_VDD_XI65/XI6/MM5_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI6/MM4 N_XI65/XI6/NET33_XI65/XI6/MM4_d N_XI65/XI6/NET34_XI65/XI6/MM4_g
+ N_VDD_XI65/XI6/MM4_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI6/MM10 N_XI65/XI6/NET35_XI65/XI6/MM10_d N_XI65/XI6/NET36_XI65/XI6/MM10_g
+ N_VDD_XI65/XI6/MM10_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI6/MM11 N_XI65/XI6/NET36_XI65/XI6/MM11_d N_XI65/XI6/NET35_XI65/XI6/MM11_g
+ N_VDD_XI65/XI6/MM11_s N_VDD_XI0/XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI7/MM2 N_XI65/XI7/NET34_XI65/XI7/MM2_d N_XI65/XI7/NET33_XI65/XI7/MM2_g
+ N_VSS_XI65/XI7/MM2_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM3 N_XI65/XI7/NET33_XI65/XI7/MM3_d N_WL<126>_XI65/XI7/MM3_g
+ N_BLN<8>_XI65/XI7/MM3_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM0 N_XI65/XI7/NET34_XI65/XI7/MM0_d N_WL<126>_XI65/XI7/MM0_g
+ N_BL<8>_XI65/XI7/MM0_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM1 N_XI65/XI7/NET33_XI65/XI7/MM1_d N_XI65/XI7/NET34_XI65/XI7/MM1_g
+ N_VSS_XI65/XI7/MM1_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM9 N_XI65/XI7/NET36_XI65/XI7/MM9_d N_WL<127>_XI65/XI7/MM9_g
+ N_BL<8>_XI65/XI7/MM9_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM6 N_XI65/XI7/NET35_XI65/XI7/MM6_d N_XI65/XI7/NET36_XI65/XI7/MM6_g
+ N_VSS_XI65/XI7/MM6_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM7 N_XI65/XI7/NET36_XI65/XI7/MM7_d N_XI65/XI7/NET35_XI65/XI7/MM7_g
+ N_VSS_XI65/XI7/MM7_s N_VSS_XI0/XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM8 N_XI65/XI7/NET35_XI65/XI7/MM8_d N_WL<127>_XI65/XI7/MM8_g
+ N_BLN<8>_XI65/XI7/MM8_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI7/MM5 N_XI65/XI7/NET34_XI65/XI7/MM5_d N_XI65/XI7/NET33_XI65/XI7/MM5_g
+ N_VDD_XI65/XI7/MM5_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI7/MM4 N_XI65/XI7/NET33_XI65/XI7/MM4_d N_XI65/XI7/NET34_XI65/XI7/MM4_g
+ N_VDD_XI65/XI7/MM4_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI7/MM10 N_XI65/XI7/NET35_XI65/XI7/MM10_d N_XI65/XI7/NET36_XI65/XI7/MM10_g
+ N_VDD_XI65/XI7/MM10_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI7/MM11 N_XI65/XI7/NET36_XI65/XI7/MM11_d N_XI65/XI7/NET35_XI65/XI7/MM11_g
+ N_VDD_XI65/XI7/MM11_s N_VDD_XI0/XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI8/MM2 N_XI65/XI8/NET34_XI65/XI8/MM2_d N_XI65/XI8/NET33_XI65/XI8/MM2_g
+ N_VSS_XI65/XI8/MM2_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM3 N_XI65/XI8/NET33_XI65/XI8/MM3_d N_WL<126>_XI65/XI8/MM3_g
+ N_BLN<7>_XI65/XI8/MM3_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM0 N_XI65/XI8/NET34_XI65/XI8/MM0_d N_WL<126>_XI65/XI8/MM0_g
+ N_BL<7>_XI65/XI8/MM0_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM1 N_XI65/XI8/NET33_XI65/XI8/MM1_d N_XI65/XI8/NET34_XI65/XI8/MM1_g
+ N_VSS_XI65/XI8/MM1_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM9 N_XI65/XI8/NET36_XI65/XI8/MM9_d N_WL<127>_XI65/XI8/MM9_g
+ N_BL<7>_XI65/XI8/MM9_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM6 N_XI65/XI8/NET35_XI65/XI8/MM6_d N_XI65/XI8/NET36_XI65/XI8/MM6_g
+ N_VSS_XI65/XI8/MM6_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM7 N_XI65/XI8/NET36_XI65/XI8/MM7_d N_XI65/XI8/NET35_XI65/XI8/MM7_g
+ N_VSS_XI65/XI8/MM7_s N_VSS_XI0/XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM8 N_XI65/XI8/NET35_XI65/XI8/MM8_d N_WL<127>_XI65/XI8/MM8_g
+ N_BLN<7>_XI65/XI8/MM8_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI8/MM5 N_XI65/XI8/NET34_XI65/XI8/MM5_d N_XI65/XI8/NET33_XI65/XI8/MM5_g
+ N_VDD_XI65/XI8/MM5_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI8/MM4 N_XI65/XI8/NET33_XI65/XI8/MM4_d N_XI65/XI8/NET34_XI65/XI8/MM4_g
+ N_VDD_XI65/XI8/MM4_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI8/MM10 N_XI65/XI8/NET35_XI65/XI8/MM10_d N_XI65/XI8/NET36_XI65/XI8/MM10_g
+ N_VDD_XI65/XI8/MM10_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI8/MM11 N_XI65/XI8/NET36_XI65/XI8/MM11_d N_XI65/XI8/NET35_XI65/XI8/MM11_g
+ N_VDD_XI65/XI8/MM11_s N_VDD_XI0/XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI9/MM2 N_XI65/XI9/NET34_XI65/XI9/MM2_d N_XI65/XI9/NET33_XI65/XI9/MM2_g
+ N_VSS_XI65/XI9/MM2_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM3 N_XI65/XI9/NET33_XI65/XI9/MM3_d N_WL<126>_XI65/XI9/MM3_g
+ N_BLN<6>_XI65/XI9/MM3_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM0 N_XI65/XI9/NET34_XI65/XI9/MM0_d N_WL<126>_XI65/XI9/MM0_g
+ N_BL<6>_XI65/XI9/MM0_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM1 N_XI65/XI9/NET33_XI65/XI9/MM1_d N_XI65/XI9/NET34_XI65/XI9/MM1_g
+ N_VSS_XI65/XI9/MM1_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM9 N_XI65/XI9/NET36_XI65/XI9/MM9_d N_WL<127>_XI65/XI9/MM9_g
+ N_BL<6>_XI65/XI9/MM9_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM6 N_XI65/XI9/NET35_XI65/XI9/MM6_d N_XI65/XI9/NET36_XI65/XI9/MM6_g
+ N_VSS_XI65/XI9/MM6_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM7 N_XI65/XI9/NET36_XI65/XI9/MM7_d N_XI65/XI9/NET35_XI65/XI9/MM7_g
+ N_VSS_XI65/XI9/MM7_s N_VSS_XI0/XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM8 N_XI65/XI9/NET35_XI65/XI9/MM8_d N_WL<127>_XI65/XI9/MM8_g
+ N_BLN<6>_XI65/XI9/MM8_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI9/MM5 N_XI65/XI9/NET34_XI65/XI9/MM5_d N_XI65/XI9/NET33_XI65/XI9/MM5_g
+ N_VDD_XI65/XI9/MM5_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI9/MM4 N_XI65/XI9/NET33_XI65/XI9/MM4_d N_XI65/XI9/NET34_XI65/XI9/MM4_g
+ N_VDD_XI65/XI9/MM4_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI9/MM10 N_XI65/XI9/NET35_XI65/XI9/MM10_d N_XI65/XI9/NET36_XI65/XI9/MM10_g
+ N_VDD_XI65/XI9/MM10_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI9/MM11 N_XI65/XI9/NET36_XI65/XI9/MM11_d N_XI65/XI9/NET35_XI65/XI9/MM11_g
+ N_VDD_XI65/XI9/MM11_s N_VDD_XI0/XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI10/MM2 N_XI65/XI10/NET34_XI65/XI10/MM2_d
+ N_XI65/XI10/NET33_XI65/XI10/MM2_g N_VSS_XI65/XI10/MM2_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI10/MM3 N_XI65/XI10/NET33_XI65/XI10/MM3_d N_WL<126>_XI65/XI10/MM3_g
+ N_BLN<5>_XI65/XI10/MM3_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI10/MM0 N_XI65/XI10/NET34_XI65/XI10/MM0_d N_WL<126>_XI65/XI10/MM0_g
+ N_BL<5>_XI65/XI10/MM0_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI10/MM1 N_XI65/XI10/NET33_XI65/XI10/MM1_d
+ N_XI65/XI10/NET34_XI65/XI10/MM1_g N_VSS_XI65/XI10/MM1_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI10/MM9 N_XI65/XI10/NET36_XI65/XI10/MM9_d N_WL<127>_XI65/XI10/MM9_g
+ N_BL<5>_XI65/XI10/MM9_s N_VSS_XI0/XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI10/MM6 N_XI65/XI10/NET35_XI65/XI10/MM6_d
+ N_XI65/XI10/NET36_XI65/XI10/MM6_g N_VSS_XI65/XI10/MM6_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI10/MM7 N_XI65/XI10/NET36_XI65/XI10/MM7_d
+ N_XI65/XI10/NET35_XI65/XI10/MM7_g N_VSS_XI65/XI10/MM7_s N_VSS_XI0/XI9/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI10/MM8 N_XI65/XI10/NET35_XI65/XI10/MM8_d N_WL<127>_XI65/XI10/MM8_g
+ N_BLN<5>_XI65/XI10/MM8_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI10/MM5 N_XI65/XI10/NET34_XI65/XI10/MM5_d
+ N_XI65/XI10/NET33_XI65/XI10/MM5_g N_VDD_XI65/XI10/MM5_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI10/MM4 N_XI65/XI10/NET33_XI65/XI10/MM4_d
+ N_XI65/XI10/NET34_XI65/XI10/MM4_g N_VDD_XI65/XI10/MM4_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI10/MM10 N_XI65/XI10/NET35_XI65/XI10/MM10_d
+ N_XI65/XI10/NET36_XI65/XI10/MM10_g N_VDD_XI65/XI10/MM10_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI10/MM11 N_XI65/XI10/NET36_XI65/XI10/MM11_d
+ N_XI65/XI10/NET35_XI65/XI10/MM11_g N_VDD_XI65/XI10/MM11_s N_VDD_XI0/XI10/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI11/MM2 N_XI65/XI11/NET34_XI65/XI11/MM2_d
+ N_XI65/XI11/NET33_XI65/XI11/MM2_g N_VSS_XI65/XI11/MM2_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI11/MM3 N_XI65/XI11/NET33_XI65/XI11/MM3_d N_WL<126>_XI65/XI11/MM3_g
+ N_BLN<4>_XI65/XI11/MM3_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI11/MM0 N_XI65/XI11/NET34_XI65/XI11/MM0_d N_WL<126>_XI65/XI11/MM0_g
+ N_BL<4>_XI65/XI11/MM0_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI11/MM1 N_XI65/XI11/NET33_XI65/XI11/MM1_d
+ N_XI65/XI11/NET34_XI65/XI11/MM1_g N_VSS_XI65/XI11/MM1_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI11/MM9 N_XI65/XI11/NET36_XI65/XI11/MM9_d N_WL<127>_XI65/XI11/MM9_g
+ N_BL<4>_XI65/XI11/MM9_s N_VSS_XI0/XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI11/MM6 N_XI65/XI11/NET35_XI65/XI11/MM6_d
+ N_XI65/XI11/NET36_XI65/XI11/MM6_g N_VSS_XI65/XI11/MM6_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI11/MM7 N_XI65/XI11/NET36_XI65/XI11/MM7_d
+ N_XI65/XI11/NET35_XI65/XI11/MM7_g N_VSS_XI65/XI11/MM7_s N_VSS_XI0/XI10/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI11/MM8 N_XI65/XI11/NET35_XI65/XI11/MM8_d N_WL<127>_XI65/XI11/MM8_g
+ N_BLN<4>_XI65/XI11/MM8_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI11/MM5 N_XI65/XI11/NET34_XI65/XI11/MM5_d
+ N_XI65/XI11/NET33_XI65/XI11/MM5_g N_VDD_XI65/XI11/MM5_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI11/MM4 N_XI65/XI11/NET33_XI65/XI11/MM4_d
+ N_XI65/XI11/NET34_XI65/XI11/MM4_g N_VDD_XI65/XI11/MM4_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI11/MM10 N_XI65/XI11/NET35_XI65/XI11/MM10_d
+ N_XI65/XI11/NET36_XI65/XI11/MM10_g N_VDD_XI65/XI11/MM10_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI11/MM11 N_XI65/XI11/NET36_XI65/XI11/MM11_d
+ N_XI65/XI11/NET35_XI65/XI11/MM11_g N_VDD_XI65/XI11/MM11_s N_VDD_XI0/XI11/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI12/MM2 N_XI65/XI12/NET34_XI65/XI12/MM2_d
+ N_XI65/XI12/NET33_XI65/XI12/MM2_g N_VSS_XI65/XI12/MM2_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI12/MM3 N_XI65/XI12/NET33_XI65/XI12/MM3_d N_WL<126>_XI65/XI12/MM3_g
+ N_BLN<3>_XI65/XI12/MM3_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI12/MM0 N_XI65/XI12/NET34_XI65/XI12/MM0_d N_WL<126>_XI65/XI12/MM0_g
+ N_BL<3>_XI65/XI12/MM0_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI12/MM1 N_XI65/XI12/NET33_XI65/XI12/MM1_d
+ N_XI65/XI12/NET34_XI65/XI12/MM1_g N_VSS_XI65/XI12/MM1_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI12/MM9 N_XI65/XI12/NET36_XI65/XI12/MM9_d N_WL<127>_XI65/XI12/MM9_g
+ N_BL<3>_XI65/XI12/MM9_s N_VSS_XI0/XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI12/MM6 N_XI65/XI12/NET35_XI65/XI12/MM6_d
+ N_XI65/XI12/NET36_XI65/XI12/MM6_g N_VSS_XI65/XI12/MM6_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI12/MM7 N_XI65/XI12/NET36_XI65/XI12/MM7_d
+ N_XI65/XI12/NET35_XI65/XI12/MM7_g N_VSS_XI65/XI12/MM7_s N_VSS_XI0/XI11/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI12/MM8 N_XI65/XI12/NET35_XI65/XI12/MM8_d N_WL<127>_XI65/XI12/MM8_g
+ N_BLN<3>_XI65/XI12/MM8_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI12/MM5 N_XI65/XI12/NET34_XI65/XI12/MM5_d
+ N_XI65/XI12/NET33_XI65/XI12/MM5_g N_VDD_XI65/XI12/MM5_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI12/MM4 N_XI65/XI12/NET33_XI65/XI12/MM4_d
+ N_XI65/XI12/NET34_XI65/XI12/MM4_g N_VDD_XI65/XI12/MM4_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI12/MM10 N_XI65/XI12/NET35_XI65/XI12/MM10_d
+ N_XI65/XI12/NET36_XI65/XI12/MM10_g N_VDD_XI65/XI12/MM10_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI12/MM11 N_XI65/XI12/NET36_XI65/XI12/MM11_d
+ N_XI65/XI12/NET35_XI65/XI12/MM11_g N_VDD_XI65/XI12/MM11_s N_VDD_XI0/XI12/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI13/MM2 N_XI65/XI13/NET34_XI65/XI13/MM2_d
+ N_XI65/XI13/NET33_XI65/XI13/MM2_g N_VSS_XI65/XI13/MM2_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI13/MM3 N_XI65/XI13/NET33_XI65/XI13/MM3_d N_WL<126>_XI65/XI13/MM3_g
+ N_BLN<2>_XI65/XI13/MM3_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI13/MM0 N_XI65/XI13/NET34_XI65/XI13/MM0_d N_WL<126>_XI65/XI13/MM0_g
+ N_BL<2>_XI65/XI13/MM0_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI13/MM1 N_XI65/XI13/NET33_XI65/XI13/MM1_d
+ N_XI65/XI13/NET34_XI65/XI13/MM1_g N_VSS_XI65/XI13/MM1_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI13/MM9 N_XI65/XI13/NET36_XI65/XI13/MM9_d N_WL<127>_XI65/XI13/MM9_g
+ N_BL<2>_XI65/XI13/MM9_s N_VSS_XI0/XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI13/MM6 N_XI65/XI13/NET35_XI65/XI13/MM6_d
+ N_XI65/XI13/NET36_XI65/XI13/MM6_g N_VSS_XI65/XI13/MM6_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI13/MM7 N_XI65/XI13/NET36_XI65/XI13/MM7_d
+ N_XI65/XI13/NET35_XI65/XI13/MM7_g N_VSS_XI65/XI13/MM7_s N_VSS_XI0/XI12/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI13/MM8 N_XI65/XI13/NET35_XI65/XI13/MM8_d N_WL<127>_XI65/XI13/MM8_g
+ N_BLN<2>_XI65/XI13/MM8_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI13/MM5 N_XI65/XI13/NET34_XI65/XI13/MM5_d
+ N_XI65/XI13/NET33_XI65/XI13/MM5_g N_VDD_XI65/XI13/MM5_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI13/MM4 N_XI65/XI13/NET33_XI65/XI13/MM4_d
+ N_XI65/XI13/NET34_XI65/XI13/MM4_g N_VDD_XI65/XI13/MM4_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI13/MM10 N_XI65/XI13/NET35_XI65/XI13/MM10_d
+ N_XI65/XI13/NET36_XI65/XI13/MM10_g N_VDD_XI65/XI13/MM10_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI13/MM11 N_XI65/XI13/NET36_XI65/XI13/MM11_d
+ N_XI65/XI13/NET35_XI65/XI13/MM11_g N_VDD_XI65/XI13/MM11_s N_VDD_XI0/XI13/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI14/MM2 N_XI65/XI14/NET34_XI65/XI14/MM2_d
+ N_XI65/XI14/NET33_XI65/XI14/MM2_g N_VSS_XI65/XI14/MM2_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI14/MM3 N_XI65/XI14/NET33_XI65/XI14/MM3_d N_WL<126>_XI65/XI14/MM3_g
+ N_BLN<1>_XI65/XI14/MM3_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI14/MM0 N_XI65/XI14/NET34_XI65/XI14/MM0_d N_WL<126>_XI65/XI14/MM0_g
+ N_BL<1>_XI65/XI14/MM0_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI14/MM1 N_XI65/XI14/NET33_XI65/XI14/MM1_d
+ N_XI65/XI14/NET34_XI65/XI14/MM1_g N_VSS_XI65/XI14/MM1_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI14/MM9 N_XI65/XI14/NET36_XI65/XI14/MM9_d N_WL<127>_XI65/XI14/MM9_g
+ N_BL<1>_XI65/XI14/MM9_s N_VSS_XI0/XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI14/MM6 N_XI65/XI14/NET35_XI65/XI14/MM6_d
+ N_XI65/XI14/NET36_XI65/XI14/MM6_g N_VSS_XI65/XI14/MM6_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI14/MM7 N_XI65/XI14/NET36_XI65/XI14/MM7_d
+ N_XI65/XI14/NET35_XI65/XI14/MM7_g N_VSS_XI65/XI14/MM7_s N_VSS_XI0/XI13/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI14/MM8 N_XI65/XI14/NET35_XI65/XI14/MM8_d N_WL<127>_XI65/XI14/MM8_g
+ N_BLN<1>_XI65/XI14/MM8_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI14/MM5 N_XI65/XI14/NET34_XI65/XI14/MM5_d
+ N_XI65/XI14/NET33_XI65/XI14/MM5_g N_VDD_XI65/XI14/MM5_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI14/MM4 N_XI65/XI14/NET33_XI65/XI14/MM4_d
+ N_XI65/XI14/NET34_XI65/XI14/MM4_g N_VDD_XI65/XI14/MM4_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI14/MM10 N_XI65/XI14/NET35_XI65/XI14/MM10_d
+ N_XI65/XI14/NET36_XI65/XI14/MM10_g N_VDD_XI65/XI14/MM10_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI14/MM11 N_XI65/XI14/NET36_XI65/XI14/MM11_d
+ N_XI65/XI14/NET35_XI65/XI14/MM11_g N_VDD_XI65/XI14/MM11_s N_VDD_XI0/XI14/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI15/MM2 N_XI65/XI15/NET34_XI65/XI15/MM2_d
+ N_XI65/XI15/NET33_XI65/XI15/MM2_g N_VSS_XI65/XI15/MM2_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI15/MM3 N_XI65/XI15/NET33_XI65/XI15/MM3_d N_WL<126>_XI65/XI15/MM3_g
+ N_BLN<0>_XI65/XI15/MM3_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI15/MM0 N_XI65/XI15/NET34_XI65/XI15/MM0_d N_WL<126>_XI65/XI15/MM0_g
+ N_BL<0>_XI65/XI15/MM0_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI15/MM1 N_XI65/XI15/NET33_XI65/XI15/MM1_d
+ N_XI65/XI15/NET34_XI65/XI15/MM1_g N_VSS_XI65/XI15/MM1_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI15/MM9 N_XI65/XI15/NET36_XI65/XI15/MM9_d N_WL<127>_XI65/XI15/MM9_g
+ N_BL<0>_XI65/XI15/MM9_s N_VSS_XI0/XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI15/MM6 N_XI65/XI15/NET35_XI65/XI15/MM6_d
+ N_XI65/XI15/NET36_XI65/XI15/MM6_g N_VSS_XI65/XI15/MM6_s N_VSS_XI0/XI15/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI15/MM7 N_XI65/XI15/NET36_XI65/XI15/MM7_d
+ N_XI65/XI15/NET35_XI65/XI15/MM7_g N_VSS_XI65/XI15/MM7_s N_VSS_XI0/XI14/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI65/XI15/MM8 N_XI65/XI15/NET35_XI65/XI15/MM8_d N_WL<127>_XI65/XI15/MM8_g
+ N_BLN<0>_XI65/XI15/MM8_s N_VSS_XI0/XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
mXI65/XI15/MM5 N_XI65/XI15/NET34_XI65/XI15/MM5_d
+ N_XI65/XI15/NET33_XI65/XI15/MM5_g N_VDD_XI65/XI15/MM5_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI15/MM4 N_XI65/XI15/NET33_XI65/XI15/MM4_d
+ N_XI65/XI15/NET34_XI65/XI15/MM4_g N_VDD_XI65/XI15/MM4_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI15/MM10 N_XI65/XI15/NET35_XI65/XI15/MM10_d
+ N_XI65/XI15/NET36_XI65/XI15/MM10_g N_VDD_XI65/XI15/MM10_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI65/XI15/MM11 N_XI65/XI15/NET36_XI65/XI15/MM11_d
+ N_XI65/XI15/NET35_XI65/XI15/MM11_g N_VDD_XI65/XI15/MM11_s N_VDD_XI0/XI15/MM5_b
+ PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
*
.include "netlist.sp.SRAM_ARRAY_1.pxi"
*
.ends
*
*
