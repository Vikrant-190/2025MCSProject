* SPICE NETLIST
***************************************

.SUBCKT test_inv3
** N=0 EP=0 IP=0 FDC=0
.ENDS
***************************************
