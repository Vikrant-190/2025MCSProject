* File: netlist.sp
* Created: Fri Jun 13 10:04:52 2025
* Program "Calibre xRC"
* Version "v2019.2_26.18"
* 
.include "netlist.sp.pex"
.subckt sram_16b_2  BL<15> BLN<15> BL<14> BLN<14> BL<13> BLN<13> BL<12> BLN<12>
+ BL<11> BLN<11> BL<10> BLN<10> BL<9> BLN<9> BL<8> BLN<8> BL<7> BLN<7> BL<6>
+ BLN<6> BL<5> BLN<5> BL<4> BLN<4> BL<3> BLN<3> BL<2> BLN<2> BL<1> BLN<1> BL<0>
+ BLN<0> VSS VDD WL0 WL1
* 
* WL1	WL1
* WL0	WL0
* VDD	VDD
* VSS	VSS
* BLN<0>	BLN<0>
* BL<0>	BL<0>
* BLN<1>	BLN<1>
* BL<1>	BL<1>
* BLN<2>	BLN<2>
* BL<2>	BL<2>
* BLN<3>	BLN<3>
* BL<3>	BL<3>
* BLN<4>	BLN<4>
* BL<4>	BL<4>
* BLN<5>	BLN<5>
* BL<5>	BL<5>
* BLN<6>	BLN<6>
* BL<6>	BL<6>
* BLN<7>	BLN<7>
* BL<7>	BL<7>
* BLN<8>	BLN<8>
* BL<8>	BL<8>
* BLN<9>	BLN<9>
* BL<9>	BL<9>
* BLN<10>	BLN<10>
* BL<10>	BL<10>
* BLN<11>	BLN<11>
* BL<11>	BL<11>
* BLN<12>	BLN<12>
* BL<12>	BL<12>
* BLN<13>	BLN<13>
* BL<13>	BL<13>
* BLN<14>	BLN<14>
* BL<14>	BL<14>
* BLN<15>	BLN<15>
* BL<15>	BL<15>
mXI0/MM2 N_XI0/NET34_XI0/MM2_d N_XI0/NET33_XI0/MM2_g N_VSS_XI0/MM2_s
+ N_VSS_XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM3 N_XI0/NET33_XI0/MM3_d N_WL0_XI0/MM3_g N_BLN<15>_XI0/MM3_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM0 N_XI0/NET34_XI0/MM0_d N_WL0_XI0/MM0_g N_BL<15>_XI0/MM0_s
+ N_VSS_XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM1 N_XI0/NET33_XI0/MM1_d N_XI0/NET34_XI0/MM1_g N_VSS_XI0/MM1_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM9 N_XI0/NET36_XI0/MM9_d N_WL1_XI0/MM9_g N_BL<15>_XI0/MM9_s
+ N_VSS_XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM6 N_XI0/NET35_XI0/MM6_d N_XI0/NET36_XI0/MM6_g N_VSS_XI0/MM6_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM7 N_XI0/NET36_XI0/MM7_d N_XI0/NET35_XI0/MM7_g N_VSS_XI0/MM7_s
+ N_VSS_XI0/MM2_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM8 N_XI0/NET35_XI0/MM8_d N_WL1_XI0/MM8_g N_BLN<15>_XI0/MM8_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI0/MM5 N_XI0/NET34_XI0/MM5_d N_XI0/NET33_XI0/MM5_g N_VDD_XI0/MM5_s
+ N_VDD_XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/MM4 N_XI0/NET33_XI0/MM4_d N_XI0/NET34_XI0/MM4_g N_VDD_XI0/MM4_s
+ N_VDD_XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/MM10 N_XI0/NET35_XI0/MM10_d N_XI0/NET36_XI0/MM10_g N_VDD_XI0/MM10_s
+ N_VDD_XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI0/MM11 N_XI0/NET36_XI0/MM11_d N_XI0/NET35_XI0/MM11_g N_VDD_XI0/MM11_s
+ N_VDD_XI0/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/MM2 N_XI1/NET34_XI1/MM2_d N_XI1/NET33_XI1/MM2_g N_VSS_XI1/MM2_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM3 N_XI1/NET33_XI1/MM3_d N_WL0_XI1/MM3_g N_BLN<14>_XI1/MM3_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM0 N_XI1/NET34_XI1/MM0_d N_WL0_XI1/MM0_g N_BL<14>_XI1/MM0_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM1 N_XI1/NET33_XI1/MM1_d N_XI1/NET34_XI1/MM1_g N_VSS_XI1/MM1_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM9 N_XI1/NET36_XI1/MM9_d N_WL1_XI1/MM9_g N_BL<14>_XI1/MM9_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM6 N_XI1/NET35_XI1/MM6_d N_XI1/NET36_XI1/MM6_g N_VSS_XI1/MM6_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM7 N_XI1/NET36_XI1/MM7_d N_XI1/NET35_XI1/MM7_g N_VSS_XI1/MM7_s
+ N_VSS_XI0/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM8 N_XI1/NET35_XI1/MM8_d N_WL1_XI1/MM8_g N_BLN<14>_XI1/MM8_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI1/MM5 N_XI1/NET34_XI1/MM5_d N_XI1/NET33_XI1/MM5_g N_VDD_XI1/MM5_s
+ N_VDD_XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/MM4 N_XI1/NET33_XI1/MM4_d N_XI1/NET34_XI1/MM4_g N_VDD_XI1/MM4_s
+ N_VDD_XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/MM10 N_XI1/NET35_XI1/MM10_d N_XI1/NET36_XI1/MM10_g N_VDD_XI1/MM10_s
+ N_VDD_XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI1/MM11 N_XI1/NET36_XI1/MM11_d N_XI1/NET35_XI1/MM11_g N_VDD_XI1/MM11_s
+ N_VDD_XI1/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI2/MM2 N_XI2/NET34_XI2/MM2_d N_XI2/NET33_XI2/MM2_g N_VSS_XI2/MM2_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM3 N_XI2/NET33_XI2/MM3_d N_WL0_XI2/MM3_g N_BLN<13>_XI2/MM3_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM0 N_XI2/NET34_XI2/MM0_d N_WL0_XI2/MM0_g N_BL<13>_XI2/MM0_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM1 N_XI2/NET33_XI2/MM1_d N_XI2/NET34_XI2/MM1_g N_VSS_XI2/MM1_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM9 N_XI2/NET36_XI2/MM9_d N_WL1_XI2/MM9_g N_BL<13>_XI2/MM9_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM6 N_XI2/NET35_XI2/MM6_d N_XI2/NET36_XI2/MM6_g N_VSS_XI2/MM6_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM7 N_XI2/NET36_XI2/MM7_d N_XI2/NET35_XI2/MM7_g N_VSS_XI2/MM7_s
+ N_VSS_XI1/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM8 N_XI2/NET35_XI2/MM8_d N_WL1_XI2/MM8_g N_BLN<13>_XI2/MM8_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI2/MM5 N_XI2/NET34_XI2/MM5_d N_XI2/NET33_XI2/MM5_g N_VDD_XI2/MM5_s
+ N_VDD_XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI2/MM4 N_XI2/NET33_XI2/MM4_d N_XI2/NET34_XI2/MM4_g N_VDD_XI2/MM4_s
+ N_VDD_XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI2/MM10 N_XI2/NET35_XI2/MM10_d N_XI2/NET36_XI2/MM10_g N_VDD_XI2/MM10_s
+ N_VDD_XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI2/MM11 N_XI2/NET36_XI2/MM11_d N_XI2/NET35_XI2/MM11_g N_VDD_XI2/MM11_s
+ N_VDD_XI2/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI3/MM2 N_XI3/NET34_XI3/MM2_d N_XI3/NET33_XI3/MM2_g N_VSS_XI3/MM2_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM3 N_XI3/NET33_XI3/MM3_d N_WL0_XI3/MM3_g N_BLN<12>_XI3/MM3_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM0 N_XI3/NET34_XI3/MM0_d N_WL0_XI3/MM0_g N_BL<12>_XI3/MM0_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM1 N_XI3/NET33_XI3/MM1_d N_XI3/NET34_XI3/MM1_g N_VSS_XI3/MM1_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM9 N_XI3/NET36_XI3/MM9_d N_WL1_XI3/MM9_g N_BL<12>_XI3/MM9_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM6 N_XI3/NET35_XI3/MM6_d N_XI3/NET36_XI3/MM6_g N_VSS_XI3/MM6_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM7 N_XI3/NET36_XI3/MM7_d N_XI3/NET35_XI3/MM7_g N_VSS_XI3/MM7_s
+ N_VSS_XI2/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM8 N_XI3/NET35_XI3/MM8_d N_WL1_XI3/MM8_g N_BLN<12>_XI3/MM8_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI3/MM5 N_XI3/NET34_XI3/MM5_d N_XI3/NET33_XI3/MM5_g N_VDD_XI3/MM5_s
+ N_VDD_XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI3/MM4 N_XI3/NET33_XI3/MM4_d N_XI3/NET34_XI3/MM4_g N_VDD_XI3/MM4_s
+ N_VDD_XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI3/MM10 N_XI3/NET35_XI3/MM10_d N_XI3/NET36_XI3/MM10_g N_VDD_XI3/MM10_s
+ N_VDD_XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI3/MM11 N_XI3/NET36_XI3/MM11_d N_XI3/NET35_XI3/MM11_g N_VDD_XI3/MM11_s
+ N_VDD_XI3/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/MM2 N_XI4/NET34_XI4/MM2_d N_XI4/NET33_XI4/MM2_g N_VSS_XI4/MM2_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM3 N_XI4/NET33_XI4/MM3_d N_WL0_XI4/MM3_g N_BLN<11>_XI4/MM3_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM0 N_XI4/NET34_XI4/MM0_d N_WL0_XI4/MM0_g N_BL<11>_XI4/MM0_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM1 N_XI4/NET33_XI4/MM1_d N_XI4/NET34_XI4/MM1_g N_VSS_XI4/MM1_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM9 N_XI4/NET36_XI4/MM9_d N_WL1_XI4/MM9_g N_BL<11>_XI4/MM9_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM6 N_XI4/NET35_XI4/MM6_d N_XI4/NET36_XI4/MM6_g N_VSS_XI4/MM6_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM7 N_XI4/NET36_XI4/MM7_d N_XI4/NET35_XI4/MM7_g N_VSS_XI4/MM7_s
+ N_VSS_XI3/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM8 N_XI4/NET35_XI4/MM8_d N_WL1_XI4/MM8_g N_BLN<11>_XI4/MM8_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI4/MM5 N_XI4/NET34_XI4/MM5_d N_XI4/NET33_XI4/MM5_g N_VDD_XI4/MM5_s
+ N_VDD_XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/MM4 N_XI4/NET33_XI4/MM4_d N_XI4/NET34_XI4/MM4_g N_VDD_XI4/MM4_s
+ N_VDD_XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/MM10 N_XI4/NET35_XI4/MM10_d N_XI4/NET36_XI4/MM10_g N_VDD_XI4/MM10_s
+ N_VDD_XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI4/MM11 N_XI4/NET36_XI4/MM11_d N_XI4/NET35_XI4/MM11_g N_VDD_XI4/MM11_s
+ N_VDD_XI4/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/MM2 N_XI5/NET34_XI5/MM2_d N_XI5/NET33_XI5/MM2_g N_VSS_XI5/MM2_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM3 N_XI5/NET33_XI5/MM3_d N_WL0_XI5/MM3_g N_BLN<10>_XI5/MM3_s
+ N_VSS_XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM0 N_XI5/NET34_XI5/MM0_d N_WL0_XI5/MM0_g N_BL<10>_XI5/MM0_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM1 N_XI5/NET33_XI5/MM1_d N_XI5/NET34_XI5/MM1_g N_VSS_XI5/MM1_s
+ N_VSS_XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM9 N_XI5/NET36_XI5/MM9_d N_WL1_XI5/MM9_g N_BL<10>_XI5/MM9_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM6 N_XI5/NET35_XI5/MM6_d N_XI5/NET36_XI5/MM6_g N_VSS_XI5/MM6_s
+ N_VSS_XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM7 N_XI5/NET36_XI5/MM7_d N_XI5/NET35_XI5/MM7_g N_VSS_XI5/MM7_s
+ N_VSS_XI4/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM8 N_XI5/NET35_XI5/MM8_d N_WL1_XI5/MM8_g N_BLN<10>_XI5/MM8_s
+ N_VSS_XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI5/MM5 N_XI5/NET34_XI5/MM5_d N_XI5/NET33_XI5/MM5_g N_VDD_XI5/MM5_s
+ N_VDD_XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/MM4 N_XI5/NET33_XI5/MM4_d N_XI5/NET34_XI5/MM4_g N_VDD_XI5/MM4_s
+ N_VDD_XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/MM10 N_XI5/NET35_XI5/MM10_d N_XI5/NET36_XI5/MM10_g N_VDD_XI5/MM10_s
+ N_VDD_XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI5/MM11 N_XI5/NET36_XI5/MM11_d N_XI5/NET35_XI5/MM11_g N_VDD_XI5/MM11_s
+ N_VDD_XI5/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/MM2 N_XI6/NET34_XI6/MM2_d N_XI6/NET33_XI6/MM2_g N_VSS_XI6/MM2_s
+ N_VSS_XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM3 N_XI6/NET33_XI6/MM3_d N_WL0_XI6/MM3_g N_BLN<9>_XI6/MM3_s
+ N_VSS_XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM0 N_XI6/NET34_XI6/MM0_d N_WL0_XI6/MM0_g N_BL<9>_XI6/MM0_s N_VSS_XI5/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM1 N_XI6/NET33_XI6/MM1_d N_XI6/NET34_XI6/MM1_g N_VSS_XI6/MM1_s
+ N_VSS_XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM9 N_XI6/NET36_XI6/MM9_d N_WL1_XI6/MM9_g N_BL<9>_XI6/MM9_s N_VSS_XI5/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM6 N_XI6/NET35_XI6/MM6_d N_XI6/NET36_XI6/MM6_g N_VSS_XI6/MM6_s
+ N_VSS_XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM7 N_XI6/NET36_XI6/MM7_d N_XI6/NET35_XI6/MM7_g N_VSS_XI6/MM7_s
+ N_VSS_XI5/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM8 N_XI6/NET35_XI6/MM8_d N_WL1_XI6/MM8_g N_BLN<9>_XI6/MM8_s
+ N_VSS_XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI6/MM5 N_XI6/NET34_XI6/MM5_d N_XI6/NET33_XI6/MM5_g N_VDD_XI6/MM5_s
+ N_VDD_XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/MM4 N_XI6/NET33_XI6/MM4_d N_XI6/NET34_XI6/MM4_g N_VDD_XI6/MM4_s
+ N_VDD_XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/MM10 N_XI6/NET35_XI6/MM10_d N_XI6/NET36_XI6/MM10_g N_VDD_XI6/MM10_s
+ N_VDD_XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI6/MM11 N_XI6/NET36_XI6/MM11_d N_XI6/NET35_XI6/MM11_g N_VDD_XI6/MM11_s
+ N_VDD_XI6/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/MM2 N_XI7/NET34_XI7/MM2_d N_XI7/NET33_XI7/MM2_g N_VSS_XI7/MM2_s
+ N_VSS_XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM3 N_XI7/NET33_XI7/MM3_d N_WL0_XI7/MM3_g N_BLN<8>_XI7/MM3_s
+ N_VSS_XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM0 N_XI7/NET34_XI7/MM0_d N_WL0_XI7/MM0_g N_BL<8>_XI7/MM0_s N_VSS_XI6/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM1 N_XI7/NET33_XI7/MM1_d N_XI7/NET34_XI7/MM1_g N_VSS_XI7/MM1_s
+ N_VSS_XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM9 N_XI7/NET36_XI7/MM9_d N_WL1_XI7/MM9_g N_BL<8>_XI7/MM9_s N_VSS_XI6/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM6 N_XI7/NET35_XI7/MM6_d N_XI7/NET36_XI7/MM6_g N_VSS_XI7/MM6_s
+ N_VSS_XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM7 N_XI7/NET36_XI7/MM7_d N_XI7/NET35_XI7/MM7_g N_VSS_XI7/MM7_s
+ N_VSS_XI6/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM8 N_XI7/NET35_XI7/MM8_d N_WL1_XI7/MM8_g N_BLN<8>_XI7/MM8_s
+ N_VSS_XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI7/MM5 N_XI7/NET34_XI7/MM5_d N_XI7/NET33_XI7/MM5_g N_VDD_XI7/MM5_s
+ N_VDD_XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/MM4 N_XI7/NET33_XI7/MM4_d N_XI7/NET34_XI7/MM4_g N_VDD_XI7/MM4_s
+ N_VDD_XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/MM10 N_XI7/NET35_XI7/MM10_d N_XI7/NET36_XI7/MM10_g N_VDD_XI7/MM10_s
+ N_VDD_XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI7/MM11 N_XI7/NET36_XI7/MM11_d N_XI7/NET35_XI7/MM11_g N_VDD_XI7/MM11_s
+ N_VDD_XI7/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/MM2 N_XI8/NET34_XI8/MM2_d N_XI8/NET33_XI8/MM2_g N_VSS_XI8/MM2_s
+ N_VSS_XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM3 N_XI8/NET33_XI8/MM3_d N_WL0_XI8/MM3_g N_BLN<7>_XI8/MM3_s
+ N_VSS_XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM0 N_XI8/NET34_XI8/MM0_d N_WL0_XI8/MM0_g N_BL<7>_XI8/MM0_s N_VSS_XI7/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM1 N_XI8/NET33_XI8/MM1_d N_XI8/NET34_XI8/MM1_g N_VSS_XI8/MM1_s
+ N_VSS_XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM9 N_XI8/NET36_XI8/MM9_d N_WL1_XI8/MM9_g N_BL<7>_XI8/MM9_s N_VSS_XI7/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM6 N_XI8/NET35_XI8/MM6_d N_XI8/NET36_XI8/MM6_g N_VSS_XI8/MM6_s
+ N_VSS_XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM7 N_XI8/NET36_XI8/MM7_d N_XI8/NET35_XI8/MM7_g N_VSS_XI8/MM7_s
+ N_VSS_XI7/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM8 N_XI8/NET35_XI8/MM8_d N_WL1_XI8/MM8_g N_BLN<7>_XI8/MM8_s
+ N_VSS_XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI8/MM5 N_XI8/NET34_XI8/MM5_d N_XI8/NET33_XI8/MM5_g N_VDD_XI8/MM5_s
+ N_VDD_XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/MM4 N_XI8/NET33_XI8/MM4_d N_XI8/NET34_XI8/MM4_g N_VDD_XI8/MM4_s
+ N_VDD_XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/MM10 N_XI8/NET35_XI8/MM10_d N_XI8/NET36_XI8/MM10_g N_VDD_XI8/MM10_s
+ N_VDD_XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI8/MM11 N_XI8/NET36_XI8/MM11_d N_XI8/NET35_XI8/MM11_g N_VDD_XI8/MM11_s
+ N_VDD_XI8/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/MM2 N_XI9/NET34_XI9/MM2_d N_XI9/NET33_XI9/MM2_g N_VSS_XI9/MM2_s
+ N_VSS_XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM3 N_XI9/NET33_XI9/MM3_d N_WL0_XI9/MM3_g N_BLN<6>_XI9/MM3_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM0 N_XI9/NET34_XI9/MM0_d N_WL0_XI9/MM0_g N_BL<6>_XI9/MM0_s N_VSS_XI8/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM1 N_XI9/NET33_XI9/MM1_d N_XI9/NET34_XI9/MM1_g N_VSS_XI9/MM1_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM9 N_XI9/NET36_XI9/MM9_d N_WL1_XI9/MM9_g N_BL<6>_XI9/MM9_s N_VSS_XI8/MM3_b
+ NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM6 N_XI9/NET35_XI9/MM6_d N_XI9/NET36_XI9/MM6_g N_VSS_XI9/MM6_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM7 N_XI9/NET36_XI9/MM7_d N_XI9/NET35_XI9/MM7_g N_VSS_XI9/MM7_s
+ N_VSS_XI8/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM8 N_XI9/NET35_XI9/MM8_d N_WL1_XI9/MM8_g N_BLN<6>_XI9/MM8_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI9/MM5 N_XI9/NET34_XI9/MM5_d N_XI9/NET33_XI9/MM5_g N_VDD_XI9/MM5_s
+ N_VDD_XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/MM4 N_XI9/NET33_XI9/MM4_d N_XI9/NET34_XI9/MM4_g N_VDD_XI9/MM4_s
+ N_VDD_XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/MM10 N_XI9/NET35_XI9/MM10_d N_XI9/NET36_XI9/MM10_g N_VDD_XI9/MM10_s
+ N_VDD_XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI9/MM11 N_XI9/NET36_XI9/MM11_d N_XI9/NET35_XI9/MM11_g N_VDD_XI9/MM11_s
+ N_VDD_XI9/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/MM2 N_XI10/NET34_XI10/MM2_d N_XI10/NET33_XI10/MM2_g N_VSS_XI10/MM2_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM3 N_XI10/NET33_XI10/MM3_d N_WL0_XI10/MM3_g N_BLN<5>_XI10/MM3_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM0 N_XI10/NET34_XI10/MM0_d N_WL0_XI10/MM0_g N_BL<5>_XI10/MM0_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM1 N_XI10/NET33_XI10/MM1_d N_XI10/NET34_XI10/MM1_g N_VSS_XI10/MM1_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM9 N_XI10/NET36_XI10/MM9_d N_WL1_XI10/MM9_g N_BL<5>_XI10/MM9_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM6 N_XI10/NET35_XI10/MM6_d N_XI10/NET36_XI10/MM6_g N_VSS_XI10/MM6_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM7 N_XI10/NET36_XI10/MM7_d N_XI10/NET35_XI10/MM7_g N_VSS_XI10/MM7_s
+ N_VSS_XI9/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM8 N_XI10/NET35_XI10/MM8_d N_WL1_XI10/MM8_g N_BLN<5>_XI10/MM8_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI10/MM5 N_XI10/NET34_XI10/MM5_d N_XI10/NET33_XI10/MM5_g N_VDD_XI10/MM5_s
+ N_VDD_XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/MM4 N_XI10/NET33_XI10/MM4_d N_XI10/NET34_XI10/MM4_g N_VDD_XI10/MM4_s
+ N_VDD_XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/MM10 N_XI10/NET35_XI10/MM10_d N_XI10/NET36_XI10/MM10_g N_VDD_XI10/MM10_s
+ N_VDD_XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI10/MM11 N_XI10/NET36_XI10/MM11_d N_XI10/NET35_XI10/MM11_g N_VDD_XI10/MM11_s
+ N_VDD_XI10/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/MM2 N_XI11/NET34_XI11/MM2_d N_XI11/NET33_XI11/MM2_g N_VSS_XI11/MM2_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM3 N_XI11/NET33_XI11/MM3_d N_WL0_XI11/MM3_g N_BLN<4>_XI11/MM3_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM0 N_XI11/NET34_XI11/MM0_d N_WL0_XI11/MM0_g N_BL<4>_XI11/MM0_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM1 N_XI11/NET33_XI11/MM1_d N_XI11/NET34_XI11/MM1_g N_VSS_XI11/MM1_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM9 N_XI11/NET36_XI11/MM9_d N_WL1_XI11/MM9_g N_BL<4>_XI11/MM9_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM6 N_XI11/NET35_XI11/MM6_d N_XI11/NET36_XI11/MM6_g N_VSS_XI11/MM6_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM7 N_XI11/NET36_XI11/MM7_d N_XI11/NET35_XI11/MM7_g N_VSS_XI11/MM7_s
+ N_VSS_XI10/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM8 N_XI11/NET35_XI11/MM8_d N_WL1_XI11/MM8_g N_BLN<4>_XI11/MM8_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI11/MM5 N_XI11/NET34_XI11/MM5_d N_XI11/NET33_XI11/MM5_g N_VDD_XI11/MM5_s
+ N_VDD_XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/MM4 N_XI11/NET33_XI11/MM4_d N_XI11/NET34_XI11/MM4_g N_VDD_XI11/MM4_s
+ N_VDD_XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/MM10 N_XI11/NET35_XI11/MM10_d N_XI11/NET36_XI11/MM10_g N_VDD_XI11/MM10_s
+ N_VDD_XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI11/MM11 N_XI11/NET36_XI11/MM11_d N_XI11/NET35_XI11/MM11_g N_VDD_XI11/MM11_s
+ N_VDD_XI11/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/MM2 N_XI12/NET34_XI12/MM2_d N_XI12/NET33_XI12/MM2_g N_VSS_XI12/MM2_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM3 N_XI12/NET33_XI12/MM3_d N_WL0_XI12/MM3_g N_BLN<3>_XI12/MM3_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM0 N_XI12/NET34_XI12/MM0_d N_WL0_XI12/MM0_g N_BL<3>_XI12/MM0_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM1 N_XI12/NET33_XI12/MM1_d N_XI12/NET34_XI12/MM1_g N_VSS_XI12/MM1_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM9 N_XI12/NET36_XI12/MM9_d N_WL1_XI12/MM9_g N_BL<3>_XI12/MM9_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM6 N_XI12/NET35_XI12/MM6_d N_XI12/NET36_XI12/MM6_g N_VSS_XI12/MM6_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM7 N_XI12/NET36_XI12/MM7_d N_XI12/NET35_XI12/MM7_g N_VSS_XI12/MM7_s
+ N_VSS_XI11/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM8 N_XI12/NET35_XI12/MM8_d N_WL1_XI12/MM8_g N_BLN<3>_XI12/MM8_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI12/MM5 N_XI12/NET34_XI12/MM5_d N_XI12/NET33_XI12/MM5_g N_VDD_XI12/MM5_s
+ N_VDD_XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/MM4 N_XI12/NET33_XI12/MM4_d N_XI12/NET34_XI12/MM4_g N_VDD_XI12/MM4_s
+ N_VDD_XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/MM10 N_XI12/NET35_XI12/MM10_d N_XI12/NET36_XI12/MM10_g N_VDD_XI12/MM10_s
+ N_VDD_XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI12/MM11 N_XI12/NET36_XI12/MM11_d N_XI12/NET35_XI12/MM11_g N_VDD_XI12/MM11_s
+ N_VDD_XI12/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/MM2 N_XI13/NET34_XI13/MM2_d N_XI13/NET33_XI13/MM2_g N_VSS_XI13/MM2_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM3 N_XI13/NET33_XI13/MM3_d N_WL0_XI13/MM3_g N_BLN<2>_XI13/MM3_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM0 N_XI13/NET34_XI13/MM0_d N_WL0_XI13/MM0_g N_BL<2>_XI13/MM0_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM1 N_XI13/NET33_XI13/MM1_d N_XI13/NET34_XI13/MM1_g N_VSS_XI13/MM1_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM9 N_XI13/NET36_XI13/MM9_d N_WL1_XI13/MM9_g N_BL<2>_XI13/MM9_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM6 N_XI13/NET35_XI13/MM6_d N_XI13/NET36_XI13/MM6_g N_VSS_XI13/MM6_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM7 N_XI13/NET36_XI13/MM7_d N_XI13/NET35_XI13/MM7_g N_VSS_XI13/MM7_s
+ N_VSS_XI12/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM8 N_XI13/NET35_XI13/MM8_d N_WL1_XI13/MM8_g N_BLN<2>_XI13/MM8_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI13/MM5 N_XI13/NET34_XI13/MM5_d N_XI13/NET33_XI13/MM5_g N_VDD_XI13/MM5_s
+ N_VDD_XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/MM4 N_XI13/NET33_XI13/MM4_d N_XI13/NET34_XI13/MM4_g N_VDD_XI13/MM4_s
+ N_VDD_XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/MM10 N_XI13/NET35_XI13/MM10_d N_XI13/NET36_XI13/MM10_g N_VDD_XI13/MM10_s
+ N_VDD_XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI13/MM11 N_XI13/NET36_XI13/MM11_d N_XI13/NET35_XI13/MM11_g N_VDD_XI13/MM11_s
+ N_VDD_XI13/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/MM2 N_XI14/NET34_XI14/MM2_d N_XI14/NET33_XI14/MM2_g N_VSS_XI14/MM2_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM3 N_XI14/NET33_XI14/MM3_d N_WL0_XI14/MM3_g N_BLN<1>_XI14/MM3_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM0 N_XI14/NET34_XI14/MM0_d N_WL0_XI14/MM0_g N_BL<1>_XI14/MM0_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM1 N_XI14/NET33_XI14/MM1_d N_XI14/NET34_XI14/MM1_g N_VSS_XI14/MM1_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM9 N_XI14/NET36_XI14/MM9_d N_WL1_XI14/MM9_g N_BL<1>_XI14/MM9_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM6 N_XI14/NET35_XI14/MM6_d N_XI14/NET36_XI14/MM6_g N_VSS_XI14/MM6_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM7 N_XI14/NET36_XI14/MM7_d N_XI14/NET35_XI14/MM7_g N_VSS_XI14/MM7_s
+ N_VSS_XI13/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM8 N_XI14/NET35_XI14/MM8_d N_WL1_XI14/MM8_g N_BLN<1>_XI14/MM8_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI14/MM5 N_XI14/NET34_XI14/MM5_d N_XI14/NET33_XI14/MM5_g N_VDD_XI14/MM5_s
+ N_VDD_XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/MM4 N_XI14/NET33_XI14/MM4_d N_XI14/NET34_XI14/MM4_g N_VDD_XI14/MM4_s
+ N_VDD_XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/MM10 N_XI14/NET35_XI14/MM10_d N_XI14/NET36_XI14/MM10_g N_VDD_XI14/MM10_s
+ N_VDD_XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI14/MM11 N_XI14/NET36_XI14/MM11_d N_XI14/NET35_XI14/MM11_g N_VDD_XI14/MM11_s
+ N_VDD_XI14/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/MM2 N_XI15/NET34_XI15/MM2_d N_XI15/NET33_XI15/MM2_g N_VSS_XI15/MM2_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM3 N_XI15/NET33_XI15/MM3_d N_WL0_XI15/MM3_g N_BLN<0>_XI15/MM3_s
+ N_VSS_XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM0 N_XI15/NET34_XI15/MM0_d N_WL0_XI15/MM0_g N_BL<0>_XI15/MM0_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM1 N_XI15/NET33_XI15/MM1_d N_XI15/NET34_XI15/MM1_g N_VSS_XI15/MM1_s
+ N_VSS_XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM9 N_XI15/NET36_XI15/MM9_d N_WL1_XI15/MM9_g N_BL<0>_XI15/MM9_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM6 N_XI15/NET35_XI15/MM6_d N_XI15/NET36_XI15/MM6_g N_VSS_XI15/MM6_s
+ N_VSS_XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM7 N_XI15/NET36_XI15/MM7_d N_XI15/NET35_XI15/MM7_g N_VSS_XI15/MM7_s
+ N_VSS_XI14/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM8 N_XI15/NET35_XI15/MM8_d N_WL1_XI15/MM8_g N_BLN<0>_XI15/MM8_s
+ N_VSS_XI15/MM3_b NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
mXI15/MM5 N_XI15/NET34_XI15/MM5_d N_XI15/NET33_XI15/MM5_g N_VDD_XI15/MM5_s
+ N_VDD_XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/MM4 N_XI15/NET33_XI15/MM4_d N_XI15/NET34_XI15/MM4_g N_VDD_XI15/MM4_s
+ N_VDD_XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/MM10 N_XI15/NET35_XI15/MM10_d N_XI15/NET36_XI15/MM10_g N_VDD_XI15/MM10_s
+ N_VDD_XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
mXI15/MM11 N_XI15/NET36_XI15/MM11_d N_XI15/NET35_XI15/MM11_g N_VDD_XI15/MM11_s
+ N_VDD_XI15/MM5_b PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
*
.include "netlist.sp.SRAM_16B_2.pxi"
*
.ends
*
*
