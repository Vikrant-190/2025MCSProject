* File: netlist.sp
* Created: Wed Jun 11 22:23:12 2025
* Program "Calibre xRC"
* Version "v2019.2_26.18"
* 
.include "netlist.sp.pex"
.subckt sram_4  WL BL VSS VDD BLN
* 
* BLN	BLN
* VDD	VDD
* VSS	VSS
* BL	BL
* WL	WL
MM0 N_NET20_MM0_d N_WL_MM0_g N_BL_MM0_s N_VSS_MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
MM1 N_NET19_MM1_d N_NET20_MM1_g N_VSS_MM1_s N_VSS_MM0_b NMOS_SRAM L=2e-08
+ W=5.4e-08 NFIN=2
MM2 N_NET20_MM2_d N_NET19_MM2_g N_VSS_MM2_s N_VSS_MM0_b NMOS_SRAM L=2e-08
+ W=5.4e-08 NFIN=2
MM3 N_NET19_MM3_d N_WL_MM3_g N_BLN_MM3_s N_VSS_MM0_b NMOS_SRAM L=2e-08 W=5.4e-08
+ NFIN=2
MM4 N_NET19_MM4_d N_NET20_MM4_g N_VDD_MM4_s N_VDD_MM4_b PMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
MM5 N_NET20_MM5_d N_NET19_MM5_g N_VDD_MM5_s N_VDD_MM4_b PMOS_SRAM L=2e-08
+ W=2.7e-08 NFIN=1
*
.include "netlist.sp.SRAM_4.pxi"
*
.ends
*
*
